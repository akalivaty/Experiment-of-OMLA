//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  OAI21_X1  g000(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g003(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT66), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207));
  NAND4_X1  g006(.A1(new_n207), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n211));
  AND2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n214), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT25), .B1(new_n209), .B2(new_n216), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n205), .A2(KEYINPUT64), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n221), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n219), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT26), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n228), .B(new_n203), .C1(new_n230), .C2(new_n212), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT28), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n237));
  OAI211_X1 g036(.A(KEYINPUT28), .B(new_n234), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n232), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n231), .B1(new_n244), .B2(new_n238), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n225), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249));
  OAI21_X1  g048(.A(G127gat), .B1(new_n249), .B2(KEYINPUT1), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G113gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G120gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(G127gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n250), .A2(new_n258), .A3(G134gat), .ZN(new_n259));
  AOI21_X1  g058(.A(G134gat), .B1(new_n250), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT68), .B1(new_n248), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n247), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n223), .A2(new_n219), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(new_n216), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n219), .B1(new_n218), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND4_X1   g067(.A1(KEYINPUT68), .A2(new_n263), .A3(new_n261), .A4(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT34), .B1(new_n272), .B2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n249), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n257), .B1(new_n255), .B2(new_n256), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n250), .A2(new_n258), .A3(G134gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n245), .A2(new_n246), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT67), .B(new_n231), .C1(new_n244), .C2(new_n238), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n279), .B1(new_n282), .B2(new_n225), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n270), .A2(new_n271), .A3(new_n273), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n273), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n268), .B(new_n261), .C1(new_n280), .C2(new_n281), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n263), .A2(KEYINPUT68), .A3(new_n261), .A4(new_n268), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n285), .B1(new_n290), .B2(new_n272), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n272), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT69), .B(G71gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G99gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G15gat), .B(G43gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n296), .B1(new_n290), .B2(new_n272), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT70), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n303), .A2(new_n295), .ZN(new_n310));
  AOI211_X1 g109(.A(new_n309), .B(new_n310), .C1(new_n290), .C2(new_n272), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n293), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g112(.A(new_n311), .B(new_n292), .C1(new_n305), .C2(new_n307), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G78gat), .B(G106gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n316), .B(G22gat), .Z(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT31), .B(G50gat), .ZN(new_n318));
  AND2_X1   g117(.A1(G228gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  OR2_X1    g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  INV_X1    g121(.A(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G141gat), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G148gat), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n321), .B(new_n322), .C1(new_n327), .C2(KEYINPUT2), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT76), .B1(new_n323), .B2(G141gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n325), .A3(G148gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n331), .A3(new_n324), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n321), .B1(new_n322), .B2(KEYINPUT2), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n332), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT73), .B(G211gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT22), .B1(new_n340), .B2(G218gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(G211gat), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G211gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT73), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G211gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n348), .A3(G218gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT22), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n345), .A3(new_n342), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n344), .A2(G218gat), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(G218gat), .B1(new_n344), .B2(new_n352), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n339), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n338), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(new_n352), .ZN(new_n358));
  INV_X1    g157(.A(G218gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n344), .A2(G218gat), .A3(new_n352), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT82), .B1(new_n362), .B2(new_n339), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n337), .B1(new_n357), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n365));
  NAND2_X1  g164(.A1(new_n332), .A2(new_n333), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT77), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT2), .B1(new_n324), .B2(new_n326), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(G155gat), .B2(G162gat), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n367), .A2(new_n368), .B1(new_n370), .B2(new_n322), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n365), .B1(new_n371), .B2(new_n338), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n320), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n365), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT3), .B1(new_n362), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n374), .B(new_n320), .C1(new_n377), .C2(new_n371), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n318), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n318), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n355), .A2(new_n356), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n362), .A2(KEYINPUT82), .A3(new_n339), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n338), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n373), .B1(new_n384), .B2(new_n337), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n378), .B(new_n381), .C1(new_n385), .C2(new_n320), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n317), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(new_n317), .A3(new_n386), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n315), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n337), .A2(KEYINPUT3), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n338), .B(new_n328), .C1(new_n335), .C2(new_n336), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n279), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n367), .A2(new_n368), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n396), .A2(new_n278), .A3(new_n277), .A4(new_n328), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n261), .B2(new_n371), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n395), .B(new_n399), .C1(new_n402), .C2(new_n398), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n279), .A2(new_n337), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n397), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n406), .B2(new_n401), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n401), .A2(KEYINPUT5), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n412));
  NAND3_X1  g211(.A1(new_n261), .A2(new_n371), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n395), .A2(new_n410), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G29gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(G1gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND3_X1  g219(.A1(new_n408), .A2(new_n414), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n408), .B2(new_n414), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n392), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(KEYINPUT6), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n414), .ZN(new_n427));
  INV_X1    g226(.A(new_n420), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(KEYINPUT81), .A3(new_n422), .A4(new_n421), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT75), .ZN(new_n434));
  INV_X1    g233(.A(G8gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n248), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n339), .B(new_n437), .C1(new_n225), .C2(new_n245), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n362), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n376), .B(new_n437), .C1(new_n282), .C2(new_n225), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n268), .A2(new_n240), .A3(new_n438), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n362), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n436), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n436), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n443), .A2(new_n444), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n441), .B(new_n447), .C1(new_n448), .C2(new_n362), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n449), .A3(KEYINPUT30), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n441), .B1(new_n448), .B2(new_n362), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n436), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n431), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT35), .B1(new_n391), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n395), .A2(new_n410), .A3(new_n413), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n411), .A2(new_n457), .B1(new_n403), .B2(new_n407), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT6), .B1(new_n458), .B2(new_n420), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT84), .B1(new_n427), .B2(new_n428), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n461), .B(new_n420), .C1(new_n408), .C2(new_n414), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT86), .B(new_n459), .C1(new_n460), .C2(new_n462), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n426), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n454), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n299), .B1(new_n298), .B2(new_n304), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n306), .A2(KEYINPUT70), .A3(new_n303), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n312), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n292), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n308), .A2(new_n293), .A3(new_n312), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n380), .A2(new_n317), .A3(new_n386), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(new_n387), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n467), .A2(new_n480), .A3(new_n454), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n469), .A2(new_n470), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n466), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n461), .B1(new_n458), .B2(new_n420), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n424), .A2(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT86), .B1(new_n486), .B2(new_n459), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n436), .B1(new_n451), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n448), .B2(new_n362), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n439), .A2(new_n440), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n362), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n489), .B1(new_n442), .B2(new_n445), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT37), .B(new_n441), .C1(new_n448), .C2(new_n362), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n447), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n498), .A2(KEYINPUT38), .B1(new_n451), .B2(new_n436), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n488), .A2(new_n426), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n395), .A2(new_n410), .A3(new_n413), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n401), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n420), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(KEYINPUT83), .A3(new_n420), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n401), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(KEYINPUT39), .C1(new_n401), .C2(new_n406), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT40), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n460), .A2(new_n462), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n511), .A2(new_n454), .A3(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n503), .A2(KEYINPUT83), .A3(new_n420), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT83), .B1(new_n503), .B2(new_n420), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT40), .B(new_n510), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n513), .A2(new_n518), .B1(new_n389), .B2(new_n388), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n500), .A2(new_n519), .B1(new_n478), .B2(new_n455), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n313), .B2(new_n314), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n476), .A2(new_n521), .A3(KEYINPUT36), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n456), .A2(new_n482), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G230gat), .A2(G233gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT96), .Z(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n531), .A2(KEYINPUT9), .ZN(new_n532));
  XNOR2_X1  g331(.A(G71gat), .B(G78gat), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT92), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(KEYINPUT92), .ZN(new_n537));
  OAI22_X1  g336(.A1(new_n532), .A2(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  INV_X1    g338(.A(G85gat), .ZN(new_n540));
  INV_X1    g339(.A(G92gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT7), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n540), .B2(new_n541), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n539), .B(new_n547), .C1(new_n540), .C2(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G99gat), .B(G106gat), .Z(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n538), .B1(new_n551), .B2(KEYINPUT95), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n550), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n552), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT10), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR3_X1    g356(.A1(new_n554), .A2(new_n556), .A3(new_n538), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n529), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n559), .A2(KEYINPUT97), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(KEYINPUT97), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n227), .ZN(new_n564));
  INV_X1    g363(.A(G204gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568));
  INV_X1    g367(.A(new_n555), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(new_n529), .ZN(new_n570));
  INV_X1    g369(.A(new_n529), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n555), .A2(KEYINPUT98), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n562), .A2(KEYINPUT99), .A3(new_n567), .A4(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n567), .B(new_n573), .C1(new_n560), .C2(new_n561), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n559), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n578), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n574), .A2(new_n577), .B1(new_n566), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G43gat), .B(G50gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n586));
  INV_X1    g385(.A(G29gat), .ZN(new_n587));
  INV_X1    g386(.A(G36gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OR3_X1    g388(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT15), .A3(new_n584), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n585), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G15gat), .B(G22gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT16), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(G1gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n435), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(G1gat), .B2(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI221_X1 g403(.A(new_n600), .B1(new_n601), .B2(new_n435), .C1(G1gat), .C2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n597), .B(KEYINPUT17), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n604), .A2(new_n605), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n612), .A2(KEYINPUT18), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n597), .B(new_n606), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n611), .B(KEYINPUT13), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(KEYINPUT18), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT89), .ZN(new_n620));
  XOR2_X1   g419(.A(G113gat), .B(G141gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G169gat), .B(G197gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n613), .A2(new_n627), .A3(new_n616), .A4(new_n617), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n583), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n609), .B1(new_n631), .B2(new_n538), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G183gat), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n633), .A2(KEYINPUT93), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(KEYINPUT93), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n634), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n345), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n633), .B(KEYINPUT93), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n635), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n646), .B2(new_n638), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n538), .A2(new_n631), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n643), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n646), .A2(new_n638), .A3(new_n644), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n608), .A2(new_n554), .ZN(new_n657));
  INV_X1    g456(.A(new_n554), .ZN(new_n658));
  AND2_X1   g457(.A1(G232gat), .A2(G233gat), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n658), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G134gat), .B(G162gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n659), .A2(KEYINPUT41), .ZN(new_n664));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n663), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n656), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n527), .A2(new_n630), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n431), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT101), .B(G1gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1324gat));
  INV_X1    g473(.A(new_n454), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n599), .B2(new_n435), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n599), .B2(new_n435), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n678), .A2(KEYINPUT102), .A3(new_n679), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n678), .A2(new_n679), .B1(G8gat), .B2(new_n676), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT102), .B1(new_n678), .B2(new_n679), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(G15gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n670), .A2(new_n684), .A3(new_n315), .ZN(new_n685));
  INV_X1    g484(.A(new_n526), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n670), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n687), .B2(new_n684), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT103), .Z(G1326gat));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n478), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NOR4_X1   g491(.A1(new_n527), .A2(new_n630), .A3(new_n656), .A4(new_n668), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n587), .A3(new_n671), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n482), .A2(new_n456), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n520), .A2(new_n526), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n668), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(KEYINPUT104), .B(KEYINPUT44), .C1(new_n527), .C2(new_n668), .ZN(new_n702));
  INV_X1    g501(.A(new_n455), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n470), .B1(new_n479), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n391), .B1(KEYINPUT87), .B2(new_n468), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n481), .A2(new_n470), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n516), .A2(KEYINPUT85), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n454), .A2(new_n512), .ZN(new_n709));
  INV_X1    g508(.A(new_n511), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n516), .A2(KEYINPUT85), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n495), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n465), .A2(new_n426), .A3(new_n466), .A4(new_n499), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n712), .B(new_n390), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT105), .B1(new_n703), .B2(new_n390), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n478), .A2(new_n455), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n524), .A2(new_n525), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT106), .B1(new_n707), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n697), .B(new_n723), .C1(new_n720), .C2(new_n717), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n701), .A2(new_n702), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(new_n630), .A3(new_n656), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n671), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n695), .B1(new_n729), .B2(new_n587), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n693), .A2(new_n588), .A3(new_n675), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n734), .A2(new_n733), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n728), .A2(new_n675), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n736), .B(new_n737), .C1(new_n738), .C2(new_n588), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT108), .Z(G1329gat));
  INV_X1    g539(.A(G43gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n728), .B2(new_n686), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n693), .A2(new_n741), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n315), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  INV_X1    g545(.A(G50gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n728), .B2(new_n478), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n693), .A2(new_n747), .A3(new_n478), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT109), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n746), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n748), .A2(new_n746), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n752), .A2(new_n753), .A3(new_n749), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n752), .B2(new_n749), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(G1331gat));
  INV_X1    g555(.A(new_n669), .ZN(new_n757));
  INV_X1    g556(.A(new_n629), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n583), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT111), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n722), .B2(new_n724), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n671), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n675), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT49), .B(G64gat), .Z(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n762), .A2(new_n769), .A3(new_n315), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n762), .B2(new_n686), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT112), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n772), .A2(new_n773), .A3(KEYINPUT50), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT50), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n762), .A2(new_n478), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT113), .B(G78gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1335gat));
  AND3_X1   g578(.A1(new_n524), .A2(new_n525), .A3(new_n719), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n718), .B1(new_n478), .B2(new_n455), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n500), .B2(new_n519), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n456), .A2(new_n482), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n651), .B1(new_n643), .B2(new_n647), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n653), .A2(new_n650), .A3(new_n654), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n787), .B2(new_n758), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT114), .B(new_n629), .C1(new_n785), .C2(new_n786), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n667), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT51), .B1(new_n783), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n574), .A2(new_n577), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n582), .A2(new_n566), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n758), .B1(new_n652), .B2(new_n655), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT114), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n787), .A2(new_n784), .A3(new_n758), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n668), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n798), .B(new_n799), .C1(new_n707), .C2(new_n721), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n791), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n671), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n794), .B1(new_n788), .B2(new_n789), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n701), .A2(new_n702), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n725), .A2(new_n726), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n431), .A2(new_n540), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n802), .B1(new_n806), .B2(new_n807), .ZN(G1336gat));
  AOI21_X1  g607(.A(new_n541), .B1(new_n806), .B2(new_n675), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n800), .A3(new_n675), .A4(new_n794), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(G92gat), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n809), .A2(KEYINPUT52), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT115), .B1(new_n810), .B2(G92gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n801), .A2(new_n814), .A3(new_n541), .A4(new_n675), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n727), .A2(new_n454), .A3(new_n803), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n813), .B(new_n815), .C1(new_n816), .C2(new_n541), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT116), .B1(new_n817), .B2(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n813), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT116), .B(KEYINPUT52), .C1(new_n809), .C2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n812), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT117), .B(new_n812), .C1(new_n818), .C2(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1337gat));
  INV_X1    g625(.A(new_n806), .ZN(new_n827));
  OAI21_X1  g626(.A(G99gat), .B1(new_n827), .B2(new_n526), .ZN(new_n828));
  INV_X1    g627(.A(G99gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n801), .A2(new_n829), .A3(new_n315), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1338gat));
  INV_X1    g630(.A(G106gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n801), .A2(new_n832), .A3(new_n478), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n827), .A2(new_n390), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n832), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n833), .B2(KEYINPUT118), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n835), .B(new_n837), .ZN(G1339gat));
  NOR2_X1   g637(.A1(new_n759), .A2(new_n794), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n610), .A2(new_n611), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n614), .A2(new_n615), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n624), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n628), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n794), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT120), .B1(new_n583), .B2(new_n844), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n557), .A2(new_n529), .A3(new_n558), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT54), .B(new_n848), .C1(new_n560), .C2(new_n561), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  INV_X1    g649(.A(new_n581), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n579), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n852), .A3(new_n566), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n849), .A2(new_n852), .A3(KEYINPUT55), .A4(new_n566), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n792), .A2(new_n855), .A3(new_n629), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n846), .A2(new_n847), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n668), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n792), .A2(new_n855), .A3(new_n845), .A4(new_n856), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT119), .B1(new_n860), .B2(new_n668), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n792), .A2(new_n855), .A3(new_n856), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n667), .A4(new_n845), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n839), .B1(new_n865), .B2(new_n787), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n391), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n671), .A3(new_n454), .ZN(new_n868));
  OAI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n758), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n671), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n253), .A3(new_n454), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n873), .B2(new_n758), .ZN(G1340gat));
  NAND2_X1  g673(.A1(new_n794), .A2(new_n251), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT122), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(new_n454), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G120gat), .B1(new_n868), .B2(new_n583), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1341gat));
  NOR3_X1   g678(.A1(new_n868), .A2(new_n257), .A3(new_n787), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n872), .A2(new_n454), .A3(new_n656), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n257), .ZN(G1342gat));
  NOR2_X1   g681(.A1(new_n668), .A2(G134gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n872), .A2(new_n454), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n868), .B2(new_n668), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n887), .A3(new_n454), .A4(new_n883), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(G1343gat));
  NOR2_X1   g688(.A1(new_n866), .A2(new_n390), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n686), .A2(new_n675), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n671), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n325), .B1(new_n894), .B2(new_n758), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n864), .A2(new_n861), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n794), .A2(new_n845), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n667), .B1(new_n898), .B2(new_n857), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n896), .B(new_n787), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n839), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n857), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n668), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n861), .A3(new_n864), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n896), .B1(new_n905), .B2(new_n787), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n478), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n892), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  INV_X1    g708(.A(new_n897), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n656), .B1(new_n910), .B2(new_n859), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n909), .B(new_n478), .C1(new_n911), .C2(new_n839), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n629), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n895), .B1(new_n913), .B2(new_n325), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT124), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g715(.A1(new_n908), .A2(new_n794), .A3(new_n912), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT57), .B1(new_n866), .B2(new_n390), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n862), .A2(new_n667), .A3(new_n845), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n656), .B1(new_n904), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n909), .B(new_n478), .C1(new_n922), .C2(new_n839), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n920), .A2(new_n794), .A3(new_n893), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G148gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n894), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n323), .A3(new_n794), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(KEYINPUT125), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1345gat));
  AOI21_X1  g733(.A(G155gat), .B1(new_n928), .B2(new_n656), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n908), .A2(G155gat), .A3(new_n912), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n656), .ZN(G1346gat));
  AOI21_X1  g736(.A(G162gat), .B1(new_n928), .B2(new_n667), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n908), .A2(new_n667), .A3(new_n912), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n671), .A2(new_n454), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n867), .A2(new_n941), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n942), .A2(new_n758), .B1(KEYINPUT126), .B2(G169gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(KEYINPUT126), .A2(G169gat), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1348gat));
  NOR2_X1   g744(.A1(new_n942), .A2(new_n583), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(new_n227), .ZN(G1349gat));
  NOR2_X1   g746(.A1(new_n942), .A2(new_n787), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n233), .ZN(new_n949));
  INV_X1    g748(.A(G183gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n948), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g751(.A1(new_n942), .A2(new_n668), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n234), .ZN(new_n955));
  XOR2_X1   g754(.A(KEYINPUT61), .B(G190gat), .Z(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n953), .B2(new_n956), .ZN(G1351gat));
  INV_X1    g756(.A(new_n890), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n526), .A2(new_n941), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(G197gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n961), .A3(new_n629), .ZN(new_n962));
  INV_X1    g761(.A(new_n959), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n920), .A2(new_n923), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n758), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(G1352gat));
  NOR4_X1   g765(.A1(new_n958), .A2(G204gat), .A3(new_n583), .A4(new_n959), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  AND4_X1   g769(.A1(new_n794), .A2(new_n920), .A3(new_n923), .A4(new_n963), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n969), .B(new_n970), .C1(new_n565), .C2(new_n971), .ZN(G1353gat));
  INV_X1    g771(.A(new_n340), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n960), .A2(new_n973), .A3(new_n656), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n920), .A2(new_n656), .A3(new_n923), .A4(new_n963), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n978), .B(new_n979), .ZN(G1354gat));
  NAND3_X1  g779(.A1(new_n960), .A2(new_n359), .A3(new_n667), .ZN(new_n981));
  OAI21_X1  g780(.A(G218gat), .B1(new_n964), .B2(new_n668), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


