//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G134), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT66), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(new_n189), .A3(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT67), .A3(G137), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n191), .A2(G137), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(G134), .B2(new_n189), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n191), .A2(KEYINPUT11), .A3(G137), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n198), .B(new_n199), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n197), .A2(KEYINPUT71), .A3(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  OAI211_X1 g026(.A(G128), .B(new_n209), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n214), .B(new_n215), .C1(KEYINPUT1), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n206), .A2(new_n207), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n220), .B(new_n221), .C1(new_n210), .C2(new_n212), .ZN(new_n222));
  INV_X1    g036(.A(new_n220), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n214), .A3(new_n215), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT70), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n220), .ZN(new_n228));
  XNOR2_X1  g042(.A(G143), .B(G146), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n224), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G131), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n203), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n219), .A2(new_n235), .A3(KEYINPUT30), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n222), .A2(KEYINPUT65), .A3(new_n224), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n218), .A2(new_n203), .A3(new_n197), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT69), .B1(new_n247), .B2(G119), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(G116), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G119), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(KEYINPUT68), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G116), .ZN(new_n254));
  AND4_X1   g068(.A1(new_n251), .A2(new_n252), .A3(new_n254), .A4(G119), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n246), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n254), .A3(G119), .ZN(new_n257));
  INV_X1    g071(.A(new_n248), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n251), .A3(G119), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n245), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n236), .A2(new_n244), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n262), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n219), .A2(new_n235), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G210), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n263), .A2(new_n265), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n264), .B1(new_n241), .B2(new_n240), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n213), .A2(new_n217), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n204), .B2(new_n205), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n277), .A2(new_n207), .B1(new_n231), .B2(new_n234), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT28), .A3(new_n264), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n271), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n187), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n219), .A2(new_n235), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n262), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n265), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(KEYINPUT28), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n265), .A2(new_n274), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n271), .A2(new_n187), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n281), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G472), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n275), .A2(new_n279), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n271), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n271), .B1(new_n278), .B2(new_n264), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n263), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT31), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n263), .A2(new_n299), .A3(new_n296), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n300), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n270), .B1(new_n275), .B2(new_n279), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n299), .B1(new_n263), .B2(new_n296), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n302), .A2(KEYINPUT32), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT73), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n301), .A2(new_n312), .A3(KEYINPUT32), .A4(new_n302), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n293), .A2(new_n305), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G128), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n216), .A2(G119), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G110), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(G128), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n318), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n324), .A2(KEYINPUT78), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(KEYINPUT78), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n323), .A2(KEYINPUT75), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(KEYINPUT75), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n319), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT24), .B(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT77), .B(G125), .ZN(new_n333));
  NOR2_X1   g147(.A1(KEYINPUT16), .A2(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G125), .A2(G140), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n333), .B2(G140), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT16), .ZN(new_n338));
  OAI211_X1 g152(.A(G146), .B(new_n335), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(G125), .A2(G140), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n211), .B1(new_n340), .B2(new_n336), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n332), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(KEYINPUT77), .A2(G125), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT77), .A2(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(G140), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n336), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n333), .A2(new_n334), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n211), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n339), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n318), .A2(new_n323), .A3(new_n321), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G110), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n350), .B(new_n352), .C1(new_n330), .C2(new_n329), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  INV_X1    g169(.A(G953), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n356), .A2(G221), .A3(G234), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n355), .B(new_n357), .Z(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n342), .A2(new_n353), .A3(new_n358), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G234), .B2(new_n291), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G902), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n360), .A2(new_n367), .A3(new_n361), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n291), .A3(new_n361), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n370), .A2(KEYINPUT25), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n363), .B(KEYINPUT74), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n370), .B2(KEYINPUT25), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n314), .A2(KEYINPUT80), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT80), .B1(new_n314), .B2(new_n374), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G214), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G101), .ZN(new_n386));
  AOI21_X1  g200(.A(G101), .B1(new_n379), .B2(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n380), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(KEYINPUT4), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT82), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n385), .A2(KEYINPUT82), .A3(new_n391), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n259), .B2(new_n260), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n316), .A3(G116), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G113), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n256), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n382), .A2(G104), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n379), .A2(G107), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n388), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT83), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n388), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI22_X1  g221(.A1(new_n264), .A2(new_n394), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT86), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT88), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n408), .A2(new_n415), .A3(new_n409), .A4(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n409), .B1(new_n408), .B2(new_n412), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n402), .A2(new_n388), .A3(new_n405), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n405), .B1(new_n402), .B2(new_n388), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n245), .B1(new_n259), .B2(new_n260), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT5), .B1(new_n250), .B2(new_n255), .ZN(new_n424));
  INV_X1    g238(.A(new_n398), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n385), .A2(new_n391), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n385), .A2(KEYINPUT82), .A3(new_n391), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n388), .A2(KEYINPUT4), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n429), .A2(new_n430), .B1(new_n431), .B2(new_n386), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n422), .A2(new_n426), .B1(new_n432), .B2(new_n262), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n419), .B1(new_n433), .B2(new_n411), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n262), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n424), .A2(new_n425), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n422), .A2(new_n436), .A3(new_n256), .ZN(new_n437));
  AND4_X1   g251(.A1(new_n419), .A2(new_n435), .A3(new_n437), .A4(new_n411), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n418), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n333), .B1(new_n213), .B2(new_n217), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n225), .B2(new_n333), .ZN(new_n441));
  INV_X1    g255(.A(G224), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G953), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n441), .B(new_n443), .Z(new_n444));
  NAND3_X1  g258(.A1(new_n417), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n399), .A2(new_n388), .A3(new_n402), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n426), .A2(new_n403), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n411), .B(KEYINPUT8), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n225), .A2(new_n333), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n440), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n440), .A2(new_n451), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n452), .A2(new_n453), .B1(new_n454), .B2(new_n443), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n443), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n441), .B(new_n457), .C1(new_n456), .C2(new_n443), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n449), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT87), .B1(new_n408), .B2(new_n412), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n433), .A2(new_n419), .A3(new_n411), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G210), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT91), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n445), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n445), .B2(new_n463), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n378), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT92), .ZN(new_n470));
  INV_X1    g284(.A(G469), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n356), .A2(G227), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n276), .A2(new_n403), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n213), .A2(new_n402), .A3(new_n388), .A4(new_n217), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n234), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n276), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n422), .A2(new_n483), .B1(new_n482), .B2(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n432), .A2(new_n231), .ZN(new_n485));
  INV_X1    g299(.A(new_n234), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n475), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n475), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n486), .B1(new_n484), .B2(new_n485), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n471), .B1(new_n494), .B2(new_n291), .ZN(new_n495));
  INV_X1    g309(.A(new_n487), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n474), .B1(new_n496), .B2(new_n491), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n404), .A2(new_n218), .A3(KEYINPUT10), .A4(new_n406), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n477), .A2(new_n482), .ZN(new_n499));
  INV_X1    g313(.A(new_n230), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n227), .B1(new_n222), .B2(new_n224), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n498), .B(new_n499), .C1(new_n394), .C2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT84), .B(new_n475), .C1(new_n503), .C2(new_n234), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n481), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT84), .B1(new_n487), .B2(new_n475), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n497), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n471), .A3(new_n291), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n471), .A4(new_n291), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n495), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G221), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT9), .B(G234), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n515), .B2(new_n291), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT81), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G478), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT96), .B1(new_n216), .B2(G143), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n208), .A2(KEYINPUT13), .A3(G128), .ZN(new_n522));
  MUX2_X1   g336(.A(KEYINPUT96), .B(new_n521), .S(new_n522), .Z(new_n523));
  AOI21_X1  g337(.A(KEYINPUT13), .B1(new_n208), .B2(G128), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT95), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n191), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n208), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n216), .A2(G143), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT97), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT97), .B1(new_n527), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n191), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n252), .A2(new_n254), .A3(G122), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n247), .A2(G122), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n532), .A2(new_n382), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n382), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n526), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n527), .A2(new_n528), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT97), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(G134), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n534), .B1(new_n531), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT14), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n532), .A2(new_n545), .A3(new_n533), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT14), .A4(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G107), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n546), .A2(KEYINPUT98), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n547), .A2(G107), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n532), .A2(new_n545), .A3(new_n533), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(KEYINPUT99), .B(new_n544), .C1(new_n549), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT98), .B1(new_n546), .B2(new_n548), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n550), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT99), .B1(new_n558), .B2(new_n544), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n538), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n514), .A2(new_n362), .A3(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n544), .B1(new_n549), .B2(new_n553), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n554), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n538), .A3(new_n561), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT100), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n571), .B(G902), .C1(new_n563), .C2(new_n568), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n520), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n561), .B1(new_n567), .B2(new_n538), .ZN(new_n574));
  AOI211_X1 g388(.A(new_n537), .B(new_n562), .C1(new_n566), .C2(new_n554), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n291), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n571), .ZN(new_n577));
  INV_X1    g391(.A(new_n520), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G952), .ZN(new_n581));
  AOI211_X1 g395(.A(G953), .B(new_n581), .C1(G234), .C2(G237), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n291), .B(new_n356), .C1(G234), .C2(G237), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT21), .B(G898), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(G113), .B(G122), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n379), .ZN(new_n587));
  INV_X1    g401(.A(G237), .ZN(new_n588));
  AND4_X1   g402(.A1(G143), .A2(new_n588), .A3(new_n356), .A4(G214), .ZN(new_n589));
  AOI21_X1  g403(.A(G143), .B1(new_n266), .B2(G214), .ZN(new_n590));
  OAI21_X1  g404(.A(G131), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(new_n356), .A3(G214), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n208), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n266), .A2(G143), .A3(G214), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n198), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(KEYINPUT17), .B(G131), .C1(new_n589), .C2(new_n590), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n349), .A2(new_n339), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n345), .A2(G146), .A3(new_n346), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n341), .ZN(new_n601));
  NAND2_X1  g415(.A1(KEYINPUT18), .A2(G131), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n594), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT18), .B(G131), .C1(new_n589), .C2(new_n590), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n587), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n597), .A2(new_n598), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n587), .B(new_n605), .C1(new_n350), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n599), .A2(KEYINPUT93), .A3(new_n587), .A4(new_n605), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(G475), .B1(new_n612), .B2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n611), .ZN(new_n614));
  OR3_X1    g428(.A1(new_n340), .A2(new_n336), .A3(KEYINPUT19), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT19), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n615), .B1(new_n337), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n211), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n591), .A2(new_n596), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n339), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n587), .B1(new_n620), .B2(new_n605), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT20), .ZN(new_n624));
  NOR2_X1   g438(.A1(G475), .A2(G902), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n623), .A2(KEYINPUT94), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n621), .B1(new_n610), .B2(new_n611), .ZN(new_n627));
  INV_X1    g441(.A(new_n625), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT20), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT94), .B1(new_n631), .B2(new_n624), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n613), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n580), .A2(new_n585), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n470), .A2(new_n518), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n377), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n390), .ZN(G3));
  OAI21_X1  g451(.A(G472), .B1(new_n309), .B2(G902), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n374), .A3(new_n303), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(new_n512), .A3(new_n517), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n519), .A2(new_n291), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n569), .B2(new_n519), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n574), .B2(new_n575), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n563), .A2(new_n644), .A3(new_n568), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(G478), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n633), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n445), .A2(new_n463), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n464), .ZN(new_n650));
  INV_X1    g464(.A(new_n585), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n445), .A2(new_n463), .A3(new_n465), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n378), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n640), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  NAND2_X1  g471(.A1(new_n569), .A2(KEYINPUT100), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n578), .B1(new_n577), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n570), .A2(new_n520), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n627), .A2(KEYINPUT20), .A3(new_n628), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n613), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n653), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n640), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n638), .A2(new_n303), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n359), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n354), .B(new_n670), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n371), .A2(new_n373), .B1(new_n364), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n470), .A2(new_n518), .A3(new_n634), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(new_n582), .ZN(new_n677));
  INV_X1    g491(.A(new_n583), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n677), .B1(new_n678), .B2(G900), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n613), .B(new_n679), .C1(new_n662), .C2(new_n663), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n659), .B2(new_n660), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n650), .A2(new_n378), .A3(new_n652), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n680), .B1(new_n573), .B2(new_n579), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n445), .A2(new_n463), .A3(new_n465), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n465), .B1(new_n445), .B2(new_n463), .ZN(new_n688));
  INV_X1    g502(.A(new_n378), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT101), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n672), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n518), .A2(new_n314), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XNOR2_X1  g511(.A(new_n679), .B(KEYINPUT39), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n518), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT40), .Z(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT102), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n285), .A2(new_n286), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n291), .B1(new_n703), .B2(new_n270), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n263), .A2(new_n265), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n270), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(G472), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n305), .A2(new_n311), .A3(new_n708), .A4(new_n313), .ZN(new_n709));
  INV_X1    g523(.A(new_n613), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT94), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n627), .A2(new_n711), .A3(KEYINPUT20), .A4(new_n628), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n662), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n631), .A2(new_n624), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n711), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n710), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n573), .B2(new_n579), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n378), .A3(new_n672), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT38), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n467), .B2(new_n468), .ZN(new_n720));
  INV_X1    g534(.A(new_n466), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n649), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n445), .A2(new_n463), .A3(new_n466), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(KEYINPUT38), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n701), .A2(new_n702), .A3(new_n709), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT103), .B(G143), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G45));
  NAND3_X1  g543(.A1(new_n647), .A2(new_n633), .A3(new_n679), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n683), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n694), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n211), .ZN(G48));
  AND2_X1   g548(.A1(new_n314), .A2(new_n374), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n471), .B1(new_n507), .B2(new_n291), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n510), .B2(new_n511), .ZN(new_n737));
  INV_X1    g551(.A(new_n516), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT104), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n516), .B(new_n736), .C1(new_n510), .C2(new_n511), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n735), .A2(new_n654), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n735), .A2(new_n665), .A3(new_n740), .A4(new_n743), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n739), .A2(new_n683), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n314), .A3(new_n634), .A4(new_n693), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  NOR3_X1   g565(.A1(new_n661), .A2(new_n683), .A3(new_n716), .ZN(new_n752));
  INV_X1    g566(.A(new_n374), .ZN(new_n753));
  INV_X1    g567(.A(new_n302), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n287), .A2(new_n288), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n271), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n306), .A2(new_n308), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(G472), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n301), .B2(new_n291), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n753), .A2(new_n758), .A3(new_n760), .A4(new_n585), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n740), .A2(new_n752), .A3(new_n743), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NAND2_X1  g577(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n647), .A2(new_n765), .A3(new_n633), .A4(new_n679), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n758), .A2(new_n760), .A3(new_n672), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n741), .A2(new_n768), .A3(new_n690), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(G125), .Z(G27));
  AND3_X1   g585(.A1(new_n303), .A2(KEYINPUT107), .A3(new_n304), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT107), .B1(new_n303), .B2(new_n304), .ZN(new_n773));
  OAI221_X1 g587(.A(new_n293), .B1(new_n309), .B2(new_n310), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n374), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n764), .A2(new_n766), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n722), .A2(new_n738), .A3(new_n378), .A4(new_n723), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n512), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(KEYINPUT42), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n735), .A2(new_n764), .A3(new_n766), .A4(new_n778), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n314), .A3(new_n374), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n780), .B(new_n782), .C1(new_n784), .C2(new_n767), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n779), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  NAND3_X1  g602(.A1(new_n735), .A2(new_n686), .A3(new_n778), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n489), .A2(new_n493), .A3(KEYINPUT45), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n488), .B2(new_n492), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n794), .A3(G469), .ZN(new_n795));
  NAND2_X1  g609(.A1(G469), .A2(G902), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n795), .A2(KEYINPUT108), .A3(KEYINPUT46), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n797), .A2(new_n798), .B1(new_n510), .B2(new_n511), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n516), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n698), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n722), .A2(new_n378), .A3(new_n723), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT110), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n716), .B(new_n647), .C1(KEYINPUT109), .C2(KEYINPUT43), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT109), .B(new_n613), .C1(new_n630), .C2(new_n632), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n642), .A2(new_n646), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n809), .B(new_n810), .C1(new_n633), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n669), .A3(new_n693), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n807), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  XNOR2_X1  g633(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n803), .A2(new_n821), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n314), .A2(new_n730), .A3(new_n374), .A4(new_n805), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT47), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n822), .B(new_n823), .C1(new_n803), .C2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT112), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  OAI211_X1 g642(.A(new_n744), .B(new_n747), .C1(new_n377), .C2(new_n635), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n633), .A2(new_n811), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n716), .B2(new_n661), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n470), .A2(new_n651), .A3(new_n640), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n674), .A2(new_n832), .A3(new_n750), .A4(new_n762), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n776), .A2(new_n768), .A3(new_n778), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n580), .A2(new_n805), .A3(new_n680), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n695), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n837), .A3(new_n789), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(KEYINPUT53), .A2(new_n834), .A3(new_n787), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n695), .B1(new_n692), .B2(new_n731), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n741), .A2(new_n768), .A3(new_n690), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n672), .A2(new_n738), .A3(new_n679), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n510), .A2(new_n511), .ZN(new_n845));
  INV_X1    g659(.A(new_n495), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n709), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n776), .A2(new_n842), .B1(new_n848), .B2(new_n752), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n686), .A2(KEYINPUT101), .A3(new_n690), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n694), .B1(new_n854), .B2(new_n732), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n512), .A2(new_n843), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n717), .A3(new_n709), .A4(new_n690), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n767), .B2(new_n769), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT113), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n841), .B2(new_n849), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT114), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n850), .B1(new_n841), .B2(new_n849), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n855), .A2(new_n858), .A3(KEYINPUT113), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n867));
  INV_X1    g681(.A(new_n862), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n840), .A2(new_n863), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n782), .B1(new_n784), .B2(new_n767), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT106), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n785), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n838), .B1(new_n874), .B2(new_n779), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n851), .A2(KEYINPUT52), .A3(new_n859), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n866), .A2(new_n875), .A3(new_n834), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n870), .A2(new_n871), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n877), .A2(new_n878), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n834), .A2(new_n787), .A3(new_n839), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n869), .A2(new_n863), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n883), .B2(KEYINPUT53), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n884), .B2(KEYINPUT54), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT50), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n813), .B2(new_n582), .ZN(new_n888));
  AOI211_X1 g702(.A(KEYINPUT115), .B(new_n677), .C1(new_n808), .C2(new_n812), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n725), .A2(new_n741), .A3(new_n689), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n753), .A2(new_n758), .A3(new_n760), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n725), .A2(new_n741), .A3(KEYINPUT116), .A4(new_n689), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n886), .B1(new_n890), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n813), .A2(new_n582), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n813), .A2(new_n887), .A3(new_n582), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n895), .A2(new_n894), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n378), .B1(new_n720), .B2(new_n724), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT116), .B1(new_n905), .B2(new_n741), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT50), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT118), .A4(KEYINPUT50), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT117), .B(new_n886), .C1(new_n890), .C2(new_n896), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n899), .A2(new_n910), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n739), .A2(new_n805), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n768), .B(new_n914), .C1(new_n888), .C2(new_n889), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n709), .A2(new_n753), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n914), .A2(new_n916), .A3(new_n582), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n716), .A3(new_n811), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n822), .B1(new_n803), .B2(new_n825), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n737), .A2(new_n517), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n806), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n903), .A2(new_n894), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n913), .A2(KEYINPUT51), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n903), .A2(new_n775), .A3(new_n914), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT48), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n749), .ZN(new_n929));
  INV_X1    g743(.A(new_n648), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n581), .B(G953), .C1(new_n917), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n913), .A2(new_n924), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT51), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT119), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n938), .B(KEYINPUT51), .C1(new_n913), .C2(new_n924), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n934), .B(KEYINPUT120), .C1(new_n937), .C2(new_n939), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n885), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n885), .A2(new_n942), .A3(new_n946), .A4(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n581), .A2(new_n356), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n737), .B(KEYINPUT49), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n517), .B(new_n689), .C1(new_n720), .C2(new_n724), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n633), .A2(new_n811), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .A4(new_n916), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n949), .A2(new_n953), .ZN(G75));
  NOR2_X1   g768(.A1(new_n356), .A2(G952), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n291), .B1(new_n870), .B2(new_n879), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT56), .B1(new_n957), .B2(G210), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n417), .A2(new_n439), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n444), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT55), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n956), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n957), .A2(new_n963), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n465), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT56), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n967), .B2(new_n969), .ZN(G51));
  AOI21_X1  g784(.A(new_n871), .B1(new_n870), .B2(new_n879), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n880), .A2(new_n971), .A3(KEYINPUT123), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n880), .B2(KEYINPUT123), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n796), .B(KEYINPUT57), .Z(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n507), .ZN(new_n976));
  INV_X1    g790(.A(new_n795), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n966), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n955), .B1(new_n976), .B2(new_n978), .ZN(G54));
  AND2_X1   g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n623), .B1(new_n966), .B2(new_n980), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n623), .A2(new_n964), .A3(new_n965), .A4(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n955), .ZN(G60));
  NAND2_X1  g797(.A1(new_n643), .A2(new_n645), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n641), .B(KEYINPUT59), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n972), .A2(new_n973), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n985), .B1(new_n885), .B2(new_n986), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n988), .A2(new_n956), .A3(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n870), .B2(new_n879), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n671), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT124), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n360), .A2(new_n361), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT125), .Z(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT124), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n993), .A2(new_n1000), .A3(new_n671), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n995), .A2(new_n999), .A3(new_n956), .A4(new_n1001), .ZN(new_n1002));
  OR2_X1    g816(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n1003));
  NAND2_X1  g817(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(G66));
  OAI21_X1  g821(.A(G953), .B1(new_n584), .B2(new_n442), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n834), .B2(G953), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n959), .B1(G898), .B2(new_n356), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  NAND2_X1  g825(.A1(new_n236), .A2(new_n244), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(new_n617), .ZN(new_n1013));
  NAND3_X1  g827(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n855), .A2(new_n770), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n727), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1018));
  INV_X1    g832(.A(new_n818), .ZN(new_n1019));
  INV_X1    g833(.A(new_n377), .ZN(new_n1020));
  INV_X1    g834(.A(new_n831), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n1021), .A2(new_n699), .A3(new_n805), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1019), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1017), .A2(new_n827), .A3(new_n1018), .A4(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1013), .B(new_n1014), .C1(new_n1024), .C2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n818), .A2(new_n1015), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT127), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n775), .A2(new_n698), .A3(new_n752), .A4(new_n803), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n827), .A2(new_n789), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1027), .A2(new_n1029), .A3(new_n787), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1030), .A2(new_n356), .ZN(new_n1031));
  INV_X1    g845(.A(G900), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n1032), .A2(new_n356), .A3(G227), .ZN(new_n1033));
  OR2_X1    g847(.A1(new_n1013), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1025), .B1(new_n1031), .B2(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  INV_X1    g851(.A(new_n834), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1037), .B1(new_n1024), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n707), .ZN(new_n1040));
  INV_X1    g854(.A(new_n272), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n884), .A2(new_n1041), .A3(new_n706), .A4(new_n1037), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1037), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n955), .B1(new_n1043), .B2(new_n272), .ZN(new_n1044));
  AND3_X1   g858(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(G57));
endmodule


