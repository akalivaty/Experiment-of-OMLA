

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761;

  XNOR2_X1 U364 ( .A(n597), .B(KEYINPUT1), .ZN(n570) );
  INV_X1 U365 ( .A(G146), .ZN(n436) );
  BUF_X1 U366 ( .A(G119), .Z(n431) );
  XNOR2_X2 U367 ( .A(n372), .B(n710), .ZN(n712) );
  AND2_X2 U368 ( .A1(n441), .A2(n443), .ZN(n356) );
  NAND2_X2 U369 ( .A1(n418), .A2(n580), .ZN(n417) );
  XNOR2_X2 U370 ( .A(n523), .B(n487), .ZN(n748) );
  XNOR2_X2 U371 ( .A(n748), .B(n478), .ZN(n715) );
  NAND2_X1 U372 ( .A1(n570), .A2(n592), .ZN(n343) );
  AND2_X2 U373 ( .A1(n346), .A2(KEYINPUT2), .ZN(n411) );
  XNOR2_X2 U374 ( .A(n389), .B(KEYINPUT45), .ZN(n346) );
  XNOR2_X2 U375 ( .A(n416), .B(n474), .ZN(n523) );
  XNOR2_X2 U376 ( .A(n417), .B(n358), .ZN(n757) );
  NOR2_X2 U377 ( .A1(n613), .A2(n700), .ZN(n602) );
  XNOR2_X2 U378 ( .A(n426), .B(n601), .ZN(n700) );
  XNOR2_X2 U379 ( .A(n345), .B(n354), .ZN(n420) );
  INV_X2 U380 ( .A(G953), .ZN(n452) );
  NOR2_X1 U381 ( .A1(n699), .A2(n577), .ZN(n419) );
  NOR2_X1 U382 ( .A1(n574), .A2(n606), .ZN(n576) );
  XNOR2_X1 U383 ( .A(n555), .B(KEYINPUT100), .ZN(n605) );
  XNOR2_X1 U384 ( .A(n567), .B(n357), .ZN(n606) );
  INV_X1 U385 ( .A(n749), .ZN(n451) );
  NOR2_X1 U386 ( .A1(n649), .A2(KEYINPUT83), .ZN(n393) );
  XNOR2_X1 U387 ( .A(n419), .B(KEYINPUT34), .ZN(n418) );
  NOR2_X1 U388 ( .A1(n368), .A2(n382), .ZN(n381) );
  BUF_X1 U389 ( .A(n699), .Z(n344) );
  XNOR2_X1 U390 ( .A(n576), .B(n575), .ZN(n699) );
  AND2_X1 U391 ( .A1(n374), .A2(n386), .ZN(n363) );
  INV_X1 U392 ( .A(n453), .ZN(n378) );
  NAND2_X1 U393 ( .A1(n453), .A2(n455), .ZN(n387) );
  XNOR2_X1 U394 ( .A(n599), .B(KEYINPUT109), .ZN(n672) );
  XNOR2_X1 U395 ( .A(n348), .B(n427), .ZN(n668) );
  OR2_X1 U396 ( .A1(n729), .A2(G902), .ZN(n402) );
  XNOR2_X1 U397 ( .A(n609), .B(KEYINPUT111), .ZN(n610) );
  XNOR2_X1 U398 ( .A(G137), .B(G140), .ZN(n487) );
  XNOR2_X2 U399 ( .A(G146), .B(G125), .ZN(n500) );
  XOR2_X1 U400 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n486) );
  AND2_X1 U401 ( .A1(n397), .A2(n396), .ZN(n395) );
  OR2_X1 U402 ( .A1(n632), .A2(n345), .ZN(n410) );
  NAND2_X1 U403 ( .A1(n589), .A2(n667), .ZN(n345) );
  AND2_X1 U404 ( .A1(n346), .A2(n447), .ZN(n355) );
  BUF_X1 U405 ( .A(n389), .Z(n347) );
  XNOR2_X1 U406 ( .A(n507), .B(n506), .ZN(n348) );
  NOR2_X2 U407 ( .A1(n711), .A2(n505), .ZN(n507) );
  XNOR2_X1 U408 ( .A(n347), .B(KEYINPUT45), .ZN(n349) );
  XNOR2_X2 U409 ( .A(G119), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X2 U410 ( .A(n449), .B(n448), .ZN(n415) );
  XNOR2_X1 U411 ( .A(G902), .B(KEYINPUT15), .ZN(n640) );
  XNOR2_X1 U412 ( .A(n561), .B(KEYINPUT22), .ZN(n562) );
  INV_X1 U413 ( .A(KEYINPUT0), .ZN(n514) );
  NAND2_X1 U414 ( .A1(n649), .A2(KEYINPUT83), .ZN(n396) );
  XOR2_X1 U415 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n539) );
  XOR2_X1 U416 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n501) );
  NOR2_X1 U417 ( .A1(n640), .A2(n450), .ZN(n447) );
  NAND2_X1 U418 ( .A1(n505), .A2(n446), .ZN(n445) );
  NAND2_X1 U419 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n446) );
  NOR2_X1 U420 ( .A1(n513), .A2(n351), .ZN(n455) );
  NOR2_X1 U421 ( .A1(G953), .A2(G237), .ZN(n540) );
  XOR2_X1 U422 ( .A(KEYINPUT67), .B(G101), .Z(n515) );
  INV_X1 U423 ( .A(n562), .ZN(n386) );
  XNOR2_X1 U424 ( .A(n498), .B(n353), .ZN(n471) );
  XNOR2_X1 U425 ( .A(G134), .B(G131), .ZN(n474) );
  AND2_X1 U426 ( .A1(n463), .A2(n761), .ZN(n462) );
  XOR2_X1 U427 ( .A(KEYINPUT24), .B(G110), .Z(n493) );
  XNOR2_X1 U428 ( .A(n431), .B(G128), .ZN(n492) );
  XNOR2_X1 U429 ( .A(n409), .B(n590), .ZN(n638) );
  INV_X1 U430 ( .A(KEYINPUT39), .ZN(n590) );
  NOR2_X1 U431 ( .A1(n588), .A2(n408), .ZN(n407) );
  NAND2_X1 U432 ( .A1(n381), .A2(n380), .ZN(n379) );
  NOR2_X1 U433 ( .A1(n625), .A2(n653), .ZN(n626) );
  XOR2_X1 U434 ( .A(n556), .B(KEYINPUT101), .Z(n671) );
  INV_X1 U435 ( .A(KEYINPUT38), .ZN(n427) );
  OR2_X1 U436 ( .A1(G237), .A2(G902), .ZN(n508) );
  INV_X1 U437 ( .A(KEYINPUT44), .ZN(n421) );
  XOR2_X1 U438 ( .A(G122), .B(G104), .Z(n544) );
  XNOR2_X1 U439 ( .A(G113), .B(G143), .ZN(n543) );
  XNOR2_X1 U440 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n538) );
  XNOR2_X1 U441 ( .A(G131), .B(G140), .ZN(n545) );
  XOR2_X1 U442 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n546) );
  XNOR2_X1 U443 ( .A(n425), .B(n457), .ZN(n424) );
  XNOR2_X1 U444 ( .A(n500), .B(KEYINPUT18), .ZN(n457) );
  XNOR2_X1 U445 ( .A(n503), .B(n501), .ZN(n425) );
  XNOR2_X1 U446 ( .A(n735), .B(n515), .ZN(n502) );
  NAND2_X1 U447 ( .A1(n445), .A2(n444), .ZN(n443) );
  NAND2_X1 U448 ( .A1(n640), .A2(KEYINPUT66), .ZN(n444) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n509) );
  NOR2_X1 U450 ( .A1(n455), .A2(n377), .ZN(n376) );
  NAND2_X1 U451 ( .A1(n570), .A2(n685), .ZN(n574) );
  XNOR2_X1 U452 ( .A(n414), .B(n440), .ZN(n518) );
  XNOR2_X1 U453 ( .A(G116), .B(G113), .ZN(n440) );
  XNOR2_X1 U454 ( .A(n413), .B(KEYINPUT71), .ZN(n414) );
  XNOR2_X1 U455 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n520) );
  XOR2_X1 U456 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n521) );
  XNOR2_X1 U457 ( .A(n517), .B(n435), .ZN(n519) );
  XNOR2_X1 U458 ( .A(n516), .B(n436), .ZN(n435) );
  XNOR2_X1 U459 ( .A(n518), .B(n504), .ZN(n732) );
  XNOR2_X1 U460 ( .A(KEYINPUT16), .B(G122), .ZN(n504) );
  INV_X1 U461 ( .A(G143), .ZN(n428) );
  XOR2_X1 U462 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n533) );
  XOR2_X1 U463 ( .A(G122), .B(G107), .Z(n530) );
  XNOR2_X1 U464 ( .A(G116), .B(G134), .ZN(n529) );
  INV_X1 U465 ( .A(KEYINPUT73), .ZN(n448) );
  XNOR2_X1 U466 ( .A(n554), .B(n553), .ZN(n558) );
  XNOR2_X1 U467 ( .A(n475), .B(n458), .ZN(n735) );
  INV_X1 U468 ( .A(G107), .ZN(n458) );
  XNOR2_X1 U469 ( .A(G104), .B(G110), .ZN(n475) );
  XNOR2_X1 U470 ( .A(n403), .B(n496), .ZN(n729) );
  XNOR2_X1 U471 ( .A(KEYINPUT81), .B(KEYINPUT23), .ZN(n494) );
  AND2_X1 U472 ( .A1(n473), .A2(G475), .ZN(n469) );
  NOR2_X1 U473 ( .A1(n638), .A2(n605), .ZN(n591) );
  AND2_X1 U474 ( .A1(n569), .A2(n430), .ZN(n649) );
  NAND2_X1 U475 ( .A1(n460), .A2(n723), .ZN(n459) );
  XNOR2_X1 U476 ( .A(n461), .B(n359), .ZN(n460) );
  INV_X1 U477 ( .A(KEYINPUT124), .ZN(n437) );
  NAND2_X1 U478 ( .A1(n439), .A2(n723), .ZN(n438) );
  XNOR2_X1 U479 ( .A(n719), .B(n718), .ZN(n439) );
  NAND2_X1 U480 ( .A1(n412), .A2(n362), .ZN(n350) );
  XOR2_X1 U481 ( .A(n514), .B(KEYINPUT84), .Z(n351) );
  INV_X1 U482 ( .A(G953), .ZN(n484) );
  AND2_X1 U483 ( .A1(n566), .A2(n643), .ZN(n352) );
  XNOR2_X1 U484 ( .A(KEYINPUT25), .B(KEYINPUT88), .ZN(n353) );
  XOR2_X1 U485 ( .A(KEYINPUT74), .B(KEYINPUT19), .Z(n354) );
  INV_X1 U486 ( .A(n593), .ZN(n465) );
  XOR2_X1 U487 ( .A(KEYINPUT6), .B(KEYINPUT102), .Z(n357) );
  XOR2_X1 U488 ( .A(KEYINPUT35), .B(KEYINPUT75), .Z(n358) );
  XOR2_X1 U489 ( .A(n642), .B(KEYINPUT62), .Z(n359) );
  INV_X1 U490 ( .A(KEYINPUT66), .ZN(n450) );
  XNOR2_X1 U491 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n360) );
  AND2_X1 U492 ( .A1(n467), .A2(n723), .ZN(n361) );
  AND2_X1 U493 ( .A1(n450), .A2(n442), .ZN(n362) );
  NOR2_X1 U494 ( .A1(G952), .A2(n452), .ZN(n731) );
  INV_X1 U495 ( .A(n731), .ZN(n723) );
  INV_X1 U496 ( .A(KEYINPUT2), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n559), .B(KEYINPUT103), .ZN(n560) );
  INV_X1 U498 ( .A(n560), .ZN(n380) );
  BUF_X1 U499 ( .A(n749), .Z(n364) );
  BUF_X1 U500 ( .A(n518), .Z(n365) );
  XNOR2_X2 U501 ( .A(n366), .B(G472), .ZN(n567) );
  NOR2_X1 U502 ( .A1(n642), .A2(G902), .ZN(n366) );
  NAND2_X1 U503 ( .A1(n668), .A2(n593), .ZN(n408) );
  NAND2_X1 U504 ( .A1(n420), .A2(n351), .ZN(n367) );
  NAND2_X1 U505 ( .A1(n420), .A2(n351), .ZN(n454) );
  NAND2_X1 U506 ( .A1(n367), .A2(n456), .ZN(n368) );
  BUF_X1 U507 ( .A(n748), .Z(n369) );
  BUF_X1 U508 ( .A(n597), .Z(n370) );
  NAND2_X1 U509 ( .A1(n383), .A2(n379), .ZN(n371) );
  NAND2_X1 U510 ( .A1(n383), .A2(n379), .ZN(n573) );
  XNOR2_X1 U511 ( .A(n732), .B(n424), .ZN(n423) );
  BUF_X1 U512 ( .A(n711), .Z(n372) );
  XNOR2_X1 U513 ( .A(n423), .B(n422), .ZN(n711) );
  BUF_X1 U514 ( .A(n415), .Z(n373) );
  NAND2_X1 U515 ( .A1(n363), .A2(n375), .ZN(n384) );
  NAND2_X1 U516 ( .A1(n367), .A2(n376), .ZN(n374) );
  NAND2_X1 U517 ( .A1(n378), .A2(n388), .ZN(n375) );
  AND2_X2 U518 ( .A1(n454), .A2(n456), .ZN(n388) );
  NAND2_X1 U519 ( .A1(n388), .A2(n387), .ZN(n577) );
  INV_X1 U520 ( .A(n456), .ZN(n377) );
  NAND2_X1 U521 ( .A1(n387), .A2(n562), .ZN(n382) );
  AND2_X2 U522 ( .A1(n384), .A2(n385), .ZN(n383) );
  NAND2_X1 U523 ( .A1(n560), .A2(n386), .ZN(n385) );
  NAND2_X2 U524 ( .A1(n390), .A2(n352), .ZN(n389) );
  XNOR2_X2 U525 ( .A(n391), .B(n421), .ZN(n390) );
  NAND2_X1 U526 ( .A1(n398), .A2(n399), .ZN(n391) );
  NAND2_X1 U527 ( .A1(n393), .A2(n392), .ZN(n394) );
  INV_X1 U528 ( .A(n758), .ZN(n392) );
  NAND2_X1 U529 ( .A1(n395), .A2(n394), .ZN(n398) );
  NAND2_X1 U530 ( .A1(n758), .A2(KEYINPUT83), .ZN(n397) );
  INV_X1 U531 ( .A(n757), .ZN(n399) );
  NAND2_X1 U532 ( .A1(n356), .A2(n350), .ZN(n433) );
  XNOR2_X2 U533 ( .A(n400), .B(G478), .ZN(n578) );
  NOR2_X2 U534 ( .A1(n726), .A2(G902), .ZN(n400) );
  XNOR2_X2 U535 ( .A(n401), .B(KEYINPUT32), .ZN(n758) );
  NOR2_X2 U536 ( .A1(n573), .A2(n572), .ZN(n401) );
  XNOR2_X2 U537 ( .A(n402), .B(n471), .ZN(n592) );
  XNOR2_X1 U538 ( .A(n491), .B(n404), .ZN(n403) );
  INV_X1 U539 ( .A(n747), .ZN(n404) );
  AND2_X1 U540 ( .A1(n405), .A2(n406), .ZN(n622) );
  NOR2_X1 U541 ( .A1(n588), .A2(n465), .ZN(n405) );
  NAND2_X1 U542 ( .A1(n407), .A2(n406), .ZN(n409) );
  XNOR2_X1 U543 ( .A(n581), .B(KEYINPUT107), .ZN(n406) );
  NAND2_X1 U544 ( .A1(n349), .A2(n451), .ZN(n412) );
  AND2_X1 U545 ( .A1(n349), .A2(n452), .ZN(n743) );
  INV_X1 U546 ( .A(n410), .ZN(n611) );
  NAND2_X1 U547 ( .A1(n355), .A2(n451), .ZN(n441) );
  NAND2_X1 U548 ( .A1(n411), .A2(n451), .ZN(n449) );
  AND2_X1 U549 ( .A1(n412), .A2(n442), .ZN(n703) );
  NAND2_X1 U550 ( .A1(n415), .A2(n433), .ZN(n641) );
  NAND2_X1 U551 ( .A1(n704), .A2(n373), .ZN(n705) );
  XNOR2_X1 U552 ( .A(n502), .B(n416), .ZN(n422) );
  XNOR2_X2 U553 ( .A(n536), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X2 U554 ( .A(n480), .B(n479), .ZN(n597) );
  INV_X1 U555 ( .A(n420), .ZN(n453) );
  NOR2_X1 U556 ( .A1(n613), .A2(n378), .ZN(n618) );
  NOR2_X2 U557 ( .A1(n592), .A2(n678), .ZN(n685) );
  NAND2_X1 U558 ( .A1(n672), .A2(n600), .ZN(n426) );
  XNOR2_X2 U559 ( .A(n429), .B(n428), .ZN(n536) );
  XNOR2_X2 U560 ( .A(G128), .B(KEYINPUT77), .ZN(n429) );
  NOR2_X1 U561 ( .A1(n568), .A2(n682), .ZN(n430) );
  NOR2_X2 U562 ( .A1(n715), .A2(G902), .ZN(n480) );
  NOR2_X1 U563 ( .A1(n371), .A2(n684), .ZN(n569) );
  XNOR2_X1 U564 ( .A(n432), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U565 ( .A1(n466), .A2(n470), .ZN(n432) );
  XNOR2_X1 U566 ( .A(n438), .B(n437), .ZN(G54) );
  XNOR2_X1 U567 ( .A(n434), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U568 ( .A1(n714), .A2(n731), .ZN(n434) );
  NAND2_X1 U569 ( .A1(n464), .A2(n462), .ZN(n749) );
  INV_X1 U570 ( .A(n665), .ZN(n463) );
  NOR2_X1 U571 ( .A1(n760), .A2(n759), .ZN(n604) );
  NAND2_X1 U572 ( .A1(n513), .A2(n351), .ZN(n456) );
  XNOR2_X1 U573 ( .A(n459), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U574 ( .A1(n720), .A2(G472), .ZN(n461) );
  XNOR2_X1 U575 ( .A(n631), .B(n360), .ZN(n464) );
  NAND2_X1 U576 ( .A1(n724), .A2(n469), .ZN(n468) );
  NAND2_X1 U577 ( .A1(n468), .A2(n361), .ZN(n466) );
  OR2_X1 U578 ( .A1(n473), .A2(G475), .ZN(n467) );
  NOR2_X1 U579 ( .A1(n724), .A2(n473), .ZN(n470) );
  AND2_X1 U580 ( .A1(G214), .A2(n540), .ZN(n472) );
  XOR2_X1 U581 ( .A(n722), .B(n721), .Z(n473) );
  XNOR2_X1 U582 ( .A(n476), .B(n436), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n502), .B(n477), .ZN(n478) );
  XNOR2_X1 U584 ( .A(n541), .B(n472), .ZN(n542) );
  XNOR2_X1 U585 ( .A(n747), .B(n542), .ZN(n550) );
  INV_X1 U586 ( .A(KEYINPUT36), .ZN(n609) );
  INV_X1 U587 ( .A(n558), .ZN(n579) );
  XNOR2_X1 U588 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n611), .B(n610), .ZN(n612) );
  XOR2_X1 U590 ( .A(KEYINPUT105), .B(n605), .Z(n657) );
  AND2_X1 U591 ( .A1(G227), .A2(n452), .ZN(n476) );
  XOR2_X1 U592 ( .A(KEYINPUT70), .B(G469), .Z(n479) );
  XOR2_X1 U593 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n483) );
  NAND2_X1 U594 ( .A1(G234), .A2(n640), .ZN(n481) );
  XNOR2_X1 U595 ( .A(KEYINPUT20), .B(n481), .ZN(n497) );
  NAND2_X1 U596 ( .A1(G221), .A2(n497), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n483), .B(n482), .ZN(n678) );
  NAND2_X1 U598 ( .A1(G234), .A2(n484), .ZN(n485) );
  XNOR2_X1 U599 ( .A(n486), .B(n485), .ZN(n531) );
  NAND2_X1 U600 ( .A1(n531), .A2(G221), .ZN(n489) );
  XNOR2_X1 U601 ( .A(n487), .B(KEYINPUT87), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n489), .B(n488), .ZN(n491) );
  INV_X1 U603 ( .A(n500), .ZN(n490) );
  XOR2_X1 U604 ( .A(KEYINPUT10), .B(n490), .Z(n747) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n495) );
  NAND2_X1 U606 ( .A1(n497), .A2(G217), .ZN(n498) );
  NAND2_X1 U607 ( .A1(n370), .A2(n685), .ZN(n499) );
  XNOR2_X2 U608 ( .A(n499), .B(KEYINPUT90), .ZN(n581) );
  NAND2_X1 U609 ( .A1(G224), .A2(n452), .ZN(n503) );
  INV_X1 U610 ( .A(n640), .ZN(n505) );
  NAND2_X1 U611 ( .A1(G210), .A2(n508), .ZN(n506) );
  XNOR2_X1 U612 ( .A(n507), .B(n506), .ZN(n589) );
  NAND2_X1 U613 ( .A1(G214), .A2(n508), .ZN(n667) );
  XNOR2_X1 U614 ( .A(n509), .B(KEYINPUT14), .ZN(n510) );
  NAND2_X1 U615 ( .A1(G952), .A2(n510), .ZN(n698) );
  NOR2_X1 U616 ( .A1(G953), .A2(n698), .ZN(n585) );
  NAND2_X1 U617 ( .A1(G902), .A2(n510), .ZN(n582) );
  INV_X1 U618 ( .A(G898), .ZN(n741) );
  NAND2_X1 U619 ( .A1(G953), .A2(n741), .ZN(n737) );
  NOR2_X1 U620 ( .A1(n582), .A2(n737), .ZN(n511) );
  NOR2_X1 U621 ( .A1(n585), .A2(n511), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n512), .B(KEYINPUT86), .ZN(n513) );
  NOR2_X1 U623 ( .A1(n581), .A2(n577), .ZN(n526) );
  XOR2_X1 U624 ( .A(n515), .B(G137), .Z(n517) );
  NAND2_X1 U625 ( .A1(n540), .A2(G210), .ZN(n516) );
  XNOR2_X1 U626 ( .A(n365), .B(n519), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U628 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U629 ( .A(n525), .B(n524), .ZN(n642) );
  NAND2_X1 U630 ( .A1(n526), .A2(n567), .ZN(n645) );
  NOR2_X1 U631 ( .A1(n567), .A2(n574), .ZN(n690) );
  INV_X1 U632 ( .A(n577), .ZN(n527) );
  NAND2_X1 U633 ( .A1(n690), .A2(n527), .ZN(n528) );
  XOR2_X1 U634 ( .A(KEYINPUT31), .B(n528), .Z(n659) );
  NAND2_X1 U635 ( .A1(n645), .A2(n659), .ZN(n557) );
  XNOR2_X1 U636 ( .A(n530), .B(n529), .ZN(n535) );
  NAND2_X1 U637 ( .A1(G217), .A2(n531), .ZN(n532) );
  XNOR2_X1 U638 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U639 ( .A(n535), .B(n534), .ZN(n537) );
  XNOR2_X1 U640 ( .A(n536), .B(n537), .ZN(n726) );
  XNOR2_X1 U641 ( .A(n539), .B(n538), .ZN(n541) );
  XNOR2_X1 U642 ( .A(n544), .B(n543), .ZN(n548) );
  XNOR2_X1 U643 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U644 ( .A(n548), .B(n547), .Z(n549) );
  XNOR2_X1 U645 ( .A(n550), .B(n549), .ZN(n722) );
  NOR2_X1 U646 ( .A1(n722), .A2(G902), .ZN(n554) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(KEYINPUT98), .Z(n552) );
  XNOR2_X1 U648 ( .A(KEYINPUT99), .B(G475), .ZN(n551) );
  XNOR2_X1 U649 ( .A(n552), .B(n551), .ZN(n553) );
  OR2_X1 U650 ( .A1(n578), .A2(n558), .ZN(n660) );
  NAND2_X1 U651 ( .A1(n558), .A2(n578), .ZN(n555) );
  NAND2_X1 U652 ( .A1(n660), .A2(n605), .ZN(n556) );
  NAND2_X1 U653 ( .A1(n557), .A2(n671), .ZN(n566) );
  INV_X1 U654 ( .A(n592), .ZN(n568) );
  BUF_X1 U655 ( .A(n570), .Z(n684) );
  INV_X1 U656 ( .A(n606), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n578), .A2(n579), .ZN(n670) );
  NOR2_X1 U658 ( .A1(n678), .A2(n670), .ZN(n559) );
  INV_X1 U659 ( .A(KEYINPUT72), .ZN(n561) );
  NOR2_X1 U660 ( .A1(n571), .A2(n371), .ZN(n563) );
  XOR2_X1 U661 ( .A(KEYINPUT82), .B(n563), .Z(n564) );
  NOR2_X1 U662 ( .A1(n684), .A2(n564), .ZN(n565) );
  NAND2_X1 U663 ( .A1(n568), .A2(n565), .ZN(n643) );
  INV_X1 U664 ( .A(n567), .ZN(n682) );
  OR2_X1 U665 ( .A1(n571), .A2(n343), .ZN(n572) );
  XNOR2_X1 U666 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n575) );
  NOR2_X1 U667 ( .A1(n579), .A2(n578), .ZN(n621) );
  XNOR2_X1 U668 ( .A(n621), .B(KEYINPUT76), .ZN(n580) );
  OR2_X1 U669 ( .A1(n452), .A2(n582), .ZN(n583) );
  NOR2_X1 U670 ( .A1(G900), .A2(n583), .ZN(n584) );
  NOR2_X1 U671 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U672 ( .A(KEYINPUT78), .B(n586), .Z(n593) );
  NAND2_X1 U673 ( .A1(n682), .A2(n667), .ZN(n587) );
  XNOR2_X1 U674 ( .A(KEYINPUT30), .B(n587), .ZN(n588) );
  XNOR2_X1 U675 ( .A(n591), .B(KEYINPUT40), .ZN(n760) );
  XOR2_X1 U676 ( .A(KEYINPUT108), .B(KEYINPUT28), .Z(n596) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U678 ( .A1(n678), .A2(n594), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n608), .A2(n682), .ZN(n595) );
  XNOR2_X1 U680 ( .A(n596), .B(n595), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n598), .A2(n370), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n601) );
  INV_X1 U683 ( .A(n670), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n667), .A2(n668), .ZN(n599) );
  XNOR2_X1 U685 ( .A(n602), .B(KEYINPUT42), .ZN(n759) );
  XNOR2_X1 U686 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n603) );
  XNOR2_X1 U687 ( .A(n604), .B(n603), .ZN(n630) );
  NOR2_X1 U688 ( .A1(n606), .A2(n657), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n632) );
  NAND2_X1 U690 ( .A1(n612), .A2(n684), .ZN(n664) );
  INV_X1 U691 ( .A(n671), .ZN(n616) );
  NOR2_X1 U692 ( .A1(KEYINPUT47), .A2(n616), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n618), .A2(n614), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n664), .A2(n615), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n616), .A2(KEYINPUT47), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n617), .B(KEYINPUT80), .ZN(n620) );
  INV_X1 U697 ( .A(n618), .ZN(n654) );
  NAND2_X1 U698 ( .A1(n654), .A2(KEYINPUT47), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n625) );
  INV_X1 U700 ( .A(n348), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n653) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n626), .ZN(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U706 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n636) );
  INV_X1 U707 ( .A(n632), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n633), .A2(n667), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n634), .A2(n684), .ZN(n635) );
  XOR2_X1 U710 ( .A(n636), .B(n635), .Z(n637) );
  NOR2_X1 U711 ( .A1(n348), .A2(n637), .ZN(n665) );
  OR2_X1 U712 ( .A1(n660), .A2(n638), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n639), .B(KEYINPUT112), .ZN(n761) );
  XNOR2_X2 U714 ( .A(n641), .B(KEYINPUT65), .ZN(n720) );
  XNOR2_X1 U715 ( .A(G101), .B(n643), .ZN(G3) );
  NOR2_X1 U716 ( .A1(n657), .A2(n645), .ZN(n644) );
  XOR2_X1 U717 ( .A(G104), .B(n644), .Z(G6) );
  NOR2_X1 U718 ( .A1(n660), .A2(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U721 ( .A(G107), .B(n648), .ZN(G9) );
  XOR2_X1 U722 ( .A(n649), .B(G110), .Z(G12) );
  XOR2_X1 U723 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n651) );
  OR2_X1 U724 ( .A1(n654), .A2(n660), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U726 ( .A(G128), .B(n652), .Z(G30) );
  XOR2_X1 U727 ( .A(G143), .B(n653), .Z(G45) );
  NOR2_X1 U728 ( .A1(n657), .A2(n654), .ZN(n655) );
  XOR2_X1 U729 ( .A(KEYINPUT114), .B(n655), .Z(n656) );
  XNOR2_X1 U730 ( .A(G146), .B(n656), .ZN(G48) );
  NOR2_X1 U731 ( .A1(n657), .A2(n659), .ZN(n658) );
  XOR2_X1 U732 ( .A(G113), .B(n658), .Z(G15) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n662) );
  XNOR2_X1 U734 ( .A(G116), .B(KEYINPUT115), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(G18) );
  XOR2_X1 U736 ( .A(G125), .B(KEYINPUT37), .Z(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(G27) );
  XOR2_X1 U738 ( .A(G140), .B(n665), .Z(n666) );
  XNOR2_X1 U739 ( .A(KEYINPUT116), .B(n666), .ZN(G42) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U743 ( .A(KEYINPUT120), .B(n673), .Z(n674) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U745 ( .A(KEYINPUT121), .B(n676), .Z(n677) );
  NOR2_X1 U746 ( .A1(n344), .A2(n677), .ZN(n695) );
  XNOR2_X1 U747 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n692) );
  XOR2_X1 U748 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n680) );
  NAND2_X1 U749 ( .A1(n678), .A2(n592), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U752 ( .A(KEYINPUT118), .B(n683), .Z(n688) );
  NOR2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U754 ( .A(KEYINPUT50), .B(n686), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n700), .A2(n693), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U760 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n700), .A2(n344), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n706) );
  INV_X1 U764 ( .A(n703), .ZN(n704) );
  NAND2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(KEYINPUT122), .B(n707), .ZN(n708) );
  NOR2_X1 U767 ( .A1(n708), .A2(G953), .ZN(n709) );
  XNOR2_X1 U768 ( .A(n709), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U769 ( .A1(n720), .A2(G210), .ZN(n713) );
  XOR2_X1 U770 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n710) );
  XNOR2_X1 U771 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U772 ( .A1(n720), .A2(G469), .ZN(n719) );
  XOR2_X1 U773 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  XNOR2_X1 U774 ( .A(n715), .B(KEYINPUT123), .ZN(n716) );
  XNOR2_X1 U775 ( .A(n717), .B(n716), .ZN(n718) );
  BUF_X2 U776 ( .A(n720), .Z(n724) );
  INV_X1 U777 ( .A(KEYINPUT59), .ZN(n721) );
  NAND2_X1 U778 ( .A1(G478), .A2(n724), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n731), .A2(n727), .ZN(G63) );
  NAND2_X1 U781 ( .A1(G217), .A2(n724), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(G66) );
  BUF_X1 U784 ( .A(n732), .Z(n733) );
  XOR2_X1 U785 ( .A(G101), .B(n733), .Z(n734) );
  XNOR2_X1 U786 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n746) );
  NAND2_X1 U788 ( .A1(G224), .A2(G953), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n738), .B(KEYINPUT61), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n739), .B(KEYINPUT125), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n742), .B(KEYINPUT126), .ZN(n744) );
  NOR2_X1 U793 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(G69) );
  XOR2_X1 U795 ( .A(n369), .B(n747), .Z(n751) );
  XNOR2_X1 U796 ( .A(n364), .B(n751), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n750), .A2(n452), .ZN(n756) );
  XNOR2_X1 U798 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(G953), .ZN(n754) );
  XOR2_X1 U801 ( .A(KEYINPUT127), .B(n754), .Z(n755) );
  NAND2_X1 U802 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U803 ( .A(n757), .B(G122), .Z(G24) );
  XOR2_X1 U804 ( .A(n758), .B(n431), .Z(G21) );
  XOR2_X1 U805 ( .A(n759), .B(G137), .Z(G39) );
  XOR2_X1 U806 ( .A(n760), .B(G131), .Z(G33) );
  XNOR2_X1 U807 ( .A(G134), .B(n761), .ZN(G36) );
endmodule

