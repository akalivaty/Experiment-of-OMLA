//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(KEYINPUT24), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n204), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT24), .A3(new_n203), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(KEYINPUT25), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n204), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n205), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT27), .B1(new_n211), .B2(KEYINPUT65), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT27), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(G183gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n225), .A3(new_n212), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT27), .B(G183gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n227), .A2(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT26), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n203), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n202), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(new_n233), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G120gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G113gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n246));
  INV_X1    g045(.A(G134gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G127gat), .ZN(new_n248));
  INV_X1    g047(.A(G127gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G134gat), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n245), .A2(new_n246), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n250), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n221), .A2(new_n240), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n221), .B2(new_n240), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT64), .Z(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT34), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT25), .B1(new_n210), .B2(new_n214), .ZN(new_n264));
  AND4_X1   g063(.A1(KEYINPUT25), .A2(new_n216), .A3(new_n217), .A4(new_n214), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n226), .A2(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n235), .A2(new_n238), .ZN(new_n267));
  OAI22_X1  g066(.A1(new_n264), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n255), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n221), .A2(new_n240), .A3(new_n256), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n269), .A2(new_n260), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT34), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  XOR2_X1   g074(.A(G15gat), .B(G43gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT66), .ZN(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n261), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n269), .B2(new_n270), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT32), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n281), .A2(KEYINPUT33), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n261), .B1(new_n257), .B2(new_n258), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT32), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT67), .A4(new_n279), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n279), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(new_n288), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n274), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n273), .B(new_n294), .C1(new_n285), .C2(new_n290), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT68), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT36), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(KEYINPUT68), .B(KEYINPUT36), .C1(new_n296), .C2(new_n297), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g102(.A1(G226gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n268), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT70), .ZN(new_n308));
  AND2_X1   g107(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n310));
  OAI21_X1  g109(.A(G218gat), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G204gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G197gat), .ZN(new_n315));
  INV_X1    g114(.A(G197gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G204gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n308), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G218gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G211gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G218gat), .ZN(new_n325));
  AND4_X1   g124(.A1(new_n315), .A2(new_n317), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT71), .B1(new_n313), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT69), .B(G211gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT22), .B1(new_n328), .B2(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n315), .A2(new_n317), .A3(new_n323), .A4(new_n325), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n321), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT29), .B1(new_n221), .B2(new_n240), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n306), .B(new_n333), .C1(new_n334), .C2(new_n305), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n220), .A2(new_n215), .B1(new_n232), .B2(new_n239), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n304), .B1(new_n337), .B2(KEYINPUT29), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n333), .B1(new_n338), .B2(new_n306), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n303), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT73), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n313), .A2(new_n326), .A3(KEYINPUT71), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n346), .A2(new_n347), .B1(new_n308), .B2(new_n320), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n305), .B1(new_n268), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n304), .B1(new_n221), .B2(new_n240), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(KEYINPUT72), .A3(new_n335), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n340), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n335), .A3(new_n344), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT30), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT30), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n355), .A2(KEYINPUT74), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT74), .B1(new_n355), .B2(new_n358), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n354), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT40), .ZN(new_n362));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT75), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(G155gat), .A3(G162gat), .ZN(new_n366));
  INV_X1    g165(.A(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G162gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(G141gat), .A2(G148gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(KEYINPUT2), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT76), .B1(new_n371), .B2(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(G141gat), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n380));
  NAND2_X1  g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OR3_X1    g181(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n376), .A2(new_n382), .B1(new_n363), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n375), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n363), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT76), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n380), .B1(new_n379), .B2(new_n381), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n364), .A2(new_n366), .A3(new_n369), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n374), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n385), .A2(new_n394), .A3(new_n255), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n389), .A2(new_n392), .A3(new_n251), .A4(new_n254), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n376), .A2(new_n382), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n399), .A2(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n256), .A2(new_n400), .A3(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n255), .B1(new_n375), .B2(new_n384), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n396), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT39), .B1(new_n415), .B2(new_n404), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n402), .B2(new_n404), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n362), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n395), .A2(new_n398), .A3(new_n403), .A4(new_n401), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n415), .B2(new_n404), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n419), .A2(KEYINPUT5), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n411), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n413), .A2(new_n417), .A3(new_n362), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n361), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT85), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT85), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n361), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT37), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n352), .A2(new_n432), .A3(new_n335), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n352), .A2(KEYINPUT86), .A3(new_n335), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n352), .A2(new_n335), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT38), .B1(new_n438), .B2(KEYINPUT37), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n345), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n355), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n344), .B1(new_n435), .B2(new_n436), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n340), .A2(KEYINPUT37), .A3(new_n353), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n398), .A2(new_n401), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n448), .A2(new_n420), .A3(new_n403), .A4(new_n395), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n419), .A2(new_n421), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n412), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n424), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT6), .B(new_n411), .C1(new_n422), .C2(new_n423), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT78), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n412), .B1(new_n449), .B2(new_n450), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(KEYINPUT6), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT87), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n456), .A3(KEYINPUT6), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n453), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n429), .A2(new_n431), .B1(new_n446), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G228gat), .ZN(new_n466));
  INV_X1    g265(.A(G233gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n333), .B1(new_n349), .B2(new_n394), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n333), .A2(KEYINPUT82), .A3(new_n349), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n348), .B2(KEYINPUT29), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n471), .A2(new_n473), .A3(new_n393), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n468), .B(new_n470), .C1(new_n474), .C2(new_n400), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n318), .B1(new_n311), .B2(new_n312), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n307), .ZN(new_n478));
  INV_X1    g277(.A(new_n307), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT80), .B(new_n479), .C1(new_n329), .C2(new_n318), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n478), .B(new_n480), .C1(new_n332), .C2(new_n327), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n349), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT81), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n484), .A3(new_n349), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n393), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n400), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n469), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n475), .B1(new_n488), .B2(new_n468), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT83), .B1(new_n489), .B2(G22gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT31), .B(G50gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G22gat), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n475), .C1(new_n488), .C2(new_n468), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT3), .B1(new_n482), .B2(KEYINPUT81), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n400), .B1(new_n498), .B2(new_n485), .ZN(new_n499));
  OAI22_X1  g298(.A1(new_n499), .A2(new_n469), .B1(new_n466), .B2(new_n467), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n495), .B1(new_n500), .B2(new_n475), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n490), .A2(new_n494), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n489), .A2(G22gat), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(KEYINPUT83), .A3(new_n496), .A4(new_n493), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n302), .B1(new_n465), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n452), .A2(new_n460), .A3(new_n462), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT79), .B1(new_n508), .B2(new_n361), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n354), .A2(new_n357), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n452), .A2(new_n460), .A3(new_n462), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT79), .ZN(new_n512));
  INV_X1    g311(.A(new_n360), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n355), .A2(KEYINPUT74), .A3(new_n358), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n505), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n296), .A2(new_n297), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n504), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT35), .B1(new_n520), .B2(new_n517), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT35), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n510), .A2(new_n522), .A3(new_n515), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n464), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n524), .A2(new_n504), .A3(new_n502), .A4(new_n519), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n507), .A2(new_n518), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G43gat), .B(G50gat), .Z(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT14), .B(G29gat), .Z(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G36gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n528), .A2(new_n529), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n534), .B(new_n537), .C1(new_n530), .C2(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  XNOR2_X1  g345(.A(G99gat), .B(G106gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548));
  INV_X1    g347(.A(G85gat), .ZN(new_n549));
  INV_X1    g348(.A(G92gat), .ZN(new_n550));
  AOI22_X1  g349(.A1(KEYINPUT8), .A2(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n547), .B1(new_n546), .B2(new_n551), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n542), .B(new_n544), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT95), .Z(new_n556));
  INV_X1    g355(.A(KEYINPUT41), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n541), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n552), .A2(new_n553), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n554), .B2(new_n561), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT96), .B1(new_n562), .B2(new_n563), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n556), .A2(new_n557), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G134gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G162gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT97), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n574), .B(new_n571), .C1(new_n566), .C2(KEYINPUT96), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n567), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n567), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G15gat), .B(G22gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT16), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(G1gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(G1gat), .B2(new_n580), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G8gat), .ZN(new_n584));
  XOR2_X1   g383(.A(G57gat), .B(G64gat), .Z(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT92), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n585), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT92), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n593), .A2(new_n585), .A3(KEYINPUT92), .A4(new_n589), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n584), .B1(KEYINPUT21), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n598), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n597), .A2(KEYINPUT93), .A3(KEYINPUT21), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT93), .B1(new_n597), .B2(KEYINPUT21), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n609));
  OR3_X1    g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n609), .B1(new_n607), .B2(new_n608), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n610), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n603), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(new_n602), .A3(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n579), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT98), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n579), .A2(new_n623), .A3(new_n620), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n597), .A2(new_n560), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n595), .B(new_n596), .C1(new_n552), .C2(new_n553), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n597), .A2(new_n560), .A3(KEYINPUT10), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n628), .ZN(new_n634));
  INV_X1    g433(.A(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n633), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n631), .A2(KEYINPUT99), .A3(new_n632), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n636), .ZN(new_n646));
  INV_X1    g445(.A(new_n639), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n641), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n625), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n584), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n542), .A2(new_n650), .A3(new_n544), .ZN(new_n651));
  NAND2_X1  g450(.A1(G229gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n559), .A2(new_n584), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n652), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n541), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n652), .B(KEYINPUT13), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT90), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G113gat), .B(G141gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G169gat), .B(G197gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT89), .B(KEYINPUT12), .Z(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n662), .A2(new_n663), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n527), .A2(new_n649), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n508), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT101), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT100), .B(G1gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n361), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(G8gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT16), .B(G8gat), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(KEYINPUT42), .B2(new_n684), .ZN(G1325gat));
  INV_X1    g485(.A(G15gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n676), .A2(new_n687), .A3(new_n519), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n676), .A2(new_n302), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(G1326gat));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  INV_X1    g490(.A(new_n675), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n526), .A2(new_n506), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n649), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n696), .A3(new_n649), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n691), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n695), .A2(new_n691), .A3(new_n697), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(G1327gat));
  NAND2_X1  g503(.A1(new_n429), .A2(new_n431), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n459), .A2(new_n463), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n443), .A2(new_n444), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT38), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n356), .B1(new_n443), .B2(new_n439), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n706), .A2(new_n708), .A3(new_n452), .A4(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n705), .A2(new_n504), .A3(new_n710), .A4(new_n502), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n300), .A2(new_n301), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n518), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n521), .A2(new_n525), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n579), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n620), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n648), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n692), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n508), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n531), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n723), .B2(new_n722), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n715), .A2(new_n721), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n531), .A3(new_n508), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(G1328gat));
  INV_X1    g528(.A(G36gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n726), .A2(new_n730), .A3(new_n361), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT46), .Z(new_n732));
  AND3_X1   g531(.A1(new_n718), .A2(new_n361), .A3(new_n721), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n730), .B2(new_n733), .ZN(G1329gat));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n302), .A3(new_n721), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n283), .A2(new_n284), .A3(new_n275), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n292), .B1(new_n286), .B2(KEYINPUT32), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT67), .B1(new_n737), .B2(new_n289), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n295), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n273), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n291), .A2(new_n274), .A3(new_n295), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n735), .A2(G43gat), .B1(new_n726), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g544(.A1(new_n716), .A2(new_n505), .A3(new_n721), .A4(new_n717), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n720), .A2(G50gat), .A3(new_n579), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n693), .A2(new_n748), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n747), .A2(new_n749), .B1(KEYINPUT105), .B2(KEYINPUT48), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1331gat));
  INV_X1    g551(.A(new_n648), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n527), .A2(new_n692), .A3(new_n625), .A4(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n508), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  INV_X1    g556(.A(new_n361), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  AOI21_X1  g562(.A(new_n587), .B1(new_n755), .B2(new_n302), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n742), .A2(G71gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n755), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n754), .A2(new_n506), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n588), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n620), .A2(new_n675), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n715), .B2(KEYINPUT107), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n526), .B2(new_n579), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n772), .A2(new_n774), .A3(KEYINPUT51), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT51), .B1(new_n772), .B2(new_n774), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n777), .A2(new_n549), .A3(new_n508), .A4(new_n753), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n771), .A2(new_n648), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n718), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n511), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G85gat), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n781), .A2(new_n779), .A3(new_n511), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n778), .B1(new_n783), .B2(new_n784), .ZN(G1336gat));
  NOR3_X1   g584(.A1(new_n758), .A2(new_n648), .A3(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n716), .A2(new_n361), .A3(new_n717), .A4(new_n780), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G92gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n772), .B2(new_n774), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n786), .B1(new_n775), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n790), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n796), .B2(KEYINPUT52), .ZN(new_n797));
  AOI211_X1 g596(.A(KEYINPUT109), .B(new_n788), .C1(new_n795), .C2(new_n790), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(G1337gat));
  NOR3_X1   g598(.A1(new_n742), .A2(G99gat), .A3(new_n648), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n777), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G99gat), .B1(new_n781), .B2(new_n712), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1338gat));
  INV_X1    g602(.A(G106gat), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n718), .A2(new_n780), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n505), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n775), .A2(new_n794), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n506), .A2(G106gat), .A3(new_n648), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n777), .A2(new_n808), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  OAI21_X1  g612(.A(G106gat), .B1(new_n781), .B2(new_n506), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n629), .A2(new_n635), .A3(new_n630), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT54), .B(new_n633), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n643), .A2(new_n823), .A3(new_n644), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n822), .A2(new_n824), .A3(KEYINPUT55), .A4(new_n647), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n640), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT111), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n828), .A3(new_n640), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n822), .A2(new_n824), .A3(new_n647), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n656), .A2(new_n657), .A3(new_n661), .A4(new_n671), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n659), .A2(new_n660), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n669), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n577), .A2(new_n578), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n817), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n578), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n576), .A3(new_n838), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n826), .A2(KEYINPUT111), .B1(new_n831), .B2(new_n830), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n843), .A2(KEYINPUT112), .A3(new_n829), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n579), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n753), .A2(new_n839), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT113), .B1(new_n648), .B2(new_n838), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n844), .A2(new_n675), .A3(new_n829), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n719), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n622), .A2(new_n692), .A3(new_n624), .A4(new_n648), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n520), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n508), .A3(new_n758), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n692), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n675), .A2(new_n243), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT114), .Z(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n857), .B2(new_n860), .ZN(G1340gat));
  NOR2_X1   g660(.A1(new_n857), .A2(new_n648), .ZN(new_n862));
  XNOR2_X1  g661(.A(KEYINPUT115), .B(G120gat), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n862), .B(new_n863), .ZN(G1341gat));
  NOR2_X1   g663(.A1(new_n857), .A2(new_n719), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(new_n249), .ZN(G1342gat));
  NAND2_X1  g665(.A1(new_n847), .A2(new_n758), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT116), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n856), .A2(new_n247), .A3(new_n508), .A4(new_n869), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT56), .Z(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n857), .B2(new_n579), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1343gat));
  NAND2_X1  g672(.A1(new_n758), .A2(new_n508), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n302), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n506), .B1(new_n854), .B2(new_n855), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n855), .ZN(new_n880));
  INV_X1    g679(.A(new_n826), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  XNOR2_X1  g681(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n830), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n830), .B2(new_n883), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n675), .B(new_n881), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n753), .A2(new_n839), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(KEYINPUT119), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n579), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT119), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n841), .B(new_n845), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n880), .B1(new_n891), .B2(new_n719), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT57), .B1(new_n892), .B2(new_n506), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n879), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G141gat), .B1(new_n894), .B2(new_n692), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n712), .A2(new_n505), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n508), .B1(new_n896), .B2(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(KEYINPUT120), .B2(new_n896), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n854), .A2(new_n855), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(new_n758), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n377), .A3(new_n675), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n895), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1344gat));
  OAI22_X1  g706(.A1(new_n889), .A2(new_n890), .B1(new_n833), .B2(new_n840), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n880), .B1(new_n908), .B2(new_n719), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n505), .A2(new_n878), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n877), .A2(new_n878), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n875), .A2(new_n753), .ZN(new_n912));
  OAI21_X1  g711(.A(G148gat), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT59), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n879), .A2(new_n893), .A3(new_n753), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n378), .A2(KEYINPUT59), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n915), .A2(KEYINPUT121), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT121), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n378), .A3(new_n753), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1345gat));
  OAI21_X1  g720(.A(G155gat), .B1(new_n894), .B2(new_n719), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n367), .A3(new_n620), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n894), .B2(new_n579), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n900), .A2(new_n368), .A3(new_n869), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  INV_X1    g726(.A(new_n520), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n758), .A2(new_n508), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n899), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n675), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n856), .A2(KEYINPUT122), .A3(new_n929), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT122), .B1(new_n856), .B2(new_n929), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n692), .A2(new_n207), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n931), .A2(new_n208), .A3(new_n753), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n934), .A2(new_n648), .A3(new_n935), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n208), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(KEYINPUT123), .B(new_n939), .C1(new_n940), .C2(new_n208), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1349gat));
  AND2_X1   g744(.A1(new_n620), .A2(new_n229), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT124), .B1(new_n931), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n934), .A2(new_n719), .A3(new_n935), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n211), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n951), .B(new_n947), .C1(new_n948), .C2(new_n211), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n931), .A2(new_n212), .A3(new_n847), .ZN(new_n954));
  INV_X1    g753(.A(new_n935), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(new_n847), .A3(new_n933), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  XOR2_X1   g759(.A(KEYINPUT126), .B(G197gat), .Z(new_n961));
  OR2_X1    g760(.A1(new_n877), .A2(new_n878), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n909), .A2(new_n910), .ZN(new_n963));
  INV_X1    g762(.A(new_n929), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n302), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n961), .B1(new_n966), .B2(new_n692), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n896), .B(new_n964), .C1(new_n854), .C2(new_n855), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT125), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n692), .A2(new_n961), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n314), .A3(new_n753), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n976), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(KEYINPUT62), .A3(new_n974), .ZN(new_n979));
  OAI21_X1  g778(.A(G204gat), .B1(new_n966), .B2(new_n648), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(G1353gat));
  NAND4_X1  g780(.A1(new_n962), .A2(new_n963), .A3(new_n620), .A4(new_n965), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n719), .A2(new_n328), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n983), .A2(new_n984), .B1(new_n969), .B2(new_n985), .ZN(G1354gat));
  OAI21_X1  g785(.A(G218gat), .B1(new_n966), .B2(new_n579), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n847), .A2(new_n322), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n969), .B2(new_n988), .ZN(G1355gat));
endmodule


