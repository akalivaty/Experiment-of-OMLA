//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  NOR2_X1   g000(.A1(KEYINPUT75), .A2(G125), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT75), .A2(G125), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G140), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(KEYINPUT16), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(new_n189), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT16), .A2(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(G146), .A3(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT74), .B1(new_n204), .B2(G128), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n206), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G110), .ZN(new_n210));
  XOR2_X1   g024(.A(G119), .B(G128), .Z(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT24), .B(G110), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n202), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G110), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n191), .A2(G140), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n193), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n215), .A2(new_n216), .B1(new_n199), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT76), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n219), .A2(new_n220), .A3(new_n201), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n219), .B2(new_n201), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n213), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n224), .B(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G902), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n213), .B(new_n227), .C1(new_n221), .C2(new_n222), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n230), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G217), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(G234), .B2(new_n230), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n229), .A2(new_n231), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n240), .A2(G902), .A3(new_n238), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n199), .A2(G143), .ZN(new_n248));
  OAI22_X1  g062(.A1(new_n245), .A2(new_n247), .B1(new_n248), .B2(G128), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT69), .B1(new_n251), .B2(new_n245), .ZN(new_n252));
  AND4_X1   g066(.A1(KEYINPUT69), .A2(new_n245), .A3(new_n247), .A4(new_n248), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G134), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n255), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n259), .B2(G134), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n256), .A2(KEYINPUT67), .A3(G137), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n256), .A2(G137), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(KEYINPUT11), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n263), .A2(new_n264), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(KEYINPUT68), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n271), .B(new_n273), .C1(G134), .C2(new_n259), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n254), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n247), .A2(new_n248), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  OR2_X1    g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n280), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n251), .B2(KEYINPUT65), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n263), .A2(new_n264), .A3(new_n269), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n264), .B1(new_n263), .B2(new_n269), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n254), .A2(new_n289), .A3(new_n275), .A4(new_n270), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n277), .A2(KEYINPUT30), .A3(new_n288), .A4(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G116), .B(G119), .ZN(new_n292));
  NAND2_X1  g106(.A1(KEYINPUT2), .A2(G113), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT2), .A2(G113), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(KEYINPUT70), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(KEYINPUT70), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n292), .B(new_n293), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n294), .B(KEYINPUT70), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n292), .B1(new_n299), .B2(new_n293), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n303));
  INV_X1    g117(.A(new_n276), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n282), .A2(new_n284), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n263), .A2(new_n269), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G131), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n307), .B2(new_n270), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n303), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n291), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n277), .A2(new_n301), .A3(new_n288), .A4(new_n290), .ZN(new_n311));
  INV_X1    g125(.A(G237), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT72), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G237), .ZN(new_n315));
  AOI21_X1  g129(.A(G953), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G210), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT26), .B(G101), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT31), .B1(new_n310), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n288), .A2(new_n301), .A3(new_n276), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n301), .B1(new_n288), .B2(new_n276), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n326), .B(new_n328), .C1(new_n311), .C2(new_n325), .ZN(new_n329));
  INV_X1    g143(.A(new_n321), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n291), .A2(new_n309), .A3(new_n302), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT31), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n311), .A4(new_n321), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G472), .A2(G902), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT32), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT32), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n339), .A3(new_n336), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n326), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n277), .A2(new_n288), .A3(new_n290), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n302), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n311), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n345), .B2(KEYINPUT28), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n330), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n332), .A2(new_n311), .A3(new_n330), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n251), .A2(KEYINPUT69), .A3(new_n245), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n355), .A2(new_n250), .B1(G131), .B2(new_n274), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n289), .B1(new_n356), .B2(new_n270), .ZN(new_n357));
  INV_X1    g171(.A(new_n290), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(KEYINPUT28), .A3(new_n301), .A4(new_n288), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n327), .B1(new_n325), .B2(new_n324), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n330), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n347), .B1(new_n350), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G472), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n243), .B1(new_n341), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n367));
  OR2_X1    g181(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n368));
  INV_X1    g182(.A(G107), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G104), .ZN(new_n370));
  AND2_X1   g184(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n369), .A2(G104), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G107), .ZN(new_n377));
  NOR2_X1   g191(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n372), .A2(new_n373), .A3(new_n375), .A4(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G101), .B1(new_n377), .B2(new_n374), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n254), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n381), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n249), .B1(new_n353), .B2(new_n354), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n307), .A2(new_n270), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(KEYINPUT12), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT12), .B1(new_n386), .B2(new_n387), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT81), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n374), .B1(new_n378), .B2(new_n377), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n372), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n373), .B1(new_n391), .B2(new_n372), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n394), .B(new_n285), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n383), .B2(new_n384), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n387), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n382), .B2(new_n398), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n380), .A2(new_n381), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(KEYINPUT79), .A3(KEYINPUT10), .A4(new_n254), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n400), .A2(new_n401), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n383), .A2(new_n384), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n383), .A2(new_n384), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n387), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n386), .A2(KEYINPUT12), .A3(new_n387), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G140), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n225), .A2(G227), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n390), .A2(new_n406), .A3(new_n414), .A4(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n405), .A2(new_n399), .A3(new_n397), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT79), .B1(new_n408), .B2(KEYINPUT10), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n387), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n406), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n417), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT80), .B(G469), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n406), .A2(new_n422), .A3(new_n418), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n411), .A2(new_n413), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n418), .B1(new_n428), .B2(new_n406), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n230), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n425), .A2(new_n426), .B1(new_n430), .B2(G469), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT9), .B(G234), .ZN(new_n432));
  OAI21_X1  g246(.A(G221), .B1(new_n432), .B2(G902), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT77), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n367), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n419), .A2(new_n424), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n437), .A2(new_n230), .A3(new_n426), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n388), .A2(new_n389), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n420), .A2(new_n387), .A3(new_n421), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n417), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n406), .A2(new_n422), .A3(new_n418), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n444), .B2(new_n230), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT82), .B(new_n436), .C1(new_n438), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n435), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT18), .A2(G131), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n316), .A2(G143), .A3(G214), .ZN(new_n450));
  AOI21_X1  g264(.A(G143), .B1(new_n316), .B2(G214), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n316), .A2(G214), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n246), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n316), .A2(G143), .A3(G214), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n448), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n218), .A2(new_n199), .ZN(new_n457));
  AND2_X1   g271(.A1(KEYINPUT75), .A2(G125), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n187), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n192), .B1(new_n459), .B2(G140), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(new_n199), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n452), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT93), .B(G104), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n465), .B(KEYINPUT95), .Z(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n450), .B2(new_n451), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n454), .A2(new_n264), .A3(new_n455), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(KEYINPUT17), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n200), .B(new_n201), .C1(new_n467), .C2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n462), .B(new_n466), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n452), .A2(new_n456), .A3(new_n461), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT19), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n193), .A2(new_n217), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n199), .B(new_n478), .C1(new_n460), .C2(new_n477), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n201), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n480), .A2(KEYINPUT92), .B1(new_n467), .B2(new_n468), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n201), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n476), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n475), .B1(new_n484), .B2(new_n465), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(KEYINPUT92), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n469), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n462), .ZN(new_n488));
  INV_X1    g302(.A(new_n465), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(KEYINPUT94), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n474), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(G475), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT94), .B1(new_n488), .B2(new_n489), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n475), .B(new_n465), .C1(new_n487), .C2(new_n462), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n473), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n492), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT96), .B(G475), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n470), .A2(new_n472), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n489), .B1(new_n503), .B2(new_n476), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n473), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n505), .B2(new_n230), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(G234), .A2(G237), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(G952), .A3(new_n225), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT21), .B(G898), .Z(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(G902), .A3(G953), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT101), .Z(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT98), .B1(new_n244), .B2(G143), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT98), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n246), .A3(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT13), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n519), .A2(new_n520), .B1(new_n244), .B2(G143), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n520), .B2(new_n519), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G134), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n244), .A2(G143), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n256), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G116), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G122), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n526), .A2(G122), .ZN(new_n529));
  OAI21_X1  g343(.A(G107), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n369), .A3(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n533), .A2(KEYINPUT97), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(KEYINPUT97), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n523), .A2(new_n525), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n532), .ZN(new_n537));
  OR3_X1    g351(.A1(new_n527), .A2(KEYINPUT99), .A3(KEYINPUT14), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n529), .B1(KEYINPUT14), .B2(new_n527), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT99), .B1(new_n527), .B2(KEYINPUT14), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n541), .B2(G107), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT100), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n519), .A2(new_n524), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G134), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n525), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n542), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n536), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n432), .A2(new_n237), .A3(G953), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n536), .B(new_n550), .C1(new_n547), .C2(new_n548), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n554), .B(new_n556), .Z(new_n557));
  NOR3_X1   g371(.A1(new_n508), .A2(new_n515), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G214), .B1(G237), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G210), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n204), .A2(G116), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n526), .A2(G119), .ZN(new_n564));
  AND2_X1   g378(.A1(KEYINPUT83), .A2(KEYINPUT5), .ZN(new_n565));
  NOR2_X1   g379(.A1(KEYINPUT83), .A2(KEYINPUT5), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n526), .A2(G119), .ZN(new_n568));
  OR2_X1    g382(.A1(KEYINPUT83), .A2(KEYINPUT5), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT83), .A2(KEYINPUT5), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n571), .A3(G113), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT84), .ZN(new_n573));
  INV_X1    g387(.A(G113), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n565), .A2(new_n566), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n568), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT84), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n567), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n578), .A3(new_n297), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n383), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n563), .A2(new_n564), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT5), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT87), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT87), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n292), .A2(new_n584), .A3(KEYINPUT5), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n576), .A3(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n404), .A2(KEYINPUT88), .A3(new_n297), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT88), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n583), .A2(new_n576), .A3(new_n585), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n380), .A2(new_n297), .A3(new_n381), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n580), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G122), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT8), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n254), .A2(new_n459), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n282), .A2(new_n284), .A3(new_n195), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT85), .B(G224), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n225), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n600), .A2(KEYINPUT89), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(KEYINPUT7), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n603), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n596), .A2(new_n597), .A3(new_n601), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT90), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n595), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n302), .B(new_n394), .C1(new_n396), .C2(new_n395), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n404), .A2(new_n297), .A3(new_n578), .A4(new_n573), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n593), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n608), .B1(new_n595), .B2(new_n607), .ZN(new_n614));
  OAI211_X1 g428(.A(KEYINPUT91), .B(new_n230), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n611), .ZN(new_n616));
  INV_X1    g430(.A(new_n593), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(KEYINPUT6), .A3(new_n612), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n596), .A2(new_n597), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n599), .B(KEYINPUT86), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT6), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n616), .A2(new_n623), .A3(new_n617), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n595), .A2(new_n607), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT90), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n612), .A3(new_n609), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT91), .B1(new_n629), .B2(new_n230), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n562), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n230), .B1(new_n613), .B2(new_n614), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT91), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n634), .A2(new_n561), .A3(new_n625), .A4(new_n615), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n560), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n366), .A2(new_n447), .A3(new_n558), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  NAND2_X1  g452(.A1(new_n335), .A2(new_n230), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n337), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n243), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n506), .B1(new_n494), .B2(new_n499), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n551), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n552), .A2(new_n553), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n552), .B2(new_n553), .ZN(new_n648));
  OAI21_X1  g462(.A(G478), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n555), .A2(new_n230), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n554), .B2(new_n555), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n643), .A2(new_n515), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n447), .A2(new_n642), .A3(new_n636), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NAND2_X1  g470(.A1(new_n643), .A2(new_n557), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n515), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n636), .A2(new_n447), .A3(new_n658), .A4(new_n642), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT35), .B(G107), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n238), .A2(G902), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n228), .A2(KEYINPUT36), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n223), .B(new_n663), .Z(new_n664));
  AOI22_X1  g478(.A1(new_n236), .A2(new_n238), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n641), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n447), .A2(new_n558), .A3(new_n666), .A4(new_n636), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  AOI21_X1  g483(.A(new_n665), .B1(new_n341), .B2(new_n365), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n512), .A2(G900), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n510), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n657), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n670), .A2(new_n447), .A3(new_n674), .A4(new_n636), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT103), .B(G128), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G30));
  XNOR2_X1  g491(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n672), .B(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n447), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n631), .A2(new_n635), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT38), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n508), .A2(new_n557), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n310), .A2(new_n322), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n321), .B1(new_n344), .B2(new_n311), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT104), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n230), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n687), .A2(KEYINPUT104), .A3(new_n688), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n341), .A2(new_n692), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n559), .A2(new_n686), .A3(new_n665), .A4(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n682), .A2(new_n684), .A3(new_n685), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NOR3_X1   g510(.A1(new_n643), .A2(new_n652), .A3(new_n673), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n670), .A2(new_n447), .A3(new_n636), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR2_X1   g513(.A1(new_n425), .A2(new_n439), .ZN(new_n700));
  INV_X1    g514(.A(new_n433), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n438), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n366), .A2(new_n653), .A3(new_n636), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND4_X1  g519(.A1(new_n366), .A2(new_n658), .A3(new_n636), .A4(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND4_X1  g521(.A1(new_n670), .A2(new_n558), .A3(new_n636), .A4(new_n702), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT106), .B(G119), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G21));
  NOR4_X1   g524(.A1(new_n438), .A2(new_n700), .A3(new_n515), .A4(new_n701), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n323), .B(new_n334), .C1(new_n346), .C2(new_n321), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n639), .A2(G472), .B1(new_n712), .B2(new_n336), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n241), .B1(new_n236), .B2(new_n238), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT107), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n686), .A2(new_n636), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(G122), .Z(G24));
  NAND2_X1  g534(.A1(new_n712), .A2(new_n336), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n640), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n665), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n636), .A3(new_n697), .A4(new_n702), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  INV_X1    g541(.A(G472), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n349), .B2(new_n363), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n338), .B2(new_n340), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n727), .B1(new_n730), .B2(new_n243), .ZN(new_n731));
  INV_X1    g545(.A(new_n340), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n339), .B1(new_n335), .B2(new_n336), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n365), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n714), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n631), .A2(new_n559), .A3(new_n635), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n643), .A2(new_n738), .A3(new_n652), .A4(new_n673), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n425), .A2(new_n426), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n430), .A2(G469), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n701), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n737), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n726), .B1(new_n736), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(new_n631), .A3(new_n559), .A4(new_n635), .ZN(new_n745));
  INV_X1    g559(.A(new_n652), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n508), .A2(new_n746), .A3(KEYINPUT42), .A4(new_n672), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(KEYINPUT109), .A3(new_n731), .A4(new_n735), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n366), .A2(new_n737), .A3(new_n697), .A4(new_n742), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n738), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n744), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NAND4_X1  g567(.A1(new_n366), .A2(new_n737), .A3(new_n674), .A4(new_n742), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n439), .B1(new_n444), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n442), .A2(KEYINPUT45), .A3(new_n443), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n439), .B2(new_n230), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n438), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n433), .A3(new_n680), .ZN(new_n764));
  INV_X1    g578(.A(new_n737), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n643), .B(KEYINPUT110), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT43), .A3(new_n746), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n508), .A2(new_n652), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(KEYINPUT43), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n665), .B1(new_n337), .B2(new_n640), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT44), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n766), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n259), .ZN(G39));
  NAND2_X1  g589(.A1(new_n763), .A2(new_n433), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n697), .A2(new_n730), .A3(new_n243), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n737), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  INV_X1    g595(.A(new_n510), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n770), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n715), .A2(new_n716), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n737), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n438), .A2(new_n700), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n778), .B1(new_n434), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT50), .ZN(new_n792));
  INV_X1    g606(.A(new_n702), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n684), .A2(new_n559), .A3(new_n793), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n785), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n792), .B1(new_n785), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n765), .A2(new_n793), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n783), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n723), .ZN(new_n800));
  INV_X1    g614(.A(new_n693), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n782), .A2(new_n798), .A3(new_n714), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n643), .A3(new_n652), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n790), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n790), .A2(KEYINPUT51), .A3(new_n797), .A4(new_n804), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n799), .A2(new_n731), .A3(new_n735), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT48), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n786), .A2(new_n636), .A3(new_n702), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n643), .A2(new_n652), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  AND4_X1   g627(.A1(G952), .A2(new_n811), .A3(new_n225), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n637), .A2(new_n667), .A3(new_n703), .A4(new_n654), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n706), .B(new_n708), .C1(new_n717), .C2(new_n718), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n737), .A2(new_n723), .A3(new_n697), .A4(new_n742), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n754), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n670), .A2(new_n447), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n508), .A2(new_n557), .A3(new_n673), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(KEYINPUT113), .A3(new_n737), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n670), .A2(new_n737), .A3(new_n447), .A4(new_n823), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n821), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n658), .A2(KEYINPUT112), .A3(new_n636), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT112), .B1(new_n658), .B2(new_n636), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n447), .A2(new_n642), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n819), .A2(new_n828), .A3(new_n752), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n742), .A2(new_n665), .A3(new_n672), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n636), .A3(new_n686), .A4(new_n693), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n675), .A2(new_n698), .A3(new_n836), .A4(new_n724), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT52), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n816), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n824), .A2(new_n827), .ZN(new_n842));
  INV_X1    g656(.A(new_n821), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n752), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n675), .A2(new_n698), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .A3(new_n724), .A4(new_n836), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n837), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n832), .A2(new_n817), .A3(new_n818), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n844), .A2(KEYINPUT53), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n840), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n841), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n839), .A2(new_n851), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(KEYINPUT54), .B2(new_n854), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n815), .A2(new_n855), .B1(G952), .B2(G953), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n714), .A2(new_n559), .A3(new_n436), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT111), .Z(new_n858));
  XOR2_X1   g672(.A(new_n788), .B(KEYINPUT49), .Z(new_n859));
  NOR3_X1   g673(.A1(new_n858), .A2(new_n859), .A3(new_n652), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n801), .A3(new_n767), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n856), .B1(new_n684), .B2(new_n861), .ZN(G75));
  AOI21_X1  g676(.A(new_n230), .B1(new_n839), .B2(new_n851), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(KEYINPUT116), .A3(G210), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n619), .A2(new_n624), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n622), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT55), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT116), .B1(new_n863), .B2(G210), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n225), .A2(G952), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT56), .B1(new_n863), .B2(G210), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n868), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n871), .A2(new_n875), .ZN(G51));
  XNOR2_X1  g690(.A(new_n854), .B(KEYINPUT54), .ZN(new_n877));
  XNOR2_X1  g691(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n439), .A2(new_n230), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n877), .A2(new_n880), .B1(new_n424), .B2(new_n419), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n759), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n881), .A2(new_n882), .B1(new_n884), .B2(new_n863), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n872), .B1(new_n883), .B2(new_n885), .ZN(G54));
  AND2_X1   g700(.A1(KEYINPUT58), .A2(G475), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n863), .A2(new_n497), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n497), .B1(new_n863), .B2(new_n887), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n872), .ZN(G60));
  OR2_X1    g704(.A1(new_n647), .A2(new_n648), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n650), .B(KEYINPUT59), .Z(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n855), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n877), .A2(new_n892), .A3(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n872), .A3(new_n895), .ZN(G63));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  XNOR2_X1  g711(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n237), .A2(new_n230), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n897), .B1(new_n854), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n900), .ZN(new_n902));
  AOI211_X1 g716(.A(KEYINPUT121), .B(new_n902), .C1(new_n839), .C2(new_n851), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n240), .B(KEYINPUT123), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n906), .B2(new_n872), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n854), .A2(new_n900), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n854), .A2(new_n897), .A3(new_n900), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n908), .B(new_n873), .C1(new_n912), .C2(new_n905), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n664), .B(KEYINPUT122), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n907), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g730(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n906), .A2(new_n872), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(KEYINPUT61), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(G66));
  AOI21_X1  g735(.A(new_n225), .B1(new_n511), .B2(new_n598), .ZN(new_n922));
  INV_X1    g736(.A(new_n850), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n225), .ZN(new_n924));
  INV_X1    g738(.A(G898), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n866), .B1(new_n925), .B2(G953), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n924), .B(new_n926), .ZN(G69));
  NAND2_X1  g741(.A1(new_n291), .A2(new_n309), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n478), .B1(new_n460), .B2(new_n477), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(G900), .A2(G953), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n764), .A2(new_n718), .A3(new_n736), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n780), .A2(new_n754), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n774), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n845), .A2(new_n724), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n933), .A2(new_n752), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n930), .B(new_n931), .C1(new_n936), .C2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n657), .B1(new_n643), .B2(new_n652), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT126), .Z(new_n939));
  NOR3_X1   g753(.A1(new_n681), .A2(new_n730), .A3(new_n243), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n737), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n780), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n935), .A2(new_n695), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n942), .A2(new_n934), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  AOI21_X1  g763(.A(G953), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n930), .B(KEYINPUT125), .Z(new_n951));
  OAI21_X1  g765(.A(new_n937), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n225), .B1(G227), .B2(G900), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G72));
  AOI21_X1  g768(.A(new_n330), .B1(new_n332), .B2(new_n311), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n948), .A2(new_n850), .A3(new_n949), .ZN(new_n956));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n350), .A2(new_n955), .A3(new_n959), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n841), .B2(new_n852), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n958), .B1(new_n936), .B2(new_n923), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n872), .B1(new_n963), .B2(new_n350), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(G57));
endmodule


