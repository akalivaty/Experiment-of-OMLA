//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT11), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(G169gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT92), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT92), .B1(new_n214), .B2(new_n208), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n213), .A2(new_n215), .B1(new_n209), .B2(new_n210), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  OR2_X1    g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT93), .B(G50gat), .Z(new_n222));
  OAI211_X1 g021(.A(new_n217), .B(new_n219), .C1(new_n222), .C2(G43gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n220), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n211), .A2(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT94), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT94), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n221), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n232), .B1(new_n235), .B2(KEYINPUT96), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(G1gat), .B2(new_n233), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT97), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT97), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n231), .A2(new_n243), .A3(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT95), .B(KEYINPUT17), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n240), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n226), .A3(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n245), .A2(KEYINPUT18), .A3(new_n246), .A4(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n231), .A2(new_n243), .A3(new_n240), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n243), .B1(new_n231), .B2(new_n240), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n253), .A2(new_n254), .B1(new_n240), .B2(new_n231), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n246), .B(KEYINPUT13), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n251), .B(new_n246), .C1(new_n254), .C2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n206), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT99), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT98), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(KEYINPUT98), .A3(new_n261), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n206), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n264), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n269), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n258), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT98), .B1(new_n260), .B2(new_n261), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n274), .A3(KEYINPUT99), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n263), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT102), .B(G85gat), .ZN(new_n277));
  INV_X1    g076(.A(G92gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G99gat), .A2(G106gat), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n277), .A2(new_n278), .B1(KEYINPUT8), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G85gat), .A2(G92gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT7), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G99gat), .B(G106gat), .Z(new_n284));
  OR2_X1    g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT103), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n284), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT100), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G57gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(G64gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G71gat), .B(G78gat), .ZN(new_n292));
  AND2_X1   g091(.A1(G71gat), .A2(G78gat), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n291), .B(new_n292), .C1(KEYINPUT9), .C2(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(G57gat), .A2(G64gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G57gat), .A2(G64gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n295), .A2(KEYINPUT9), .A3(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(new_n292), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n288), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n284), .B2(new_n283), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n285), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n286), .A2(KEYINPUT10), .A3(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G230gat), .A2(G233gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n303), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G120gat), .B(G148gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT106), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G204gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n318), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n308), .A2(new_n311), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n276), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT77), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G141gat), .ZN(new_n329));
  INV_X1    g128(.A(G141gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G148gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n334), .B(KEYINPUT2), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n327), .A2(new_n332), .A3(new_n333), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339));
  NOR2_X1   g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G141gat), .B(G148gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(KEYINPUT2), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n338), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT78), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n338), .A2(new_n346), .A3(new_n343), .A4(new_n339), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n338), .A2(new_n343), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n350));
  INV_X1    g149(.A(G113gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(G120gat), .ZN(new_n352));
  INV_X1    g151(.A(G120gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n352), .B(new_n354), .C1(G113gat), .C2(new_n353), .ZN(new_n355));
  XOR2_X1   g154(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n356));
  NOR2_X1   g155(.A1(G127gat), .A2(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G127gat), .A2(G134gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n355), .B(new_n356), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n357), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(KEYINPUT71), .A3(new_n358), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n359), .B2(new_n357), .ZN(new_n364));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n362), .B(new_n364), .C1(KEYINPUT1), .C2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(KEYINPUT3), .A2(new_n349), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT79), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n348), .A2(new_n370), .A3(new_n367), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n360), .A2(new_n366), .ZN(new_n375));
  OR3_X1    g174(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n349), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT4), .B1(new_n375), .B2(new_n349), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(KEYINPUT82), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n377), .A2(KEYINPUT82), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n374), .A2(KEYINPUT5), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  NAND2_X1  g186(.A1(new_n376), .A2(new_n377), .ZN(new_n388));
  INV_X1    g187(.A(new_n371), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n370), .B1(new_n348), .B2(new_n367), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n373), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n372), .A2(KEYINPUT80), .A3(new_n373), .A4(new_n388), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n375), .B(new_n349), .ZN(new_n396));
  INV_X1    g195(.A(new_n373), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT5), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n382), .B(new_n387), .C1(new_n395), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  INV_X1    g200(.A(new_n387), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n393), .B2(new_n394), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(new_n381), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT6), .B(new_n402), .C1(new_n403), .C2(new_n381), .ZN(new_n406));
  XNOR2_X1  g205(.A(G197gat), .B(G204gat), .ZN(new_n407));
  INV_X1    g206(.A(G211gat), .ZN(new_n408));
  INV_X1    g207(.A(G218gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(KEYINPUT22), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G211gat), .B(G218gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(G183gat), .ZN(new_n417));
  INV_X1    g216(.A(G183gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(KEYINPUT27), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT67), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G190gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT66), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT66), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G190gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(KEYINPUT27), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT67), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT28), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430));
  NOR2_X1   g229(.A1(G169gat), .A2(G176gat), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT26), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT69), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n422), .A2(new_n424), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT68), .B1(new_n417), .B2(new_n419), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n416), .A2(G183gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT68), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n429), .B(new_n437), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT25), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT24), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n425), .A2(new_n418), .B1(new_n450), .B2(new_n446), .ZN(new_n451));
  NAND3_X1  g250(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT65), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n449), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n431), .A2(KEYINPUT23), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT23), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(G169gat), .B2(G176gat), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n455), .A2(new_n434), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n447), .A2(KEYINPUT24), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n452), .B1(G183gat), .B2(G190gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n454), .A2(new_n458), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n415), .B1(new_n448), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n465), .B(KEYINPUT76), .Z(new_n466));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n445), .B2(new_n447), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n429), .A2(new_n437), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n442), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n441), .B1(new_n426), .B2(new_n440), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n425), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT28), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n470), .A2(KEYINPUT70), .A3(new_n474), .A4(new_n446), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n464), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT75), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n464), .B1(new_n468), .B2(new_n475), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT75), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT29), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n413), .B(new_n466), .C1(new_n483), .C2(new_n415), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n415), .A3(new_n482), .ZN(new_n485));
  INV_X1    g284(.A(new_n413), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n415), .A2(KEYINPUT29), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n448), .B2(new_n464), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G8gat), .B(G36gat), .Z(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(G64gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(new_n278), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n405), .A2(new_n406), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n493), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT37), .B1(new_n484), .B2(new_n489), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n466), .B1(new_n483), .B2(new_n415), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n502), .B2(new_n486), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n413), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n494), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n500), .A2(new_n497), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT88), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT88), .B1(new_n506), .B2(new_n507), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n496), .B(new_n501), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n484), .A2(new_n489), .A3(new_n493), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n511), .A3(KEYINPUT30), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n513), .A3(new_n494), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n380), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n373), .B1(new_n516), .B2(new_n372), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT39), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n402), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR3_X1    g318(.A1(new_n396), .A2(KEYINPUT84), .A3(new_n397), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT84), .B1(new_n396), .B2(new_n397), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT39), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT85), .Z(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n523), .B2(new_n517), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT86), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT40), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n515), .A2(new_n527), .A3(new_n404), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G50gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n339), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n349), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT29), .B1(new_n345), .B2(new_n347), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(new_n486), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G22gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(G22gat), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n531), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT83), .B1(new_n534), .B2(new_n486), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(G228gat), .A3(G233gat), .ZN(new_n543));
  XOR2_X1   g342(.A(G78gat), .B(G106gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT31), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n543), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n538), .A2(new_n531), .A3(new_n539), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n546), .B1(new_n550), .B2(new_n540), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n510), .A2(new_n530), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n405), .A2(new_n406), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n559));
  XNOR2_X1  g358(.A(G15gat), .B(G43gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G71gat), .ZN(new_n561));
  INV_X1    g360(.A(G99gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n375), .B1(new_n476), .B2(new_n477), .ZN(new_n564));
  INV_X1    g363(.A(new_n375), .ZN(new_n565));
  AOI211_X1 g364(.A(new_n565), .B(new_n464), .C1(new_n468), .C2(new_n475), .ZN(new_n566));
  INV_X1    g365(.A(G227gat), .ZN(new_n567));
  INV_X1    g366(.A(G233gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n564), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n563), .B1(new_n571), .B2(KEYINPUT33), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT32), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT34), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n478), .A2(new_n565), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n481), .A2(new_n375), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT34), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n569), .B1(new_n575), .B2(new_n576), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n574), .B2(new_n579), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n572), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT34), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n578), .B1(new_n577), .B2(KEYINPUT32), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n572), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n559), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(KEYINPUT36), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n584), .A2(KEYINPUT74), .A3(new_n558), .A4(new_n590), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n553), .A2(new_n557), .A3(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT89), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT89), .B1(new_n584), .B2(new_n590), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI221_X4 g401(.A(KEYINPUT35), .B1(new_n405), .B2(new_n406), .C1(new_n512), .C2(new_n514), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n552), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n584), .A2(new_n590), .A3(new_n552), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT91), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n512), .A2(new_n514), .B1(new_n406), .B2(new_n405), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT91), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n584), .A2(new_n552), .A3(new_n609), .A4(new_n590), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT35), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n599), .B1(new_n597), .B2(new_n598), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n584), .A2(KEYINPUT89), .A3(new_n590), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n552), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n512), .A2(new_n514), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n555), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT90), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n605), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n324), .B1(new_n596), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n299), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(KEYINPUT21), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G127gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n240), .B1(KEYINPUT21), .B2(new_n622), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT101), .B(G155gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n630), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n288), .A2(new_n250), .A3(new_n248), .ZN(new_n635));
  NAND3_X1  g434(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n286), .A2(new_n287), .A3(new_n231), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT104), .B(G134gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G162gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n641), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n642), .B2(new_n645), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT105), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n621), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT107), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n621), .A2(new_n654), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n556), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g457(.A(new_n616), .B1(new_n653), .B2(new_n655), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n234), .B2(new_n232), .ZN(new_n660));
  NOR2_X1   g459(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n232), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT42), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(KEYINPUT42), .B2(new_n662), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n656), .A2(new_n666), .A3(new_n602), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n595), .B1(new_n653), .B2(new_n655), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT108), .ZN(G1326gat));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n656), .B2(new_n554), .ZN(new_n672));
  AOI211_X1 g471(.A(KEYINPUT109), .B(new_n552), .C1(new_n653), .C2(new_n655), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n655), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n654), .B1(new_n621), .B2(new_n651), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n554), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT109), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n656), .A2(new_n671), .A3(new_n554), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n674), .A2(new_n681), .A3(G22gat), .ZN(new_n682));
  AOI21_X1  g481(.A(G22gat), .B1(new_n674), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n553), .A2(new_n557), .A3(new_n595), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT113), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n620), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n605), .A2(new_n612), .A3(new_n619), .A4(KEYINPUT113), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n685), .B1(new_n690), .B2(new_n649), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n596), .A2(new_n620), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n648), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n634), .B(KEYINPUT111), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n323), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT112), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n555), .ZN(new_n699));
  INV_X1    g498(.A(new_n634), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n621), .A2(new_n700), .A3(new_n648), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n209), .A3(new_n556), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n704), .ZN(G1328gat));
  OAI21_X1  g504(.A(G36gat), .B1(new_n698), .B2(new_n616), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n210), .A3(new_n515), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT46), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(new_n602), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(G43gat), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n701), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n595), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n694), .A2(new_n713), .A3(new_n697), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(G43gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n716), .ZN(new_n718));
  AOI211_X1 g517(.A(new_n718), .B(new_n712), .C1(new_n714), .C2(G43gat), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n719), .ZN(G1330gat));
  NAND4_X1  g519(.A1(new_n691), .A2(new_n554), .A3(new_n693), .A4(new_n697), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT115), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  INV_X1    g523(.A(new_n222), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n701), .A2(new_n725), .A3(new_n554), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT48), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n721), .A2(new_n222), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(new_n727), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n726), .A2(new_n728), .B1(KEYINPUT48), .B2(new_n730), .ZN(G1331gat));
  INV_X1    g530(.A(new_n651), .ZN(new_n732));
  INV_X1    g531(.A(new_n276), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n690), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n322), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n556), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g537(.A1(new_n735), .A2(new_n616), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n735), .B2(new_n595), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n710), .A2(G71gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n735), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n736), .A2(new_n554), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n634), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n694), .A2(new_n322), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n555), .A3(new_n277), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n688), .A2(new_n689), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n596), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n648), .A3(new_n751), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n755), .A2(new_n758), .A3(new_n648), .A4(new_n751), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n556), .A3(new_n322), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n753), .B1(new_n761), .B2(new_n277), .ZN(G1336gat));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n757), .A2(new_n515), .A3(new_n322), .A4(new_n759), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(new_n278), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n515), .A2(G92gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n752), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n763), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n278), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n769), .B(KEYINPUT52), .C1(new_n752), .C2(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1337gat));
  NOR3_X1   g570(.A1(new_n752), .A2(new_n562), .A3(new_n595), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n760), .A2(new_n602), .A3(new_n322), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n562), .ZN(G1338gat));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n554), .A3(new_n322), .A4(new_n759), .ZN(new_n775));
  INV_X1    g574(.A(G106gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(KEYINPUT53), .ZN(new_n779));
  AND4_X1   g578(.A1(new_n322), .A2(new_n691), .A3(new_n693), .A4(new_n751), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n552), .A2(new_n776), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(KEYINPUT53), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n777), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n777), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n515), .A2(new_n555), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n246), .B1(new_n245), .B2(new_n251), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT117), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n255), .A2(new_n257), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(KEYINPUT117), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n205), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT99), .B1(new_n271), .B2(new_n274), .ZN(new_n795));
  NOR4_X1   g594(.A1(new_n269), .A2(new_n272), .A3(new_n273), .A4(new_n264), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n322), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n304), .A2(new_n310), .A3(new_n305), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n310), .B1(new_n304), .B2(new_n305), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n306), .A2(new_n803), .A3(new_n307), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n318), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n798), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n320), .B1(new_n801), .B2(new_n803), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(KEYINPUT55), .C1(new_n801), .C2(new_n800), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n321), .A3(new_n808), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n797), .A2(KEYINPUT119), .B1(new_n276), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n270), .A2(new_n275), .B1(new_n205), .B2(new_n793), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n322), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n649), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n809), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n812), .A3(KEYINPUT118), .A4(new_n648), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n648), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n809), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n814), .A2(new_n820), .A3(KEYINPUT120), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n695), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n322), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n651), .A2(new_n826), .A3(new_n276), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n788), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n607), .A2(new_n610), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n351), .A3(new_n733), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n552), .A3(new_n602), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n276), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1340gat));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n353), .A3(new_n322), .ZN(new_n835));
  OAI21_X1  g634(.A(G120gat), .B1(new_n832), .B2(new_n826), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1341gat));
  AOI21_X1  g636(.A(G127gat), .B1(new_n830), .B2(new_n634), .ZN(new_n838));
  INV_X1    g637(.A(G127gat), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n832), .A2(new_n839), .A3(new_n695), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n838), .A2(new_n840), .ZN(G1342gat));
  NAND2_X1  g640(.A1(new_n828), .A2(new_n829), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(G134gat), .A3(new_n649), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  OAI21_X1  g645(.A(G134gat), .B1(new_n832), .B2(new_n649), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  NOR2_X1   g647(.A1(new_n713), .A2(new_n788), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n825), .A2(new_n827), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n554), .ZN(new_n852));
  INV_X1    g651(.A(new_n827), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n797), .B1(new_n276), .B2(new_n809), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n649), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n634), .B1(new_n820), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(KEYINPUT57), .B(new_n554), .C1(new_n853), .C2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n733), .B(new_n849), .C1(new_n852), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G141gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n552), .B1(new_n825), .B2(new_n827), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n849), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n330), .A3(new_n733), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1344gat));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n328), .A3(new_n322), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n849), .B1(new_n852), .B2(new_n858), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n826), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n328), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n861), .A2(new_n850), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n855), .B1(new_n809), .B2(new_n818), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n827), .B1(new_n877), .B2(new_n634), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n878), .B2(new_n554), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n322), .A3(new_n849), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n871), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n870), .B1(new_n874), .B2(new_n883), .ZN(G1345gat));
  NOR3_X1   g683(.A1(new_n872), .A2(new_n335), .A3(new_n695), .ZN(new_n885));
  AOI21_X1  g684(.A(G155gat), .B1(new_n863), .B2(new_n634), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n872), .B2(new_n649), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n336), .A3(new_n648), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n556), .A2(new_n616), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n602), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT125), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(KEYINPUT125), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n851), .A2(new_n552), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n276), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n556), .B1(new_n825), .B2(new_n827), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n829), .A2(new_n515), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(KEYINPUT122), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n897), .A2(new_n903), .A3(new_n899), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n276), .A2(G169gat), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(KEYINPUT124), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT124), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n896), .B1(new_n907), .B2(new_n908), .ZN(G1348gat));
  NOR3_X1   g708(.A1(new_n895), .A2(new_n315), .A3(new_n826), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n322), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n315), .ZN(G1349gat));
  OAI21_X1  g711(.A(G183gat), .B1(new_n895), .B2(new_n695), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n439), .A2(new_n442), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n634), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n901), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n905), .A2(new_n648), .A3(new_n425), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n895), .A2(new_n649), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(G190gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n919), .B2(G190gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(G1351gat));
  NOR2_X1   g722(.A1(new_n616), .A2(new_n552), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n897), .A2(new_n595), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(G197gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n733), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n595), .A2(new_n891), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n875), .B2(new_n880), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n733), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n926), .ZN(G1352gat));
  NOR2_X1   g730(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n826), .A2(G204gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g733(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  AOI211_X1 g736(.A(new_n826), .B(new_n928), .C1(new_n875), .C2(new_n880), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n936), .B(new_n937), .C1(new_n317), .C2(new_n938), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n925), .A2(new_n408), .A3(new_n634), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n929), .A2(new_n634), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n943));
  AOI211_X1 g742(.A(new_n943), .B(new_n408), .C1(new_n929), .C2(new_n634), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n942), .B2(new_n944), .ZN(G1354gat));
  NAND3_X1  g744(.A1(new_n929), .A2(G218gat), .A3(new_n648), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n897), .A2(new_n595), .A3(new_n924), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n409), .B1(new_n947), .B2(new_n649), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1355gat));
endmodule


