//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT65), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n211), .B(new_n212), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n207), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(G58), .A2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n228), .A2(G50), .A3(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n210), .B(new_n222), .C1(new_n225), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  XNOR2_X1  g0049(.A(KEYINPUT73), .B(G200), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT68), .B(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n258), .B1(G226), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n260), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G222), .A2(G1698), .ZN(new_n273));
  XOR2_X1   g0073(.A(KEYINPUT69), .B(G223), .Z(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(G1698), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n251), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n265), .A2(new_n276), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(G190), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n280), .A2(new_n224), .A3(G1), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n223), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n261), .B2(G20), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n286), .B2(G50), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g0088(.A(KEYINPUT8), .B(G58), .Z(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n269), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G150), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n204), .A2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n295), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n291), .B2(new_n293), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT71), .B1(new_n306), .B2(new_n301), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n288), .B1(new_n308), .B2(new_n285), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n279), .B1(new_n309), .B2(KEYINPUT9), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  AOI211_X1 g0111(.A(new_n311), .B(new_n288), .C1(new_n308), .C2(new_n285), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n308), .A2(new_n285), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n311), .B1(new_n314), .B2(new_n288), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(new_n279), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n278), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G169), .B2(new_n278), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n309), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n281), .A2(new_n203), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n295), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n201), .B2(new_n299), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n330));
  INV_X1    g0130(.A(new_n286), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n327), .B(new_n330), .C1(new_n203), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT11), .B1(new_n329), .B2(new_n285), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G238), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n257), .B1(new_n263), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT3), .B(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n214), .A2(G1698), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n339), .C1(G226), .C2(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n260), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT13), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n347));
  NOR2_X1   g0147(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n343), .B(new_n350), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n346), .A2(new_n349), .B1(new_n320), .B2(new_n351), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n335), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n334), .B1(new_n344), .B2(new_n355), .C1(new_n356), .C2(new_n351), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n202), .A2(new_n203), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n226), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n298), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n338), .B2(G20), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n366), .B2(G68), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n285), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT76), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(new_n267), .A3(G33), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT76), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n224), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n203), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n363), .A3(new_n224), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n362), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT77), .B1(new_n379), .B2(KEYINPUT16), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n269), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n371), .B1(new_n267), .B2(G33), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n268), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT7), .B1(new_n383), .B2(G20), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(G68), .A3(new_n378), .ZN(new_n385));
  INV_X1    g0185(.A(new_n362), .ZN(new_n386));
  AND4_X1   g0186(.A1(KEYINPUT77), .A2(new_n385), .A3(KEYINPUT16), .A4(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n370), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n294), .A2(new_n281), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n331), .B2(new_n294), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n257), .B1(new_n263), .B2(new_n214), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  MUX2_X1   g0193(.A(G223), .B(G226), .S(G1698), .Z(new_n394));
  AOI22_X1  g0194(.A1(new_n383), .A2(new_n394), .B1(G33), .B2(G87), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(G190), .C1(new_n260), .C2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n260), .ZN(new_n397));
  OAI21_X1  g0197(.A(G200), .B1(new_n397), .B2(new_n392), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n388), .A2(new_n391), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT17), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n388), .A2(new_n402), .A3(new_n391), .A4(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n393), .B1(new_n260), .B2(new_n395), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G169), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n320), .B2(new_n405), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n382), .A2(new_n268), .ZN(new_n408));
  AOI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n372), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n409), .B2(new_n363), .ZN(new_n410));
  INV_X1    g0210(.A(new_n378), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT16), .B(new_n386), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT77), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n385), .A2(KEYINPUT77), .A3(KEYINPUT16), .A4(new_n386), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n369), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n407), .B1(new_n416), .B2(new_n390), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n407), .B(KEYINPUT18), .C1(new_n416), .C2(new_n390), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n404), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n285), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n292), .A2(new_n299), .B1(new_n224), .B2(new_n266), .ZN(new_n424));
  XOR2_X1   g0224(.A(KEYINPUT15), .B(G87), .Z(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n295), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(KEYINPUT72), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n426), .A2(KEYINPUT72), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n281), .A2(new_n266), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n331), .B2(new_n266), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n258), .B1(G244), .B2(new_n264), .ZN(new_n434));
  NOR2_X1   g0234(.A1(G232), .A2(G1698), .ZN(new_n435));
  INV_X1    g0235(.A(G1698), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(G238), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n338), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n259), .C1(G107), .C2(new_n338), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n250), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n433), .B(new_n441), .C1(new_n356), .C2(new_n440), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n345), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n432), .B(new_n443), .C1(G179), .C2(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR4_X1   g0245(.A1(new_n325), .A2(new_n358), .A3(new_n422), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n253), .A2(G1), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n252), .B2(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT80), .ZN(new_n450));
  INV_X1    g0250(.A(G41), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT5), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT80), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n448), .C1(new_n252), .C2(KEYINPUT5), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n259), .A2(new_n255), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n450), .A2(new_n452), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n216), .A2(new_n436), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G264), .B2(new_n436), .ZN(new_n458));
  INV_X1    g0258(.A(G303), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n375), .A2(new_n458), .B1(new_n459), .B2(new_n338), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n259), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n449), .A2(KEYINPUT80), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n454), .A2(new_n452), .ZN(new_n464));
  OAI211_X1 g0264(.A(G270), .B(new_n260), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(G190), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n281), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n282), .B(new_n423), .C1(G1), .C2(new_n269), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n467), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n224), .C1(G33), .C2(new_n215), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(new_n285), .C1(new_n224), .C2(G116), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT20), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n474), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n476), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n470), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n466), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n355), .B1(new_n462), .B2(new_n465), .ZN(new_n483));
  OR3_X1    g0283(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT85), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n383), .A2(KEYINPUT22), .A3(new_n224), .A4(G87), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT22), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n224), .A2(G87), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n271), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n269), .A2(new_n467), .A3(G20), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n224), .B2(G107), .ZN(new_n493));
  INV_X1    g0293(.A(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT23), .A3(G20), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n487), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n487), .A2(KEYINPUT24), .A3(new_n490), .A4(new_n496), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n285), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n282), .A2(G107), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT25), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n469), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G264), .B(new_n260), .C1(new_n463), .C2(new_n464), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n216), .A2(G1698), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(G250), .B2(G1698), .ZN(new_n510));
  INV_X1    g0310(.A(G294), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n375), .A2(new_n510), .B1(new_n269), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n259), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n508), .A2(new_n320), .A3(new_n456), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n456), .A3(new_n513), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n345), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G250), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n259), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n448), .A2(KEYINPUT81), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n253), .B2(G1), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(KEYINPUT82), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n522), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n269), .A2(new_n451), .ZN(new_n526));
  OAI21_X1  g0326(.A(G250), .B1(new_n526), .B2(new_n223), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n523), .A2(new_n528), .B1(G45), .B2(new_n256), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n336), .A2(new_n436), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G244), .B2(new_n436), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n375), .A2(new_n531), .B1(new_n269), .B2(new_n467), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n259), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G169), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n529), .A2(G179), .A3(new_n533), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n383), .A2(new_n224), .A3(G68), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT19), .B1(new_n295), .B2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(G87), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n215), .A3(new_n494), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n224), .B1(new_n341), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n539), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n285), .ZN(new_n546));
  INV_X1    g0346(.A(new_n425), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n281), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n505), .A2(new_n425), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n546), .A2(KEYINPUT83), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT83), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n537), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n515), .A2(G200), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n508), .A2(G190), .A3(new_n456), .A4(new_n513), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(new_n501), .A3(new_n506), .A4(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n251), .B1(new_n529), .B2(new_n533), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n505), .A2(G87), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n546), .A2(new_n560), .A3(new_n548), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n559), .B(new_n562), .C1(new_n356), .C2(new_n534), .ZN(new_n563));
  AND4_X1   g0363(.A1(new_n517), .A2(new_n554), .A3(new_n557), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n298), .A2(G77), .ZN(new_n565));
  XNOR2_X1  g0365(.A(G97), .B(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT6), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n215), .A2(KEYINPUT6), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n566), .B1(new_n567), .B2(KEYINPUT6), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n565), .B1(new_n571), .B2(new_n224), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n494), .B1(new_n364), .B2(new_n365), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n285), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n282), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n505), .B2(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(new_n260), .C1(new_n463), .C2(new_n464), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n338), .A2(KEYINPUT4), .A3(G244), .A4(new_n436), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n338), .B2(G250), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n471), .B(new_n579), .C1(new_n581), .C2(new_n436), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT4), .B1(new_n383), .B2(G244), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n259), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n578), .A2(new_n584), .A3(new_n456), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(G200), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n578), .A2(new_n584), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G190), .A3(new_n456), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n320), .A3(new_n456), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n574), .A2(new_n576), .B1(new_n585), .B2(new_n345), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n586), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n462), .A2(new_n465), .ZN(new_n592));
  INV_X1    g0392(.A(new_n470), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n477), .A2(new_n476), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n474), .B2(new_n473), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n595), .B2(new_n479), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(new_n596), .A3(G169), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n592), .A2(new_n596), .A3(KEYINPUT21), .A4(G169), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(G179), .A3(new_n465), .A4(new_n462), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n486), .A2(new_n564), .A3(new_n591), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n447), .A2(new_n603), .ZN(G372));
  NAND2_X1  g0404(.A1(new_n354), .A2(new_n444), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n404), .A3(new_n357), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n421), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT88), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n606), .A2(KEYINPUT88), .A3(new_n421), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n319), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n534), .A2(new_n356), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n612), .A2(new_n561), .A3(new_n558), .ZN(new_n613));
  INV_X1    g0413(.A(new_n551), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n537), .B2(KEYINPUT86), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT86), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n535), .A2(new_n616), .A3(new_n536), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n613), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n590), .A2(new_n589), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n617), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n554), .A2(new_n589), .A3(new_n563), .A4(new_n590), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n517), .A2(KEYINPUT87), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n507), .A2(new_n516), .A3(new_n629), .A4(new_n514), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n602), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n623), .A2(new_n557), .A3(new_n563), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n632), .A3(new_n591), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n446), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n611), .A2(new_n324), .A3(new_n635), .ZN(G369));
  AND2_X1   g0436(.A1(new_n600), .A2(new_n601), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n599), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n485), .B2(new_n484), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n280), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n261), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n481), .A2(new_n647), .ZN(new_n648));
  MUX2_X1   g0448(.A(new_n639), .B(new_n638), .S(new_n648), .Z(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n517), .A2(new_n557), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n507), .A2(new_n646), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n517), .A2(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n646), .B1(new_n628), .B2(new_n630), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n602), .A2(new_n646), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n252), .ZN(new_n662));
  INV_X1    g0462(.A(new_n208), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n541), .A2(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n230), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n619), .B1(new_n618), .B2(new_n621), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n623), .B1(new_n624), .B2(KEYINPUT26), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n637), .A2(new_n599), .A3(new_n517), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n632), .A2(new_n591), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n646), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT29), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n646), .B1(new_n627), .B2(new_n633), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(KEYINPUT29), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n515), .A2(new_n534), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n587), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n462), .A2(G179), .A3(new_n465), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n682), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n680), .A3(KEYINPUT30), .A4(new_n587), .ZN(new_n685));
  AOI21_X1  g0485(.A(G179), .B1(new_n529), .B2(new_n533), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n592), .A2(new_n585), .A3(new_n515), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n646), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI221_X1 g0493(.A(new_n691), .B1(new_n689), .B2(new_n693), .C1(new_n603), .C2(new_n646), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n678), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n669), .B1(new_n697), .B2(G1), .ZN(G364));
  AOI21_X1  g0498(.A(new_n261), .B1(new_n640), .B2(G45), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n664), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n651), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(G330), .B2(new_n649), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n223), .B1(G20), .B2(new_n345), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G283), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n224), .A2(G190), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n251), .A2(G179), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n224), .A2(new_n356), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n251), .A2(G179), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n706), .A2(new_n710), .B1(new_n714), .B2(new_n459), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G179), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT94), .Z(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(G329), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n320), .A2(new_n355), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n711), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n320), .A2(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n711), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(G326), .A2(new_n723), .B1(new_n726), .B2(G322), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(new_n707), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT33), .B(G317), .Z(new_n729));
  OAI211_X1 g0529(.A(new_n727), .B(new_n271), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n707), .A2(new_n724), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT91), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n730), .B1(G311), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n224), .B1(new_n716), .B2(G190), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n720), .B(new_n738), .C1(new_n511), .C2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n717), .ZN(new_n744));
  XOR2_X1   g0544(.A(KEYINPUT92), .B(G159), .Z(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT32), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n338), .B1(new_n725), .B2(new_n202), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n722), .A2(new_n201), .B1(new_n728), .B2(new_n203), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n714), .A2(new_n540), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(G77), .B2(new_n737), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n709), .A2(G107), .ZN(new_n753));
  INV_X1    g0553(.A(new_n742), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G97), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n750), .A2(new_n752), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n705), .B1(new_n743), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n704), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n245), .A2(G45), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n383), .A2(new_n663), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n763), .B(new_n764), .C1(G45), .C2(new_n230), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n338), .A2(new_n208), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(KEYINPUT90), .B2(G355), .ZN(new_n767));
  OR2_X1    g0567(.A1(G355), .A2(KEYINPUT90), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n767), .A2(new_n768), .B1(new_n467), .B2(new_n663), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n762), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n757), .A2(new_n770), .A3(new_n664), .A4(new_n700), .ZN(new_n771));
  INV_X1    g0571(.A(new_n760), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n649), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n703), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(G396));
  XOR2_X1   g0575(.A(new_n444), .B(KEYINPUT96), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n442), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n631), .A2(new_n591), .A3(new_n632), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n647), .B(new_n778), .C1(new_n779), .C2(new_n626), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n433), .A2(new_n647), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n781), .B1(new_n444), .B2(new_n647), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n780), .B1(new_n677), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT97), .ZN(new_n784));
  OR3_X1    g0584(.A1(new_n783), .A2(new_n784), .A3(new_n695), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n783), .B2(new_n695), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n701), .B1(new_n783), .B2(new_n695), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n705), .A2(new_n759), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n701), .B1(G77), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n718), .A2(new_n791), .B1(new_n714), .B2(new_n494), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n722), .A2(new_n459), .B1(new_n728), .B2(new_n706), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n338), .B(new_n793), .C1(G294), .C2(new_n726), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n794), .B(new_n755), .C1(new_n540), .C2(new_n710), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n792), .B(new_n795), .C1(G116), .C2(new_n737), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT95), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT95), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G137), .A2(new_n723), .B1(new_n726), .B2(G143), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n300), .B2(new_n728), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n737), .B2(new_n745), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT34), .Z(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n718), .A2(new_n803), .B1(new_n714), .B2(new_n201), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n375), .B(new_n804), .C1(G68), .C2(new_n709), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(new_n202), .C2(new_n742), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n797), .A2(new_n798), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n790), .B1(new_n807), .B2(new_n704), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n782), .B2(new_n759), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n788), .A2(new_n809), .ZN(G384));
  AOI21_X1  g0610(.A(new_n693), .B1(new_n688), .B2(new_n646), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n603), .B2(new_n646), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n688), .A2(new_n690), .A3(new_n646), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n335), .A2(new_n646), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT98), .Z(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n358), .A2(new_n817), .B1(new_n354), .B2(new_n647), .ZN(new_n818));
  AND4_X1   g0618(.A1(KEYINPUT40), .A2(new_n814), .A3(new_n782), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT99), .ZN(new_n820));
  INV_X1    g0620(.A(new_n644), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n416), .B2(new_n390), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n400), .A2(new_n417), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT37), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n400), .A2(new_n417), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n820), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n822), .B1(new_n404), .B2(new_n421), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n824), .A2(new_n820), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT38), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g0631(.A1(new_n825), .A2(new_n400), .A3(new_n417), .A4(new_n822), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n285), .B1(new_n379), .B2(new_n368), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n414), .B2(new_n415), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n821), .B1(new_n834), .B2(new_n390), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n407), .B1(new_n834), .B2(new_n390), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(new_n400), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n832), .B1(KEYINPUT37), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n835), .B1(new_n404), .B2(new_n421), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n831), .A2(KEYINPUT102), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT102), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n824), .A2(new_n826), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT99), .ZN(new_n845));
  INV_X1    g0645(.A(new_n822), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n422), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n830), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n840), .ZN(new_n849));
  INV_X1    g0649(.A(new_n835), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n422), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n837), .A2(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n826), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n843), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n819), .B1(new_n842), .B2(new_n855), .ZN(new_n856));
  AND4_X1   g0656(.A1(new_n782), .A2(new_n812), .A3(new_n818), .A4(new_n813), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n840), .B1(new_n838), .B2(new_n839), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n854), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT40), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n856), .A2(G330), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n814), .A2(G330), .A3(new_n446), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n814), .A2(new_n446), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT102), .B1(new_n831), .B2(new_n841), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n849), .A2(new_n843), .A3(new_n854), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n860), .B1(new_n868), .B2(new_n819), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n862), .A2(new_n863), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT101), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n676), .B(new_n446), .C1(KEYINPUT29), .C2(new_n677), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n872), .A2(new_n324), .A3(new_n611), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n871), .B(new_n873), .Z(new_n874));
  NOR2_X1   g0674(.A1(new_n421), .A2(new_n821), .ZN(new_n875));
  INV_X1    g0675(.A(new_n818), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n776), .A2(new_n646), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n780), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n875), .B1(new_n879), .B2(new_n859), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT100), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n824), .A2(new_n820), .A3(new_n826), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n883), .A2(new_n827), .A3(new_n828), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n882), .B(new_n854), .C1(new_n884), .C2(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n841), .B1(new_n840), .B2(new_n848), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT100), .B1(new_n888), .B2(new_n882), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n354), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n647), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n880), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n874), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n874), .A2(new_n893), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n894), .B(new_n895), .C1(new_n261), .C2(new_n640), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT35), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n571), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n571), .A2(new_n897), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n898), .A2(G116), .A3(new_n225), .A4(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT36), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n230), .A2(new_n266), .A3(new_n359), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n203), .A2(G50), .ZN(new_n903));
  OAI211_X1 g0703(.A(G1), .B(new_n280), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n896), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT103), .ZN(G367));
  NOR2_X1   g0706(.A1(new_n562), .A2(new_n647), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n618), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n623), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT104), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n659), .A2(new_n652), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n577), .A2(new_n646), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n591), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT42), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n620), .B1(new_n916), .B2(new_n517), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n647), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n914), .A2(KEYINPUT42), .A3(new_n916), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n912), .B(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n657), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n916), .B1(new_n620), .B2(new_n647), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n923), .B(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n664), .B(KEYINPUT41), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n914), .B1(new_n656), .B2(new_n659), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n924), .B1(new_n650), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n660), .A2(new_n925), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT45), .Z(new_n933));
  NOR2_X1   g0733(.A1(new_n660), .A2(new_n925), .ZN(new_n934));
  OR2_X1    g0734(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n934), .B2(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n933), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n931), .A2(new_n939), .A3(new_n697), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n929), .B1(new_n940), .B2(new_n697), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n927), .B1(new_n941), .B2(new_n700), .ZN(new_n942));
  INV_X1    g0742(.A(new_n764), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n761), .B1(new_n208), .B2(new_n547), .C1(new_n240), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n701), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n726), .A2(G150), .ZN(new_n946));
  XOR2_X1   g0746(.A(KEYINPUT107), .B(G137), .Z(new_n947));
  INV_X1    g0747(.A(G143), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n946), .B1(new_n947), .B2(new_n717), .C1(new_n948), .C2(new_n722), .ZN(new_n949));
  INV_X1    g0749(.A(new_n728), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n271), .B(new_n949), .C1(new_n950), .C2(new_n745), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n713), .A2(G58), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n737), .A2(G50), .B1(G77), .B2(new_n709), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n742), .A2(new_n203), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n736), .A2(new_n706), .B1(new_n710), .B2(new_n215), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G311), .A2(new_n723), .B1(new_n726), .B2(G303), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n717), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n957), .A2(new_n383), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n714), .A2(new_n467), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n962), .A2(KEYINPUT46), .B1(new_n511), .B2(new_n728), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT46), .B2(new_n962), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT106), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n961), .B1(new_n494), .B2(new_n742), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n964), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(KEYINPUT106), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n956), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT47), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n705), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n945), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n910), .B2(new_n772), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n942), .A2(new_n974), .ZN(G387));
  NAND3_X1  g0775(.A1(new_n654), .A2(new_n655), .A3(new_n760), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n764), .B1(new_n236), .B2(new_n253), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n666), .B2(new_n766), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n289), .A2(new_n201), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n981));
  AOI21_X1  g0781(.A(G45), .B1(G68), .B2(G77), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n980), .A2(new_n666), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n978), .A2(new_n983), .B1(new_n494), .B2(new_n663), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n701), .B1(new_n984), .B2(new_n762), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n714), .A2(new_n266), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n294), .B2(new_n950), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n737), .A2(G68), .B1(G97), .B2(new_n709), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n754), .A2(new_n425), .ZN(new_n989));
  INV_X1    g0789(.A(G159), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n722), .A2(new_n990), .B1(new_n725), .B2(new_n201), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n375), .B(new_n991), .C1(G150), .C2(new_n744), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(KEYINPUT108), .B(G322), .Z(new_n994));
  AOI22_X1  g0794(.A1(new_n723), .A2(new_n994), .B1(new_n726), .B2(G317), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n791), .B2(new_n728), .C1(new_n736), .C2(new_n459), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT48), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n706), .B2(new_n742), .C1(new_n511), .C2(new_n714), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n383), .B1(G326), .B2(new_n744), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n710), .B2(new_n467), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n993), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n985), .B1(new_n1003), .B2(new_n704), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n931), .A2(new_n700), .B1(new_n976), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n931), .A2(new_n697), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n664), .B(KEYINPUT110), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n931), .A2(new_n697), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(G393));
  OR3_X1    g0810(.A1(new_n939), .A2(new_n924), .A3(KEYINPUT111), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT111), .B1(new_n939), .B2(new_n924), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n939), .A2(new_n924), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n699), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n925), .A2(new_n772), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n761), .B1(new_n215), .B2(new_n208), .C1(new_n943), .C2(new_n248), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n701), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT51), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n722), .A2(new_n300), .B1(new_n725), .B2(new_n990), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n737), .A2(new_n289), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n1019), .B2(new_n1020), .C1(new_n203), .C2(new_n714), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n728), .A2(new_n201), .B1(new_n717), .B2(new_n948), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n375), .B(new_n1023), .C1(G87), .C2(new_n709), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n266), .B2(new_n742), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n737), .A2(G294), .B1(G283), .B2(new_n713), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n728), .A2(new_n459), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n338), .B(new_n1027), .C1(new_n744), .C2(new_n994), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n753), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n722), .A2(new_n959), .B1(new_n725), .B2(new_n791), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT52), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n467), .B2(new_n742), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1022), .A2(new_n1025), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1018), .B1(new_n1033), .B2(new_n704), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1015), .B1(new_n1016), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1014), .A2(new_n1006), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(new_n940), .A3(new_n1007), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(G390));
  OAI21_X1  g0838(.A(new_n701), .B1(new_n294), .B2(new_n789), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n338), .B1(new_n950), .B2(G107), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n467), .B2(new_n725), .C1(new_n706), .C2(new_n722), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n751), .B(new_n1041), .C1(G97), .C2(new_n737), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n718), .A2(new_n511), .B1(new_n710), .B2(new_n203), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT116), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n266), .C2(new_n742), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT54), .B(G143), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n736), .A2(new_n1047), .B1(new_n728), .B2(new_n947), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G159), .B2(new_n754), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  NAND2_X1  g0850(.A1(new_n713), .A2(G150), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT53), .Z(new_n1052));
  AOI22_X1  g0852(.A1(G128), .A2(new_n723), .B1(new_n726), .B2(G132), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n719), .A2(G125), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n271), .B1(new_n709), .B2(G50), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1045), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1039), .B1(new_n1058), .B2(new_n704), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n885), .A2(new_n881), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n882), .B1(new_n858), .B2(new_n854), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n888), .B2(new_n882), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1062), .B2(new_n881), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1059), .B1(new_n1063), .B2(new_n759), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n877), .B1(new_n677), .B2(new_n778), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n892), .B1(new_n1066), .B2(new_n876), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1060), .B(new_n1067), .C1(new_n1062), .C2(new_n881), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n877), .B1(new_n675), .B2(new_n778), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(new_n876), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n892), .B(KEYINPUT112), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n868), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n694), .A2(G330), .A3(new_n782), .A4(new_n818), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1068), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1071), .B1(new_n1069), .B2(new_n876), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n866), .B2(new_n867), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n890), .B2(new_n1067), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n857), .A2(G330), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1074), .B(new_n700), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1065), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AND4_X1   g0881(.A1(new_n324), .A2(new_n872), .A3(new_n611), .A4(new_n863), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n694), .A2(G330), .A3(new_n782), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n876), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1066), .B1(new_n1084), .B2(new_n1078), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n812), .A2(new_n782), .A3(G330), .A4(new_n813), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n876), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n1073), .A3(new_n1069), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1082), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT113), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n1074), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n1007), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n1091), .A3(new_n1090), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1081), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G378));
  NOR2_X1   g0898(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1074), .B(new_n1100), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1082), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT118), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n325), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n309), .A2(new_n644), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n319), .A2(KEYINPUT118), .A3(new_n324), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT118), .B1(new_n319), .B2(new_n324), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1103), .B(new_n323), .C1(new_n313), .C2(new_n318), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n862), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n880), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n892), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1063), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1115), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n869), .A2(G330), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n869), .B2(G330), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n814), .A2(KEYINPUT40), .A3(new_n782), .A4(new_n818), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n866), .B2(new_n867), .ZN(new_n1125));
  INV_X1    g0925(.A(G330), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n1125), .A2(new_n860), .A3(new_n1115), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n893), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1102), .A2(KEYINPUT57), .A3(new_n1122), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT119), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1123), .A2(new_n893), .A3(new_n1127), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1119), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(KEYINPUT57), .A4(new_n1102), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT57), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1101), .A2(new_n1082), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1128), .A2(new_n1122), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1130), .A2(new_n1007), .A3(new_n1135), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1133), .A2(new_n700), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n701), .B1(G50), .B2(new_n789), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n710), .A2(new_n202), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1143), .A2(new_n383), .A3(new_n662), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n706), .B2(new_n718), .C1(new_n547), .C2(new_n736), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G97), .A2(new_n950), .B1(new_n726), .B2(G107), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n467), .B2(new_n722), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1145), .A2(new_n954), .A3(new_n986), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n201), .B1(G33), .B2(G41), .C1(new_n383), .C2(new_n662), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G128), .A2(new_n726), .B1(new_n950), .B2(G132), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n722), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G137), .B2(new_n737), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n300), .B2(new_n742), .C1(new_n714), .C2(new_n1047), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n709), .A2(new_n745), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n744), .C2(G124), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1151), .B1(KEYINPUT58), .B2(new_n1148), .C1(new_n1157), .C2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1142), .B1(new_n1162), .B2(new_n704), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1115), .B2(new_n759), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1141), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1140), .A2(new_n1165), .ZN(G375));
  INV_X1    g0966(.A(new_n1082), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1099), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n928), .A3(new_n1090), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n718), .A2(new_n459), .B1(new_n714), .B2(new_n215), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n725), .A2(new_n706), .B1(new_n728), .B2(new_n467), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n338), .B(new_n1171), .C1(G294), .C2(new_n723), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1172), .B(new_n989), .C1(new_n266), .C2(new_n710), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1170), .B(new_n1173), .C1(G107), .C2(new_n737), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n375), .B(new_n1143), .C1(new_n754), .C2(G50), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n719), .A2(G128), .B1(G159), .B2(new_n713), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n300), .C2(new_n736), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT120), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n950), .A2(new_n1046), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n803), .B2(new_n722), .C1(new_n725), .C2(new_n947), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1177), .B2(KEYINPUT120), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1174), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n701), .B1(G68), .B2(new_n789), .C1(new_n1182), .C2(new_n705), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n876), .B2(new_n758), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1100), .B2(new_n700), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1169), .A2(new_n1185), .ZN(G381));
  NAND3_X1  g0986(.A1(new_n1140), .A2(new_n1097), .A3(new_n1165), .ZN(new_n1187));
  OR4_X1    g0987(.A1(G396), .A2(G387), .A3(G384), .A4(G393), .ZN(new_n1188));
  OR4_X1    g0988(.A1(G390), .A2(new_n1187), .A3(G381), .A4(new_n1188), .ZN(G407));
  OAI211_X1 g0989(.A(G407), .B(G213), .C1(G343), .C2(new_n1187), .ZN(G409));
  XOR2_X1   g0990(.A(G390), .B(G387), .Z(new_n1191));
  XNOR2_X1  g0991(.A(G393), .B(new_n774), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1191), .A2(KEYINPUT127), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1191), .B2(KEYINPUT127), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1140), .A2(G378), .A3(new_n1165), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT121), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT121), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1128), .A2(new_n1122), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n700), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1133), .A2(new_n928), .A3(new_n1102), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n1164), .A3(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1204), .A2(KEYINPUT122), .A3(new_n1097), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT122), .B1(new_n1204), .B2(new_n1097), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1198), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT123), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1168), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1099), .A2(new_n1167), .A3(KEYINPUT60), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1211), .A2(new_n1007), .A3(new_n1090), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1185), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT124), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G384), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n788), .A2(KEYINPUT124), .A3(new_n809), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1214), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1213), .A2(new_n1185), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT125), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1221), .B(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1198), .B(KEYINPUT123), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n645), .A2(G213), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1209), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT62), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1207), .A2(new_n1225), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n645), .A2(G213), .A3(G2897), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1221), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT61), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1207), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT62), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1197), .B1(new_n1227), .B2(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1237));
  NAND2_X1  g1037(.A1(new_n1226), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1209), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1231), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1207), .A2(KEYINPUT63), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1194), .A2(new_n1195), .A3(KEYINPUT61), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1236), .A2(new_n1243), .ZN(G405));
  XNOR2_X1  g1044(.A(G375), .B(G378), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(new_n1223), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1221), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1196), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1197), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(G402));
endmodule


