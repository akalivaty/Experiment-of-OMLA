//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n651, new_n653, new_n654,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  AOI22_X1  g031(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n462), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n471), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n469), .A2(G137), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND4_X1  g052(.A1(new_n472), .A2(new_n468), .A3(G2105), .A4(new_n465), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n470), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n478), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n472), .A2(new_n468), .A3(new_n470), .A4(new_n465), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(G136), .B2(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n472), .A2(new_n468), .A3(new_n487), .A4(new_n465), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n486), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(G114), .B2(new_n470), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n478), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n491), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(G62), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(G50), .A2(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n510), .B2(G88), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n503), .A2(new_n504), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n506), .A2(new_n515), .ZN(G166));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(KEYINPUT71), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n512), .B2(new_n513), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n519), .A2(new_n521), .A3(G543), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT72), .B(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n499), .A2(new_n500), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  OR3_X1    g101(.A1(new_n525), .A2(KEYINPUT70), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT70), .B1(new_n525), .B2(new_n526), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n524), .A2(new_n529), .A3(KEYINPUT73), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n525), .A2(new_n514), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n533), .B1(G89), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT73), .B1(new_n524), .B2(new_n529), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n498), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n522), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(G90), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  OAI21_X1  g119(.A(G56), .B1(new_n499), .B2(new_n500), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n498), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n519), .A2(new_n521), .A3(G543), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n508), .B2(new_n509), .ZN(new_n553));
  INV_X1    g128(.A(new_n546), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n548), .B(G651), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n517), .A2(new_n518), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n510), .A2(new_n556), .A3(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT76), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND3_X1  g140(.A1(new_n510), .A2(new_n556), .A3(G91), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(G65), .B1(new_n499), .B2(new_n500), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n498), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n519), .A2(new_n521), .A3(G53), .A4(G543), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n524), .A2(new_n529), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n578), .A2(new_n530), .A3(new_n535), .ZN(G286));
  OR2_X1    g154(.A1(new_n506), .A2(new_n515), .ZN(G303));
  NAND2_X1  g155(.A1(new_n522), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT77), .B1(new_n534), .B2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n510), .A2(new_n556), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n587), .ZN(G288));
  OAI21_X1  g163(.A(G61), .B1(new_n499), .B2(new_n500), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(KEYINPUT78), .A3(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n534), .A2(G86), .ZN(new_n598));
  AND2_X1   g173(.A1(G48), .A2(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n556), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT78), .B1(new_n591), .B2(G651), .ZN(new_n602));
  AOI211_X1 g177(.A(new_n593), .B(new_n498), .C1(new_n589), .C2(new_n590), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n598), .B(new_n600), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(G72), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G60), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n525), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n534), .A2(G85), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n519), .A2(new_n521), .A3(G47), .A4(G543), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n612), .A2(KEYINPUT80), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(KEYINPUT80), .B1(new_n612), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n611), .B1(new_n615), .B2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n549), .A2(KEYINPUT81), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n549), .A2(KEYINPUT81), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n619), .A2(G54), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n584), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n510), .A2(G66), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT82), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n630), .A2(G79), .A3(G543), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT83), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G66), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n632), .B(KEYINPUT83), .C1(new_n525), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G651), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n626), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n621), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n618), .B1(new_n638), .B2(G868), .ZN(G284));
  OAI21_X1  g214(.A(new_n618), .B1(new_n638), .B2(G868), .ZN(G321));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  NOR2_X1   g216(.A1(G286), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n568), .A2(new_n569), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n566), .B1(new_n643), .B2(new_n498), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n642), .B1(new_n641), .B2(new_n648), .ZN(G297));
  AOI21_X1  g224(.A(new_n642), .B1(new_n641), .B2(new_n648), .ZN(G280));
  INV_X1    g225(.A(G559), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n638), .B1(new_n651), .B2(G860), .ZN(G148));
  NAND2_X1  g227(.A1(new_n638), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G868), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g230(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n656));
  XNOR2_X1  g231(.A(G323), .B(new_n656), .ZN(G282));
  NAND2_X1  g232(.A1(new_n489), .A2(new_n474), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT12), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT13), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n484), .A2(G135), .ZN(new_n662));
  INV_X1    g237(.A(G123), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n470), .A2(G111), .ZN(new_n664));
  OAI21_X1  g239(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n665));
  OAI22_X1  g240(.A1(new_n478), .A2(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(G2096), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(G2096), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n661), .A2(new_n669), .A3(new_n670), .ZN(G156));
  INV_X1    g246(.A(G14), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2427), .B(G2438), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2430), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT15), .B(G2435), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(KEYINPUT14), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2443), .B(G2446), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1341), .B(G1348), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n672), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n683), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n679), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n686), .A2(new_n690), .ZN(G401));
  XNOR2_X1  g266(.A(G2084), .B(G2090), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT87), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2067), .B(G2678), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n695), .A2(KEYINPUT17), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT18), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G2100), .ZN(new_n700));
  INV_X1    g275(.A(G2100), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n696), .A2(KEYINPUT18), .ZN(new_n704));
  XOR2_X1   g279(.A(G2072), .B(G2078), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2096), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n703), .A2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(G227));
  XNOR2_X1  g286(.A(G1991), .B(G1996), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G1961), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G1966), .ZN(new_n715));
  INV_X1    g290(.A(G1966), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G1961), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT89), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1956), .B(G2474), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(G1961), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n714), .A2(G1966), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n718), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT19), .ZN(new_n726));
  AND2_X1   g301(.A1(G1971), .A2(G1976), .ZN(new_n727));
  NOR2_X1   g302(.A1(G1971), .A2(G1976), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  INV_X1    g305(.A(G1976), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G1971), .A2(G1976), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n732), .A2(KEYINPUT19), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT90), .B1(new_n725), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n723), .B1(new_n721), .B2(new_n722), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n729), .A2(new_n734), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n739), .A2(new_n740), .A3(new_n720), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT20), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n737), .A2(new_n738), .A3(new_n719), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n720), .B1(new_n718), .B2(new_n724), .ZN(new_n747));
  OAI211_X1 g322(.A(KEYINPUT91), .B(new_n735), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n719), .B1(new_n737), .B2(new_n738), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n729), .A2(new_n734), .A3(KEYINPUT91), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n749), .B(new_n750), .C1(new_n725), .C2(new_n741), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n736), .A2(new_n742), .A3(KEYINPUT20), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n745), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n745), .A2(new_n752), .A3(KEYINPUT92), .A4(new_n753), .ZN(new_n757));
  XNOR2_X1  g332(.A(G1981), .B(G1986), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n756), .B2(new_n757), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n762), .ZN(new_n764));
  INV_X1    g339(.A(new_n758), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n736), .A2(new_n742), .A3(KEYINPUT20), .ZN(new_n766));
  AOI21_X1  g341(.A(KEYINPUT20), .B1(new_n736), .B2(new_n742), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(KEYINPUT92), .B1(new_n768), .B2(new_n752), .ZN(new_n769));
  INV_X1    g344(.A(new_n757), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n764), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n713), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n771), .A2(new_n764), .A3(new_n772), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n775), .A2(new_n712), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(G229));
  INV_X1    g354(.A(G16), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n780), .ZN(new_n782));
  INV_X1    g357(.A(G2072), .ZN(new_n783));
  NOR2_X1   g358(.A1(G29), .A2(G33), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  INV_X1    g360(.A(G139), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n483), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n463), .A2(new_n465), .A3(G127), .ZN(new_n788));
  NAND2_X1  g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n470), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT25), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n787), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G29), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n785), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n782), .A2(G1961), .B1(new_n783), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT31), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(G11), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(G11), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n801), .A2(G28), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n795), .B1(new_n801), .B2(G28), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n799), .B(new_n800), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n667), .B2(G29), .ZN(new_n805));
  INV_X1    g380(.A(G2084), .ZN(new_n806));
  INV_X1    g381(.A(G34), .ZN(new_n807));
  AOI21_X1  g382(.A(G29), .B1(new_n807), .B2(KEYINPUT24), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(KEYINPUT24), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n476), .B2(new_n795), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n797), .B(new_n805), .C1(new_n806), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n795), .A2(G32), .ZN(new_n812));
  INV_X1    g387(.A(new_n478), .ZN(new_n813));
  NAND3_X1  g388(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT97), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n816), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT26), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT26), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n815), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  AOI22_X1  g396(.A1(G129), .A2(new_n813), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n474), .A2(G105), .ZN(new_n823));
  INV_X1    g398(.A(G141), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n483), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n812), .B1(new_n828), .B2(new_n795), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT27), .B(G1996), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n780), .A2(G19), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n559), .B2(new_n780), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1341), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n810), .A2(new_n806), .ZN(new_n835));
  OAI221_X1 g410(.A(new_n835), .B1(new_n796), .B2(new_n783), .C1(new_n782), .C2(G1961), .ZN(new_n836));
  NOR4_X1   g411(.A1(new_n811), .A2(new_n831), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(G4), .A2(G16), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n638), .B2(G16), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1348), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n795), .A2(G27), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G164), .B2(new_n795), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G2078), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n795), .A2(G26), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT28), .ZN(new_n845));
  INV_X1    g420(.A(G128), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n470), .A2(G116), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n478), .A2(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G140), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n483), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n845), .B1(new_n852), .B2(new_n795), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G2067), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n840), .A2(new_n843), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n837), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n795), .A2(G35), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT99), .Z(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(G162), .B2(new_n795), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT29), .Z(new_n860));
  INV_X1    g435(.A(G2090), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT100), .Z(new_n863));
  NOR2_X1   g438(.A1(G168), .A2(new_n780), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n780), .B2(G21), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT98), .B(G1966), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n780), .A2(G20), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT23), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n647), .B2(new_n780), .ZN(new_n870));
  INV_X1    g445(.A(G1956), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  OAI22_X1  g448(.A1(new_n865), .A2(new_n866), .B1(new_n860), .B2(new_n861), .ZN(new_n874));
  NOR4_X1   g449(.A1(new_n856), .A2(new_n863), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n606), .A2(G16), .ZN(new_n877));
  NOR2_X1   g452(.A1(G6), .A2(G16), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(KEYINPUT32), .B(G1981), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n883));
  INV_X1    g458(.A(new_n881), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n884), .A3(new_n879), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n780), .A2(G22), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(G166), .B2(new_n780), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n730), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n780), .A2(G23), .ZN(new_n890));
  INV_X1    g465(.A(G288), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(new_n780), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT33), .B(G1976), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n886), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT34), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n882), .A2(new_n885), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT95), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n612), .A2(new_n613), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT80), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n902), .A2(new_n614), .B1(G651), .B2(new_n610), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G16), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G16), .B2(G24), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n906), .A2(G1986), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(G1986), .ZN(new_n908));
  NOR2_X1   g483(.A1(G25), .A2(G29), .ZN(new_n909));
  OR2_X1    g484(.A1(G95), .A2(G2105), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n910), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n911));
  INV_X1    g486(.A(G119), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n478), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G131), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n483), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n909), .B1(new_n916), .B2(G29), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT35), .B(G1991), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT94), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n917), .B(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n907), .A2(new_n908), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n899), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n895), .A2(new_n898), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT34), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT36), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT36), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n876), .B1(new_n926), .B2(new_n928), .ZN(G311));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n922), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n875), .B1(new_n930), .B2(new_n931), .ZN(G150));
  NAND2_X1  g507(.A1(new_n638), .A2(G559), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT38), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n545), .A2(new_n546), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n548), .B1(new_n935), .B2(G651), .ZN(new_n936));
  AND4_X1   g511(.A1(G43), .A2(new_n519), .A3(new_n521), .A4(G543), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G67), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n508), .B2(new_n509), .ZN(new_n940));
  AND2_X1   g515(.A1(G80), .A2(G543), .ZN(new_n941));
  OAI21_X1  g516(.A(G651), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n519), .A2(new_n521), .A3(G55), .A4(G543), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n510), .A2(new_n556), .A3(G93), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n555), .A2(new_n557), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n938), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n551), .B2(new_n558), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n934), .B(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT39), .ZN(new_n952));
  AOI21_X1  g527(.A(G860), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n952), .B2(new_n951), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(G860), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT37), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(G145));
  INV_X1    g532(.A(KEYINPUT25), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n791), .B(new_n958), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n470), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n815), .A2(new_n820), .A3(new_n817), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n820), .B1(new_n815), .B2(new_n817), .ZN(new_n963));
  INV_X1    g538(.A(G129), .ZN(new_n964));
  OAI22_X1  g539(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n478), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n787), .A2(new_n961), .B1(new_n965), .B2(new_n825), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n793), .A2(new_n826), .A3(new_n822), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n469), .A2(G131), .A3(new_n470), .A4(new_n472), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n469), .A2(G119), .A3(G2105), .A4(new_n472), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT102), .A4(new_n911), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n913), .B2(new_n915), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n970), .A2(new_n972), .A3(new_n659), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n659), .B1(new_n970), .B2(new_n972), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n966), .B(new_n967), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n967), .A2(new_n966), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n970), .A2(new_n972), .ZN(new_n977));
  INV_X1    g552(.A(new_n659), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n970), .A2(new_n972), .A3(new_n659), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G164), .A2(new_n852), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n484), .A2(G142), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n813), .A2(G130), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n470), .A2(KEYINPUT101), .A3(G118), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT101), .B1(new_n470), .B2(G118), .ZN(new_n987));
  OR2_X1    g562(.A1(G106), .A2(G2105), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G2104), .A3(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n984), .B(new_n985), .C1(new_n986), .C2(new_n989), .ZN(new_n990));
  OAI22_X1  g565(.A1(new_n491), .A2(new_n496), .B1(new_n849), .B2(new_n851), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n983), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n983), .B2(new_n991), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n982), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n668), .A2(G160), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n667), .A2(new_n476), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n996), .A2(new_n997), .A3(G162), .ZN(new_n998));
  AOI21_X1  g573(.A(G162), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n992), .A2(new_n993), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(new_n975), .A3(new_n981), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n995), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT103), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n995), .A2(KEYINPUT103), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1000), .B1(new_n995), .B2(new_n1002), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G37), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g586(.A1(new_n948), .A2(G868), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G288), .B(G166), .ZN(new_n1013));
  NAND3_X1  g588(.A1(G290), .A2(new_n601), .A3(new_n605), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G290), .B1(new_n605), .B2(new_n601), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(G303), .B(G288), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n606), .A2(new_n903), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n1014), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT104), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1022), .B(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT106), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1022), .B(new_n1023), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n653), .B(new_n950), .Z(new_n1030));
  OAI21_X1  g605(.A(new_n647), .B1(new_n621), .B2(new_n637), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n636), .A2(new_n633), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n619), .A2(G54), .A3(new_n620), .ZN(new_n1033));
  NAND4_X1  g608(.A1(G299), .A2(new_n1032), .A3(new_n1033), .A4(new_n626), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT41), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1031), .A2(new_n1034), .A3(KEYINPUT41), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1037), .B1(new_n1030), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1026), .A2(new_n1029), .A3(new_n1042), .ZN(new_n1043));
  OR3_X1    g618(.A1(new_n1025), .A2(new_n1042), .A3(KEYINPUT106), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1012), .B1(new_n1045), .B2(G868), .ZN(G295));
  AOI21_X1  g621(.A(new_n1012), .B1(new_n1045), .B2(G868), .ZN(G331));
  AND3_X1   g622(.A1(new_n947), .A2(G301), .A3(new_n949), .ZN(new_n1048));
  AOI21_X1  g623(.A(G301), .B1(new_n947), .B2(new_n949), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1048), .A2(new_n1049), .A3(G286), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n945), .B1(new_n938), .B2(new_n946), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n551), .A2(new_n948), .A3(new_n558), .ZN(new_n1052));
  OAI21_X1  g627(.A(G171), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n947), .A2(new_n949), .A3(G301), .ZN(new_n1054));
  AOI21_X1  g629(.A(G168), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1035), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT108), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1021), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1041), .ZN(new_n1060));
  OAI21_X1  g635(.A(G286), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1053), .A2(G168), .A3(new_n1054), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT108), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n1035), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G37), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1036), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1069), .A2(new_n1064), .B1(new_n1059), .B2(new_n1041), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1058), .B1(new_n1070), .B2(new_n1057), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT43), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1040), .B(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT109), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT109), .B(KEYINPUT41), .C1(new_n1031), .C2(new_n1034), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1063), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1021), .B1(new_n1079), .B2(new_n1069), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT43), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n1067), .A4(new_n1066), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1072), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1080), .A2(new_n1067), .A3(new_n1066), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT44), .B1(new_n1086), .B2(new_n1081), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1068), .A2(new_n1071), .A3(KEYINPUT43), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(G397));
  INV_X1    g664(.A(new_n496), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n489), .A2(new_n490), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1384), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT111), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT45), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1094), .B2(KEYINPUT111), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n467), .A2(G40), .A3(new_n473), .A4(new_n475), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(G1996), .A3(new_n827), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1101), .A2(KEYINPUT114), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(KEYINPUT114), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1100), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n852), .B(G2067), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1996), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n828), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1102), .A2(new_n1103), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n916), .A2(new_n918), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n916), .A2(new_n918), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1104), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(G290), .A2(G1986), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT112), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n1104), .ZN(new_n1116));
  AND2_X1   g691(.A1(G290), .A2(G1986), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1100), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1113), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1099), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n861), .ZN(new_n1124));
  INV_X1    g699(.A(G1384), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n491), .B2(new_n496), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT50), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT50), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n1125), .C1(new_n491), .C2(new_n496), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1099), .B1(new_n1094), .B2(KEYINPUT45), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1126), .A2(new_n1097), .ZN(new_n1135));
  AOI21_X1  g710(.A(G1971), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n506), .B2(new_n515), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT55), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n1141));
  OAI211_X1 g716(.A(KEYINPUT55), .B(G8), .C1(new_n506), .C2(new_n515), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1137), .A2(KEYINPUT117), .A3(G8), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  OAI21_X1  g722(.A(G8), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT116), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n1155));
  INV_X1    g730(.A(G1981), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n596), .A2(new_n1156), .A3(new_n598), .A4(new_n600), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT118), .B(G86), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n534), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n600), .B(new_n1159), .C1(new_n602), .C2(new_n603), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(G1981), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1157), .A2(new_n1161), .A3(KEYINPUT49), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT49), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g738(.A(G8), .B1(new_n1126), .B2(new_n1099), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1164), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT52), .B1(G288), .B2(new_n731), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n534), .A2(KEYINPUT77), .A3(G87), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1170), .A2(G1976), .A3(new_n581), .A4(new_n582), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1171), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT52), .B1(new_n1173), .B2(new_n1164), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1155), .B1(new_n1165), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1175), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1163), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1157), .A2(new_n1161), .A3(KEYINPUT49), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n1166), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1180), .A3(KEYINPUT119), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1127), .A2(new_n1123), .A3(new_n1130), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(G2090), .ZN(new_n1184));
  OAI21_X1  g759(.A(G8), .B1(new_n1184), .B2(new_n1136), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1149), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1099), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1188), .A2(new_n806), .B1(new_n866), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(G8), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1190), .A2(new_n1191), .A3(G286), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1154), .A2(new_n1182), .A3(new_n1187), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1196), .A2(new_n1194), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1148), .A2(new_n1186), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1154), .A2(new_n1192), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT53), .ZN(new_n1201));
  INV_X1    g776(.A(G2078), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1134), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1135), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1134), .A2(KEYINPUT53), .A3(new_n1202), .A4(new_n1135), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1188), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n714), .ZN(new_n1209));
  AOI21_X1  g784(.A(G301), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  AND4_X1   g785(.A1(new_n1154), .A2(new_n1182), .A3(new_n1187), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT51), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1191), .B1(new_n1190), .B2(G168), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1214), .A2(new_n806), .A3(new_n1123), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1189), .A2(new_n866), .ZN(new_n1216));
  AOI21_X1  g791(.A(G168), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1212), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1215), .A2(G168), .A3(new_n1216), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1220), .A2(G8), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1221), .A2(KEYINPUT51), .ZN(new_n1222));
  OAI21_X1  g797(.A(KEYINPUT62), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(KEYINPUT51), .B1(new_n1221), .B2(new_n1217), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1213), .A2(new_n1212), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1211), .A2(new_n1223), .A3(new_n1227), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n1154), .A2(new_n1196), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n891), .A2(new_n731), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1157), .B1(new_n1165), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1229), .B1(new_n1166), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1200), .A2(new_n1228), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1234));
  AOI22_X1  g809(.A1(new_n1176), .A2(new_n1181), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1235));
  INV_X1    g810(.A(new_n1205), .ZN(new_n1236));
  NOR2_X1   g811(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1237));
  NOR3_X1   g812(.A1(new_n1237), .A2(new_n1203), .A3(new_n1201), .ZN(new_n1238));
  XNOR2_X1  g813(.A(G301), .B(KEYINPUT54), .ZN(new_n1239));
  NOR3_X1   g814(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1209), .A2(new_n1206), .A3(new_n1205), .ZN(new_n1241));
  AOI22_X1  g816(.A1(new_n1240), .A2(new_n1209), .B1(new_n1241), .B2(new_n1239), .ZN(new_n1242));
  NAND4_X1  g817(.A1(new_n1234), .A2(new_n1154), .A3(new_n1235), .A4(new_n1242), .ZN(new_n1243));
  XOR2_X1   g818(.A(KEYINPUT58), .B(G1341), .Z(new_n1244));
  OAI21_X1  g819(.A(new_n1244), .B1(new_n1126), .B2(new_n1099), .ZN(new_n1245));
  INV_X1    g820(.A(KEYINPUT122), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g822(.A(KEYINPUT45), .B(new_n1125), .C1(new_n491), .C2(new_n496), .ZN(new_n1248));
  NAND4_X1  g823(.A1(new_n1135), .A2(new_n1123), .A3(new_n1107), .A4(new_n1248), .ZN(new_n1249));
  OAI211_X1 g824(.A(KEYINPUT122), .B(new_n1244), .C1(new_n1126), .C2(new_n1099), .ZN(new_n1250));
  NAND3_X1  g825(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1251), .A2(new_n559), .ZN(new_n1252));
  NOR2_X1   g827(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g829(.A(new_n1251), .B(new_n559), .C1(KEYINPUT123), .C2(KEYINPUT59), .ZN(new_n1255));
  AOI22_X1  g830(.A1(new_n1254), .A2(new_n1255), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1256));
  INV_X1    g831(.A(KEYINPUT61), .ZN(new_n1257));
  XOR2_X1   g832(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n1258));
  NOR2_X1   g833(.A1(new_n573), .A2(new_n574), .ZN(new_n1259));
  INV_X1    g834(.A(KEYINPUT121), .ZN(new_n1260));
  OAI21_X1  g835(.A(new_n1260), .B1(new_n567), .B2(new_n570), .ZN(new_n1261));
  OAI211_X1 g836(.A(KEYINPUT121), .B(new_n566), .C1(new_n643), .C2(new_n498), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g838(.A(new_n1258), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g839(.A1(new_n647), .A2(KEYINPUT57), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g841(.A(KEYINPUT56), .B(G2072), .ZN(new_n1267));
  NAND3_X1  g842(.A1(new_n1134), .A2(new_n1135), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g843(.A1(new_n1183), .A2(new_n871), .ZN(new_n1269));
  AND3_X1   g844(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g845(.A(new_n1266), .B1(new_n1269), .B2(new_n1268), .ZN(new_n1271));
  OAI21_X1  g846(.A(new_n1257), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g847(.A1(new_n1272), .A2(KEYINPUT124), .ZN(new_n1273));
  INV_X1    g848(.A(KEYINPUT124), .ZN(new_n1274));
  OAI211_X1 g849(.A(new_n1274), .B(new_n1257), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1275));
  AOI21_X1  g850(.A(new_n1256), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g851(.A(new_n1271), .ZN(new_n1277));
  NAND3_X1  g852(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1278));
  NAND3_X1  g853(.A1(new_n1277), .A2(KEYINPUT61), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g854(.A1(new_n1279), .A2(KEYINPUT125), .ZN(new_n1280));
  INV_X1    g855(.A(KEYINPUT125), .ZN(new_n1281));
  NAND4_X1  g856(.A1(new_n1277), .A2(new_n1281), .A3(KEYINPUT61), .A4(new_n1278), .ZN(new_n1282));
  NAND2_X1  g857(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g858(.A1(new_n1126), .A2(new_n1099), .ZN(new_n1284));
  INV_X1    g859(.A(G2067), .ZN(new_n1285));
  NAND2_X1  g860(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g861(.A(KEYINPUT60), .B(new_n1286), .C1(new_n1188), .C2(G1348), .ZN(new_n1287));
  NOR2_X1   g862(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1288));
  NAND2_X1  g863(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1289));
  NAND2_X1  g864(.A1(new_n1289), .A2(new_n638), .ZN(new_n1290));
  INV_X1    g865(.A(new_n638), .ZN(new_n1291));
  NAND3_X1  g866(.A1(new_n1287), .A2(KEYINPUT126), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g867(.A(new_n1288), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g868(.A(G1348), .ZN(new_n1294));
  AOI22_X1  g869(.A1(new_n1208), .A2(new_n1294), .B1(new_n1285), .B2(new_n1284), .ZN(new_n1295));
  NOR2_X1   g870(.A1(new_n1295), .A2(KEYINPUT60), .ZN(new_n1296));
  OAI211_X1 g871(.A(new_n1276), .B(new_n1283), .C1(new_n1293), .C2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g872(.A(new_n1277), .B1(new_n1295), .B2(new_n1291), .ZN(new_n1298));
  NAND2_X1  g873(.A1(new_n1298), .A2(new_n1278), .ZN(new_n1299));
  AOI21_X1  g874(.A(new_n1243), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g875(.A(new_n1122), .B1(new_n1233), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g876(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1302));
  XNOR2_X1  g877(.A(new_n1302), .B(KEYINPUT46), .ZN(new_n1303));
  NOR2_X1   g878(.A1(new_n1106), .A2(new_n827), .ZN(new_n1304));
  OAI21_X1  g879(.A(new_n1303), .B1(new_n1104), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g880(.A1(new_n1305), .A2(KEYINPUT47), .ZN(new_n1306));
  NOR2_X1   g881(.A1(new_n1305), .A2(KEYINPUT47), .ZN(new_n1307));
  XNOR2_X1  g882(.A(new_n1116), .B(KEYINPUT48), .ZN(new_n1308));
  OAI22_X1  g883(.A1(new_n1306), .A2(new_n1307), .B1(new_n1113), .B2(new_n1308), .ZN(new_n1309));
  OR2_X1    g884(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1310));
  NAND2_X1  g885(.A1(new_n852), .A2(new_n1285), .ZN(new_n1311));
  AOI21_X1  g886(.A(new_n1104), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NOR2_X1   g887(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g888(.A1(new_n1301), .A2(new_n1313), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g889(.A(KEYINPUT127), .ZN(new_n1316));
  OAI21_X1  g890(.A(new_n457), .B1(new_n709), .B2(new_n710), .ZN(new_n1317));
  AOI21_X1  g891(.A(new_n1317), .B1(new_n686), .B2(new_n690), .ZN(new_n1318));
  NAND3_X1  g892(.A1(new_n778), .A2(new_n1010), .A3(new_n1318), .ZN(new_n1319));
  AOI211_X1 g893(.A(new_n1316), .B(new_n1319), .C1(new_n1072), .C2(new_n1082), .ZN(new_n1320));
  INV_X1    g894(.A(new_n1319), .ZN(new_n1321));
  AOI21_X1  g895(.A(KEYINPUT127), .B1(new_n1083), .B2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g896(.A1(new_n1320), .A2(new_n1322), .ZN(G308));
  NAND2_X1  g897(.A1(new_n1083), .A2(new_n1321), .ZN(G225));
endmodule


