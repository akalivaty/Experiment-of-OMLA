//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G107), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n188), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n187), .A2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n192), .B2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n189), .B1(new_n191), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n193), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n188), .A4(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n204), .B(G101), .C1(new_n192), .C2(new_n196), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G119), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT69), .A3(G116), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT2), .B(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n208), .A3(new_n209), .A4(new_n211), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n214), .A2(new_n220), .A3(KEYINPUT70), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT70), .B1(new_n214), .B2(new_n220), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n203), .B(new_n205), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n191), .A2(new_n188), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n194), .A2(KEYINPUT81), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n202), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n202), .A2(new_n227), .A3(KEYINPUT82), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n207), .A2(G119), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT5), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n215), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n212), .B2(new_n233), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n235), .A2(new_n220), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n223), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n223), .A2(new_n237), .A3(new_n239), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT85), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT0), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n250), .A2(KEYINPUT65), .A3(G146), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT65), .B1(new_n250), .B2(G146), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n247), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n250), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n248), .B2(G143), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n250), .A2(KEYINPUT65), .A3(G146), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n247), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n250), .A2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n249), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT0), .B(G128), .Z(new_n264));
  AOI22_X1  g078(.A1(new_n254), .A2(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT86), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G125), .ZN(new_n268));
  INV_X1    g082(.A(G125), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT86), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n272));
  OAI21_X1  g086(.A(G128), .B1(new_n255), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n259), .A2(new_n271), .B1(new_n273), .B2(new_n263), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n269), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n268), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G224), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n268), .A2(new_n270), .A3(new_n278), .A4(new_n275), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n241), .A2(new_n283), .A3(KEYINPUT6), .A4(new_n242), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n241), .A2(KEYINPUT6), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n244), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT7), .B1(new_n278), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n287), .B2(new_n278), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n268), .A2(new_n270), .A3(new_n275), .A4(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n239), .B(KEYINPUT8), .ZN(new_n291));
  INV_X1    g105(.A(new_n237), .ZN(new_n292));
  INV_X1    g106(.A(new_n228), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(new_n236), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n290), .A2(new_n295), .A3(new_n242), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n276), .B1(new_n297), .B2(new_n279), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n286), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT88), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n286), .A2(new_n299), .A3(new_n301), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G221), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n202), .A2(KEYINPUT82), .A3(new_n227), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT82), .B1(new_n202), .B2(new_n227), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n249), .B(new_n271), .C1(new_n251), .C2(new_n252), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n272), .B1(G143), .B2(new_n248), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n263), .B1(new_n316), .B2(new_n246), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n314), .A2(KEYINPUT10), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT67), .B(G131), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT11), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G137), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(G137), .ZN(new_n327));
  INV_X1    g141(.A(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT11), .A3(G134), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n326), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n331));
  INV_X1    g145(.A(G131), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  INV_X1    g149(.A(new_n315), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n246), .B1(new_n249), .B2(KEYINPUT1), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n259), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n335), .B1(new_n339), .B2(new_n228), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n254), .A2(new_n261), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n264), .A2(new_n263), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n203), .A2(new_n341), .A3(new_n342), .A4(new_n205), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n322), .A2(new_n334), .A3(new_n340), .A4(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n274), .B1(new_n312), .B2(new_n313), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n293), .B1(new_n336), .B2(new_n338), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT12), .B1(new_n347), .B2(new_n333), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT12), .ZN(new_n349));
  AOI211_X1 g163(.A(new_n349), .B(new_n334), .C1(new_n345), .C2(new_n346), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n344), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G140), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n277), .A2(G227), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n230), .A2(new_n231), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n319), .A2(KEYINPUT10), .A3(new_n321), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n343), .B(new_n340), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n358), .B2(new_n333), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n333), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n351), .A2(new_n354), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G469), .B1(new_n362), .B2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n344), .A2(new_n361), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n354), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n344), .B(new_n355), .C1(new_n348), .C2(new_n350), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT83), .B(G469), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n311), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G214), .B1(G237), .B2(G902), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT84), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n300), .A2(KEYINPUT88), .A3(new_n302), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n306), .A2(new_n370), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G217), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n308), .A2(new_n376), .A3(G953), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G128), .B(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n246), .A2(G143), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT95), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT13), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT13), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT95), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n379), .B1(new_n385), .B2(G134), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(G134), .A3(new_n379), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT94), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G122), .ZN(new_n390));
  INV_X1    g204(.A(G122), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT94), .ZN(new_n392));
  OAI21_X1  g206(.A(G116), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n391), .A2(G116), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n190), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(KEYINPUT94), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n389), .A2(G122), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n207), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G107), .B1(new_n399), .B2(new_n394), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n387), .A2(new_n388), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT14), .B1(new_n391), .B2(G116), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n207), .A3(G122), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G107), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n250), .A2(G128), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n407), .A2(new_n380), .A3(G134), .ZN(new_n408));
  AOI21_X1  g222(.A(G134), .B1(new_n407), .B2(new_n380), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n406), .A2(new_n396), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n378), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n190), .B1(new_n393), .B2(new_n395), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n399), .A2(G107), .A3(new_n394), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n385), .A2(G134), .A3(new_n379), .ZN(new_n415));
  OAI22_X1  g229(.A1(new_n413), .A2(new_n414), .B1(new_n415), .B2(new_n386), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n406), .A2(new_n396), .A3(new_n410), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n377), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT96), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n310), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n420), .B1(new_n419), .B2(new_n310), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n310), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT96), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n421), .A3(new_n423), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT97), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT97), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G113), .B(G122), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(new_n187), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G125), .B(G140), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT16), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT16), .ZN(new_n440));
  INV_X1    g254(.A(G140), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT77), .A4(G125), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(G125), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(KEYINPUT16), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n439), .A2(G146), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n269), .A2(G140), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT19), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT19), .B1(new_n444), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n248), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G237), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n277), .A3(G214), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n250), .ZN(new_n454));
  NOR2_X1   g268(.A1(G237), .A2(G953), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(G143), .A3(G214), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n323), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n454), .A2(new_n460), .A3(new_n323), .A4(new_n456), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT91), .B1(new_n457), .B2(new_n458), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n451), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n444), .A2(new_n447), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n438), .A2(new_n248), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT18), .A2(G131), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n457), .B2(new_n470), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n457), .A2(new_n472), .A3(new_n470), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n437), .B1(new_n464), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n454), .A2(new_n456), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  INV_X1    g293(.A(new_n475), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n479), .B(new_n468), .C1(new_n480), .C2(new_n473), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n463), .A2(new_n482), .A3(new_n459), .A4(new_n461), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n445), .B(new_n442), .C1(new_n465), .C2(new_n440), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n248), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n457), .A2(KEYINPUT17), .A3(new_n458), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n446), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n436), .B(new_n481), .C1(new_n484), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n477), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(G475), .A2(G902), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT92), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n497), .A3(new_n492), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n489), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n483), .A2(new_n446), .A3(new_n486), .A4(new_n487), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n436), .B1(new_n501), .B2(new_n481), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n310), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT93), .B(G475), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n277), .A2(G952), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(G234), .B2(G237), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n310), .B(new_n277), .C1(G234), .C2(G237), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT21), .B(G898), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n434), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n375), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n221), .A2(new_n222), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n328), .A2(G134), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n332), .B1(new_n518), .B2(new_n327), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n331), .B2(new_n323), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n319), .A2(new_n321), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n260), .B1(new_n259), .B2(new_n247), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n333), .B(new_n342), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(KEYINPUT30), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n327), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G131), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n330), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT68), .B1(new_n274), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT68), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n520), .A2(new_n318), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n529), .A2(new_n531), .B1(new_n265), .B2(new_n333), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n517), .B(new_n525), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n521), .A2(new_n516), .A3(new_n524), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n455), .A2(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT27), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT31), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n534), .A2(new_n542), .A3(new_n535), .A4(new_n539), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n535), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n274), .A2(new_n528), .A3(KEYINPUT68), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n530), .B1(new_n520), .B2(new_n318), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n524), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n517), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n521), .A2(new_n516), .A3(KEYINPUT28), .A4(new_n524), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n552));
  INV_X1    g366(.A(new_n539), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n541), .B(new_n543), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(G472), .A2(G902), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT73), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n561), .A3(new_n557), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n556), .A2(new_n557), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n521), .A2(new_n524), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n517), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(new_n535), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n535), .A2(new_n567), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT28), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n571), .A2(KEYINPUT29), .A3(new_n539), .A4(new_n545), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n551), .A2(new_n539), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n534), .A2(new_n535), .A3(new_n553), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n310), .B(new_n572), .C1(new_n575), .C2(KEYINPUT29), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n564), .A2(KEYINPUT32), .B1(G472), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n563), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n376), .B1(G234), .B2(new_n310), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n486), .A2(new_n446), .ZN(new_n581));
  INV_X1    g395(.A(G110), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT24), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT24), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G110), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT75), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n583), .B2(new_n585), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(G119), .B(G128), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT23), .B1(new_n246), .B2(G119), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT76), .B1(new_n246), .B2(G119), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n210), .A2(G128), .ZN(new_n594));
  OR2_X1    g408(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n589), .A2(new_n590), .B1(new_n597), .B2(G110), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n581), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n587), .A2(new_n588), .ZN(new_n600));
  INV_X1    g414(.A(new_n590), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n593), .A2(new_n596), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n600), .A2(new_n601), .B1(new_n602), .B2(new_n582), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n446), .A2(new_n467), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n603), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT78), .ZN(new_n606));
  INV_X1    g420(.A(new_n604), .ZN(new_n607));
  OAI22_X1  g421(.A1(new_n589), .A2(new_n590), .B1(G110), .B2(new_n597), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n599), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT22), .B(G137), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n613), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n599), .B(new_n615), .C1(new_n605), .C2(new_n609), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n310), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT25), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n614), .A2(KEYINPUT25), .A3(new_n310), .A4(new_n616), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n580), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n614), .A2(new_n616), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n622), .A2(G902), .A3(new_n579), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n578), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT79), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n624), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n563), .B2(new_n577), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT79), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n515), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n200), .ZN(G3));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n416), .A2(new_n417), .A3(new_n377), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n377), .B1(new_n416), .B2(new_n417), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n416), .B2(new_n417), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(KEYINPUT33), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT33), .B1(new_n401), .B2(new_n411), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n637), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n419), .A2(new_n642), .A3(new_n633), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n422), .A2(G902), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n646), .A2(new_n647), .B1(new_n422), .B2(new_n427), .ZN(new_n648));
  INV_X1    g462(.A(new_n645), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n647), .B(new_n649), .C1(new_n640), .C2(new_n643), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n511), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n506), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n301), .B1(new_n286), .B2(new_n299), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n305), .B1(new_n656), .B2(KEYINPUT98), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n655), .B(new_n373), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n556), .A2(new_n310), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n559), .A2(new_n662), .A3(new_n562), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n370), .A2(new_n624), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND3_X1  g482(.A1(new_n490), .A2(new_n494), .A3(new_n492), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n496), .A2(new_n669), .B1(new_n503), .B2(new_n504), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n434), .A2(new_n511), .A3(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n672), .B(new_n373), .C1(new_n658), .C2(new_n657), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n665), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G107), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NAND2_X1  g492(.A1(new_n619), .A2(new_n620), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n579), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n613), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n610), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n579), .A2(G902), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n434), .A3(new_n512), .ZN(new_n686));
  OR3_X1    g500(.A1(new_n375), .A2(new_n663), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  AND2_X1   g503(.A1(new_n370), .A2(new_n685), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n556), .A2(new_n561), .A3(new_n557), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n561), .B1(new_n556), .B2(new_n557), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT32), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n576), .A2(G472), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n556), .A2(KEYINPUT32), .A3(new_n557), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n690), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n286), .A2(new_n299), .A3(new_n301), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n698), .B1(new_n303), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n508), .B1(new_n509), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n433), .A2(new_n432), .A3(new_n670), .A4(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n702), .A2(new_n703), .A3(new_n373), .A4(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n373), .B(new_n707), .C1(new_n658), .C2(new_n657), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT102), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n697), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n246), .ZN(G30));
  INV_X1    g526(.A(new_n534), .ZN(new_n713));
  INV_X1    g527(.A(new_n535), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n539), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n516), .B1(new_n524), .B2(new_n521), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n714), .B2(KEYINPUT74), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n553), .A3(new_n569), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n310), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G472), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n695), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n693), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n496), .A2(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n434), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n679), .A2(new_n579), .B1(new_n683), .B2(new_n682), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n373), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n705), .B(KEYINPUT39), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n370), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n727), .B1(KEYINPUT40), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n306), .A2(new_n374), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT38), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n306), .A2(KEYINPUT38), .A3(new_n374), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n363), .A2(new_n369), .ZN(new_n736));
  INV_X1    g550(.A(new_n311), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n728), .ZN(new_n739));
  OR3_X1    g553(.A1(new_n738), .A2(KEYINPUT40), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n723), .A2(new_n730), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G143), .ZN(G45));
  AOI21_X1  g556(.A(new_n372), .B1(new_n700), .B2(new_n701), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n427), .A2(new_n422), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n649), .B1(new_n640), .B2(new_n643), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(KEYINPUT100), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n506), .B(new_n706), .C1(new_n650), .C2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n578), .A2(new_n743), .A3(new_n690), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G146), .ZN(G48));
  INV_X1    g564(.A(G469), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n367), .A2(KEYINPUT103), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n347), .A2(KEYINPUT12), .A3(new_n333), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n318), .B1(new_n230), .B2(new_n231), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n339), .A2(new_n228), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n333), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n349), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n359), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n355), .B1(new_n344), .B2(new_n361), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n310), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n753), .B1(new_n761), .B2(G469), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n737), .B(new_n369), .C1(new_n752), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT104), .ZN(new_n764));
  INV_X1    g578(.A(new_n368), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT103), .B1(new_n367), .B2(new_n751), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n753), .A3(G469), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n737), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n629), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n659), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT41), .B(G113), .Z(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G15));
  NOR2_X1   g590(.A1(new_n773), .A2(new_n673), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n207), .ZN(G18));
  AOI21_X1  g592(.A(new_n686), .B1(new_n563), .B2(new_n577), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n743), .A3(new_n764), .A4(new_n771), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  INV_X1    g595(.A(new_n557), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n541), .A2(new_n543), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n571), .A2(new_n545), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n553), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n782), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n662), .A3(new_n624), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT105), .ZN(new_n789));
  INV_X1    g603(.A(G472), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n556), .B2(new_n310), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n786), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT105), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n624), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n373), .B(new_n725), .C1(new_n658), .C2(new_n657), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n772), .A2(new_n795), .A3(new_n653), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G122), .ZN(G24));
  NOR4_X1   g613(.A1(new_n791), .A2(new_n747), .A3(new_n726), .A4(new_n786), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n743), .A3(new_n764), .A4(new_n771), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G125), .ZN(G27));
  NOR2_X1   g616(.A1(new_n564), .A2(KEYINPUT32), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n624), .B(new_n748), .C1(new_n696), .C2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n305), .A2(new_n304), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n656), .ZN(new_n807));
  INV_X1    g621(.A(new_n374), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n373), .B(new_n370), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n372), .B1(new_n306), .B2(new_n374), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT106), .B1(new_n812), .B2(new_n370), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n805), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n809), .A2(new_n810), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(KEYINPUT106), .A3(new_n370), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n625), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n818));
  AOI22_X1  g632(.A1(KEYINPUT42), .A2(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G131), .ZN(G33));
  OAI211_X1 g634(.A(new_n629), .B(new_n707), .C1(new_n811), .C2(new_n813), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT107), .B(G134), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(G36));
  INV_X1    g637(.A(KEYINPUT44), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n691), .A2(new_n692), .A3(new_n791), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n724), .B1(new_n746), .B2(new_n650), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT43), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT43), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n724), .B(new_n828), .C1(new_n746), .C2(new_n650), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n685), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n824), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT110), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n833), .B(new_n824), .C1(new_n825), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n373), .B1(new_n807), .B2(new_n808), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n827), .A2(new_n685), .A3(new_n829), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(KEYINPUT44), .A3(new_n663), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n812), .A2(KEYINPUT109), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT108), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n751), .A2(new_n310), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n344), .A2(new_n361), .A3(new_n355), .ZN(new_n845));
  INV_X1    g659(.A(new_n358), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n758), .A2(new_n754), .B1(new_n846), .B2(new_n334), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n847), .B2(new_n355), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT45), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n751), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(KEYINPUT45), .B(new_n845), .C1(new_n847), .C2(new_n355), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n843), .B1(new_n852), .B2(KEYINPUT46), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n766), .B1(new_n852), .B2(KEYINPUT46), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT46), .ZN(new_n855));
  OAI21_X1  g669(.A(G469), .B1(new_n362), .B2(KEYINPUT45), .ZN(new_n856));
  INV_X1    g670(.A(new_n851), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(KEYINPUT108), .B(new_n855), .C1(new_n858), .C2(new_n844), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(new_n737), .A3(new_n728), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n835), .A2(new_n842), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(G137), .ZN(G39));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n737), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT47), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n860), .A2(KEYINPUT47), .A3(new_n737), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n578), .A2(new_n836), .A3(new_n624), .A4(new_n747), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(G140), .ZN(G42));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n801), .A2(new_n749), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n711), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n370), .A2(new_n726), .A3(new_n706), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n722), .A2(new_n796), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n873), .A2(new_n711), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n800), .B1(new_n811), .B2(new_n813), .ZN(new_n882));
  INV_X1    g696(.A(new_n697), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n670), .A2(new_n430), .A3(new_n706), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT114), .Z(new_n885));
  NOR2_X1   g699(.A1(new_n836), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n821), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n731), .A2(new_n372), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n724), .A2(new_n426), .A3(new_n429), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n724), .B1(new_n648), .B2(new_n651), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(KEYINPUT113), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n890), .A2(KEYINPUT113), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n511), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n889), .A2(new_n665), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n780), .A2(new_n687), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n631), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n772), .B(new_n629), .C1(new_n660), .C2(new_n674), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(new_n798), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n888), .A2(new_n819), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n872), .B1(new_n881), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n814), .A2(KEYINPUT42), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n817), .A2(new_n818), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n815), .A2(new_n816), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n904), .A2(new_n800), .B1(new_n883), .B2(new_n886), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n902), .A2(new_n903), .A3(new_n905), .A4(new_n821), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n780), .A2(new_n687), .A3(new_n895), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n629), .A2(KEYINPUT79), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n629), .A2(KEYINPUT79), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n514), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n907), .A2(new_n910), .A3(new_n798), .A4(new_n898), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n801), .A2(new_n749), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n708), .A2(new_n710), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n883), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n915), .A3(new_n877), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n879), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n874), .A2(KEYINPUT52), .A3(new_n877), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n912), .A2(KEYINPUT53), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n901), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT54), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n901), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT51), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n772), .A2(new_n812), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT116), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n722), .A2(new_n624), .A3(new_n508), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n652), .A2(new_n506), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n827), .A2(new_n508), .A3(new_n829), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n772), .A2(new_n812), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n792), .A2(new_n685), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n372), .A2(new_n772), .A3(new_n734), .A4(new_n733), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n795), .A2(new_n934), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT50), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n933), .B(new_n938), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n769), .A2(new_n311), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n866), .A2(new_n867), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n838), .A2(new_n841), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n949), .A3(new_n940), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n926), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n945), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n937), .B1(new_n953), .B2(new_n943), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(new_n950), .A3(KEYINPUT51), .A4(new_n933), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n624), .B1(new_n696), .B2(new_n803), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n935), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT117), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT48), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(KEYINPUT48), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n772), .A2(new_n743), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n507), .B1(new_n962), .B2(new_n940), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n961), .B(new_n963), .C1(new_n957), .C2(new_n959), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n930), .A2(new_n931), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n891), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n952), .A2(new_n955), .A3(new_n966), .ZN(new_n967));
  OAI22_X1  g781(.A1(new_n925), .A2(new_n967), .B1(G952), .B2(G953), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n624), .A2(new_n373), .A3(new_n737), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT111), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n826), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT49), .ZN(new_n972));
  OAI221_X1 g786(.A(new_n971), .B1(new_n970), .B2(new_n969), .C1(new_n972), .C2(new_n769), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n769), .A2(new_n972), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT112), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n973), .A2(new_n975), .A3(new_n723), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n968), .B1(new_n735), .B2(new_n976), .ZN(G75));
  AND2_X1   g791(.A1(G210), .A2(G902), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n881), .A2(new_n900), .A3(new_n872), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT53), .B1(new_n912), .B2(new_n919), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT56), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n244), .A2(new_n284), .A3(new_n285), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(new_n282), .Z(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT55), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n981), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n277), .A2(G952), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n981), .A2(new_n982), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(KEYINPUT118), .A3(new_n985), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT118), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT56), .B1(new_n921), .B2(new_n978), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n986), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n992), .B2(new_n995), .ZN(G51));
  XOR2_X1   g810(.A(new_n858), .B(KEYINPUT119), .Z(new_n997));
  AND4_X1   g811(.A1(KEYINPUT120), .A2(new_n921), .A3(G902), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n310), .B1(new_n901), .B2(new_n920), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT120), .B1(new_n999), .B2(new_n997), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n844), .B(KEYINPUT57), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n901), .A2(new_n920), .A3(new_n923), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n923), .B1(new_n901), .B2(new_n920), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n759), .A2(new_n760), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n988), .B1(new_n1001), .B2(new_n1008), .ZN(G54));
  AND2_X1   g823(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n999), .A2(new_n490), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n490), .B1(new_n999), .B2(new_n1010), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1011), .A2(new_n1012), .A3(new_n988), .ZN(G60));
  NAND2_X1  g827(.A1(G478), .A2(G902), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT59), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n644), .B(new_n1015), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n989), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n644), .B1(new_n925), .B2(new_n1015), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(G63));
  INV_X1    g833(.A(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G217), .A2(G902), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT122), .ZN(new_n1022));
  XNOR2_X1  g836(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n901), .B2(new_n920), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n682), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n622), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n989), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1020), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g845(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1032), .A2(KEYINPUT61), .A3(new_n989), .A4(new_n1027), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1031), .A2(new_n1033), .ZN(G66));
  NAND2_X1  g848(.A1(G224), .A2(G953), .ZN(new_n1035));
  OAI22_X1  g849(.A1(new_n911), .A2(G953), .B1(new_n510), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n983), .B1(G898), .B2(new_n277), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT123), .Z(new_n1038));
  XNOR2_X1  g852(.A(new_n1036), .B(new_n1038), .ZN(G69));
  NOR2_X1   g853(.A1(new_n956), .A2(new_n796), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n861), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n819), .A2(new_n821), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n870), .A2(new_n862), .A3(new_n874), .ZN(new_n1043));
  OR3_X1    g857(.A1(new_n1042), .A2(new_n1043), .A3(G953), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n525), .B1(new_n532), .B2(new_n533), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n448), .A2(new_n449), .ZN(new_n1046));
  XNOR2_X1  g860(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1044), .B(new_n1047), .C1(new_n704), .C2(new_n277), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT62), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n874), .A2(KEYINPUT125), .A3(new_n1049), .A4(new_n741), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n729), .B1(new_n892), .B2(new_n893), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n812), .B(new_n1051), .C1(new_n908), .C2(new_n909), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n862), .A2(KEYINPUT126), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(KEYINPUT126), .B1(new_n862), .B2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n913), .A2(new_n915), .A3(new_n741), .ZN(new_n1056));
  AOI22_X1  g870(.A1(new_n1056), .A2(KEYINPUT62), .B1(new_n868), .B2(new_n869), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT125), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1058), .B1(new_n1056), .B2(KEYINPUT62), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g874(.A(new_n277), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g875(.A(KEYINPUT127), .ZN(new_n1062));
  XNOR2_X1  g876(.A(new_n1047), .B(KEYINPUT124), .ZN(new_n1063));
  AND3_X1   g877(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g878(.A(new_n1062), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1048), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n277), .B1(G227), .B2(G900), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g882(.A(new_n1067), .ZN(new_n1069));
  OAI211_X1 g883(.A(new_n1069), .B(new_n1048), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1068), .A2(new_n1070), .ZN(G72));
  OR3_X1    g885(.A1(new_n1055), .A2(new_n1060), .A3(new_n911), .ZN(new_n1072));
  NAND2_X1  g886(.A1(G472), .A2(G902), .ZN(new_n1073));
  XOR2_X1   g887(.A(new_n1073), .B(KEYINPUT63), .Z(new_n1074));
  AOI21_X1  g888(.A(new_n715), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g889(.A(new_n1074), .ZN(new_n1076));
  NOR2_X1   g890(.A1(new_n574), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g891(.A1(new_n921), .A2(new_n715), .A3(new_n1077), .ZN(new_n1078));
  NOR3_X1   g892(.A1(new_n1042), .A2(new_n1043), .A3(new_n911), .ZN(new_n1079));
  OAI21_X1  g893(.A(new_n574), .B1(new_n1079), .B2(new_n1076), .ZN(new_n1080));
  NAND2_X1  g894(.A1(new_n1080), .A2(new_n989), .ZN(new_n1081));
  NOR3_X1   g895(.A1(new_n1075), .A2(new_n1078), .A3(new_n1081), .ZN(G57));
endmodule


