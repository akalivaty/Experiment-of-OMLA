

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U554 ( .A(n710), .Z(n711) );
  AND2_X2 U555 ( .A1(n523), .A2(G2104), .ZN(n884) );
  NOR2_X1 U556 ( .A1(n649), .A2(n648), .ZN(n650) );
  AND2_X1 U557 ( .A1(n741), .A2(n754), .ZN(n742) );
  NOR2_X1 U558 ( .A1(G651), .A2(n586), .ZN(n788) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X1 U560 ( .A(n519), .B(KEYINPUT66), .Z(n520) );
  XNOR2_X1 U561 ( .A(n520), .B(KEYINPUT17), .ZN(n710) );
  AND2_X1 U562 ( .A1(G137), .A2(n710), .ZN(n530) );
  INV_X1 U563 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U564 ( .A1(G101), .A2(n884), .ZN(n521) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n521), .Z(n528) );
  NAND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X2 U567 ( .A(n522), .B(KEYINPUT65), .ZN(n880) );
  NAND2_X1 U568 ( .A1(G113), .A2(n880), .ZN(n526) );
  NOR2_X1 U569 ( .A1(n523), .A2(G2104), .ZN(n524) );
  XNOR2_X1 U570 ( .A(n524), .B(KEYINPUT64), .ZN(n550) );
  NAND2_X1 U571 ( .A1(G125), .A2(n550), .ZN(n525) );
  AND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U574 ( .A1(n530), .A2(n529), .ZN(G160) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n792) );
  NAND2_X1 U576 ( .A1(n792), .A2(G89), .ZN(n531) );
  XNOR2_X1 U577 ( .A(KEYINPUT4), .B(n531), .ZN(n535) );
  XNOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .ZN(n532) );
  XNOR2_X1 U579 ( .A(n532), .B(KEYINPUT67), .ZN(n586) );
  INV_X1 U580 ( .A(G651), .ZN(n537) );
  NOR2_X1 U581 ( .A1(n586), .A2(n537), .ZN(n793) );
  NAND2_X1 U582 ( .A1(n793), .A2(G76), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT77), .B(n533), .Z(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U585 ( .A(n536), .B(KEYINPUT5), .ZN(n545) );
  NAND2_X1 U586 ( .A1(G51), .A2(n788), .ZN(n542) );
  NOR2_X1 U587 ( .A1(G543), .A2(n537), .ZN(n539) );
  XNOR2_X1 U588 ( .A(KEYINPUT70), .B(KEYINPUT1), .ZN(n538) );
  XNOR2_X1 U589 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X2 U590 ( .A(KEYINPUT69), .B(n540), .ZN(n789) );
  NAND2_X1 U591 ( .A1(G63), .A2(n789), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U593 ( .A(KEYINPUT6), .B(n543), .Z(n544) );
  NAND2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U595 ( .A(n546), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U596 ( .A(G168), .B(KEYINPUT8), .Z(n547) );
  XNOR2_X1 U597 ( .A(KEYINPUT78), .B(n547), .ZN(G286) );
  NAND2_X1 U598 ( .A1(n880), .A2(G114), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G138), .A2(n710), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n555) );
  BUF_X1 U601 ( .A(n550), .Z(n881) );
  NAND2_X1 U602 ( .A1(n881), .A2(G126), .ZN(n553) );
  NAND2_X1 U603 ( .A1(n884), .A2(G102), .ZN(n551) );
  XNOR2_X1 U604 ( .A(KEYINPUT86), .B(n551), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U607 ( .A(KEYINPUT87), .ZN(n556) );
  XNOR2_X1 U608 ( .A(n557), .B(n556), .ZN(G164) );
  NAND2_X1 U609 ( .A1(G53), .A2(n788), .ZN(n559) );
  NAND2_X1 U610 ( .A1(G65), .A2(n789), .ZN(n558) );
  NAND2_X1 U611 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U612 ( .A(KEYINPUT71), .B(n560), .ZN(n564) );
  NAND2_X1 U613 ( .A1(G91), .A2(n792), .ZN(n562) );
  NAND2_X1 U614 ( .A1(G78), .A2(n793), .ZN(n561) );
  AND2_X1 U615 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U616 ( .A1(n564), .A2(n563), .ZN(G299) );
  NAND2_X1 U617 ( .A1(G52), .A2(n788), .ZN(n566) );
  NAND2_X1 U618 ( .A1(G64), .A2(n789), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U620 ( .A1(G90), .A2(n792), .ZN(n568) );
  NAND2_X1 U621 ( .A1(G77), .A2(n793), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U624 ( .A1(n571), .A2(n570), .ZN(G171) );
  INV_X1 U625 ( .A(G171), .ZN(G301) );
  NAND2_X1 U626 ( .A1(G50), .A2(n788), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G62), .A2(n789), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U629 ( .A1(G88), .A2(n792), .ZN(n575) );
  NAND2_X1 U630 ( .A1(G75), .A2(n793), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U632 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U633 ( .A(n578), .B(KEYINPUT82), .ZN(G166) );
  XOR2_X1 U634 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  NAND2_X1 U635 ( .A1(G86), .A2(n792), .ZN(n580) );
  NAND2_X1 U636 ( .A1(G48), .A2(n788), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U638 ( .A1(n793), .A2(G73), .ZN(n581) );
  XOR2_X1 U639 ( .A(KEYINPUT2), .B(n581), .Z(n582) );
  NOR2_X1 U640 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U641 ( .A1(G61), .A2(n789), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n585), .A2(n584), .ZN(G305) );
  NAND2_X1 U643 ( .A1(G87), .A2(n586), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U646 ( .A1(n789), .A2(n589), .ZN(n591) );
  NAND2_X1 U647 ( .A1(n788), .A2(G49), .ZN(n590) );
  NAND2_X1 U648 ( .A1(n591), .A2(n590), .ZN(G288) );
  NAND2_X1 U649 ( .A1(G85), .A2(n792), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G72), .A2(n793), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U652 ( .A(KEYINPUT68), .B(n594), .Z(n598) );
  NAND2_X1 U653 ( .A1(n789), .A2(G60), .ZN(n596) );
  NAND2_X1 U654 ( .A1(G47), .A2(n788), .ZN(n595) );
  AND2_X1 U655 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U656 ( .A1(n598), .A2(n597), .ZN(G290) );
  NAND2_X1 U657 ( .A1(G79), .A2(n793), .ZN(n600) );
  NAND2_X1 U658 ( .A1(G54), .A2(n788), .ZN(n599) );
  NAND2_X1 U659 ( .A1(n600), .A2(n599), .ZN(n606) );
  NAND2_X1 U660 ( .A1(n792), .A2(G92), .ZN(n601) );
  XNOR2_X1 U661 ( .A(n601), .B(KEYINPUT74), .ZN(n603) );
  NAND2_X1 U662 ( .A1(G66), .A2(n789), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U664 ( .A(KEYINPUT75), .B(n604), .Z(n605) );
  NOR2_X1 U665 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n607), .Z(n992) );
  NOR2_X1 U667 ( .A1(G164), .A2(G1384), .ZN(n728) );
  NAND2_X1 U668 ( .A1(G40), .A2(G160), .ZN(n608) );
  XOR2_X1 U669 ( .A(n608), .B(KEYINPUT90), .Z(n727) );
  NAND2_X1 U670 ( .A1(n728), .A2(n727), .ZN(n624) );
  BUF_X2 U671 ( .A(n624), .Z(n662) );
  NAND2_X1 U672 ( .A1(n662), .A2(G1341), .ZN(n609) );
  XNOR2_X1 U673 ( .A(n609), .B(KEYINPUT96), .ZN(n619) );
  NAND2_X1 U674 ( .A1(n792), .A2(G81), .ZN(n610) );
  XNOR2_X1 U675 ( .A(n610), .B(KEYINPUT12), .ZN(n612) );
  NAND2_X1 U676 ( .A1(G68), .A2(n793), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U678 ( .A(n613), .B(KEYINPUT13), .ZN(n615) );
  NAND2_X1 U679 ( .A1(G43), .A2(n788), .ZN(n614) );
  NAND2_X1 U680 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U681 ( .A1(n789), .A2(G56), .ZN(n616) );
  XOR2_X1 U682 ( .A(KEYINPUT14), .B(n616), .Z(n617) );
  NOR2_X2 U683 ( .A1(n618), .A2(n617), .ZN(n1012) );
  NAND2_X1 U684 ( .A1(n619), .A2(n1012), .ZN(n623) );
  INV_X1 U685 ( .A(KEYINPUT26), .ZN(n621) );
  INV_X1 U686 ( .A(n624), .ZN(n644) );
  NAND2_X1 U687 ( .A1(n644), .A2(G1996), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X2 U689 ( .A1(n623), .A2(n622), .ZN(n631) );
  NAND2_X1 U690 ( .A1(n992), .A2(n631), .ZN(n630) );
  AND2_X1 U691 ( .A1(G1348), .A2(n624), .ZN(n625) );
  XNOR2_X1 U692 ( .A(KEYINPUT97), .B(n625), .ZN(n627) );
  NAND2_X1 U693 ( .A1(n644), .A2(G2067), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U695 ( .A(KEYINPUT98), .B(n628), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n633) );
  OR2_X1 U697 ( .A1(n631), .A2(n992), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n638) );
  NAND2_X1 U699 ( .A1(n644), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U700 ( .A(n634), .B(KEYINPUT27), .ZN(n636) );
  INV_X1 U701 ( .A(G1956), .ZN(n967) );
  NOR2_X1 U702 ( .A1(n967), .A2(n644), .ZN(n635) );
  NOR2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n639) );
  INV_X1 U704 ( .A(G299), .ZN(n803) );
  NAND2_X1 U705 ( .A1(n639), .A2(n803), .ZN(n637) );
  NAND2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U707 ( .A1(n639), .A2(n803), .ZN(n640) );
  XOR2_X1 U708 ( .A(n640), .B(KEYINPUT28), .Z(n641) );
  NAND2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U710 ( .A(n643), .B(KEYINPUT29), .ZN(n649) );
  XNOR2_X1 U711 ( .A(G1961), .B(KEYINPUT94), .ZN(n977) );
  NAND2_X1 U712 ( .A1(n662), .A2(n977), .ZN(n646) );
  XOR2_X1 U713 ( .A(G2078), .B(KEYINPUT25), .Z(n947) );
  NAND2_X1 U714 ( .A1(n644), .A2(n947), .ZN(n645) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U716 ( .A(n647), .B(KEYINPUT95), .Z(n654) );
  NOR2_X1 U717 ( .A1(G301), .A2(n654), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT99), .ZN(n659) );
  NAND2_X1 U719 ( .A1(G8), .A2(n662), .ZN(n703) );
  NOR2_X1 U720 ( .A1(G1966), .A2(n703), .ZN(n674) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n662), .ZN(n671) );
  NOR2_X1 U722 ( .A1(n674), .A2(n671), .ZN(n651) );
  NAND2_X1 U723 ( .A1(G8), .A2(n651), .ZN(n652) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n652), .ZN(n653) );
  NOR2_X1 U725 ( .A1(G168), .A2(n653), .ZN(n656) );
  AND2_X1 U726 ( .A1(G301), .A2(n654), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U728 ( .A(KEYINPUT31), .B(n657), .Z(n658) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n672) );
  NAND2_X1 U730 ( .A1(n672), .A2(G286), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n660), .B(KEYINPUT100), .ZN(n667) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n703), .ZN(n661) );
  XOR2_X1 U733 ( .A(KEYINPUT101), .B(n661), .Z(n664) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n662), .ZN(n663) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n665), .A2(G303), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n668), .A2(G8), .ZN(n669) );
  XNOR2_X1 U739 ( .A(KEYINPUT32), .B(n669), .ZN(n693) );
  XNOR2_X1 U740 ( .A(KEYINPUT103), .B(G1981), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n670), .B(G305), .ZN(n1006) );
  AND2_X1 U742 ( .A1(n693), .A2(n1006), .ZN(n681) );
  NAND2_X1 U743 ( .A1(G8), .A2(n671), .ZN(n676) );
  INV_X1 U744 ( .A(n672), .ZN(n673) );
  NOR2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n694) );
  NAND2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n996) );
  AND2_X1 U748 ( .A1(n694), .A2(n996), .ZN(n679) );
  NOR2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NAND2_X1 U750 ( .A1(n994), .A2(KEYINPUT33), .ZN(n677) );
  NOR2_X1 U751 ( .A1(n703), .A2(n677), .ZN(n688) );
  INV_X1 U752 ( .A(n688), .ZN(n678) );
  AND2_X1 U753 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U754 ( .A1(n681), .A2(n680), .ZN(n692) );
  INV_X1 U755 ( .A(n1006), .ZN(n690) );
  INV_X1 U756 ( .A(n996), .ZN(n684) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n1014) );
  XNOR2_X1 U758 ( .A(KEYINPUT102), .B(n1014), .ZN(n682) );
  NOR2_X1 U759 ( .A1(n994), .A2(n682), .ZN(n683) );
  OR2_X1 U760 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U761 ( .A1(n703), .A2(n685), .ZN(n686) );
  NOR2_X1 U762 ( .A1(KEYINPUT33), .A2(n686), .ZN(n687) );
  OR2_X1 U763 ( .A1(n688), .A2(n687), .ZN(n689) );
  OR2_X1 U764 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U765 ( .A1(n692), .A2(n691), .ZN(n708) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n702) );
  NOR2_X1 U767 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U768 ( .A1(G8), .A2(n695), .ZN(n700) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n696) );
  XOR2_X1 U770 ( .A(n696), .B(KEYINPUT24), .Z(n697) );
  NOR2_X1 U771 ( .A1(n703), .A2(n697), .ZN(n698) );
  XOR2_X1 U772 ( .A(KEYINPUT93), .B(n698), .Z(n704) );
  INV_X1 U773 ( .A(n704), .ZN(n699) );
  AND2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n706) );
  OR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n709) );
  INV_X1 U779 ( .A(n709), .ZN(n743) );
  NAND2_X1 U780 ( .A1(G95), .A2(n884), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G131), .A2(n711), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U783 ( .A1(G107), .A2(n880), .ZN(n715) );
  NAND2_X1 U784 ( .A1(G119), .A2(n881), .ZN(n714) );
  NAND2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n890) );
  INV_X1 U787 ( .A(G1991), .ZN(n953) );
  NOR2_X1 U788 ( .A1(n890), .A2(n953), .ZN(n726) );
  NAND2_X1 U789 ( .A1(G141), .A2(n711), .ZN(n719) );
  NAND2_X1 U790 ( .A1(G129), .A2(n881), .ZN(n718) );
  NAND2_X1 U791 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U792 ( .A1(n884), .A2(G105), .ZN(n720) );
  XOR2_X1 U793 ( .A(KEYINPUT38), .B(n720), .Z(n721) );
  NOR2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n724) );
  NAND2_X1 U795 ( .A1(n880), .A2(G117), .ZN(n723) );
  NAND2_X1 U796 ( .A1(n724), .A2(n723), .ZN(n862) );
  AND2_X1 U797 ( .A1(G1996), .A2(n862), .ZN(n725) );
  NOR2_X1 U798 ( .A1(n726), .A2(n725), .ZN(n926) );
  INV_X1 U799 ( .A(n727), .ZN(n729) );
  NOR2_X1 U800 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U801 ( .A(KEYINPUT91), .B(n730), .Z(n758) );
  XOR2_X1 U802 ( .A(KEYINPUT92), .B(n758), .Z(n731) );
  NOR2_X1 U803 ( .A1(n926), .A2(n731), .ZN(n751) );
  INV_X1 U804 ( .A(n751), .ZN(n741) );
  XNOR2_X1 U805 ( .A(G2067), .B(KEYINPUT37), .ZN(n756) );
  NAND2_X1 U806 ( .A1(G104), .A2(n884), .ZN(n733) );
  NAND2_X1 U807 ( .A1(G140), .A2(n711), .ZN(n732) );
  NAND2_X1 U808 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U809 ( .A(KEYINPUT34), .B(n734), .ZN(n739) );
  NAND2_X1 U810 ( .A1(G116), .A2(n880), .ZN(n736) );
  NAND2_X1 U811 ( .A1(G128), .A2(n881), .ZN(n735) );
  NAND2_X1 U812 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U813 ( .A(KEYINPUT35), .B(n737), .Z(n738) );
  NOR2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n740), .ZN(n875) );
  NOR2_X1 U816 ( .A1(n756), .A2(n875), .ZN(n924) );
  NAND2_X1 U817 ( .A1(n758), .A2(n924), .ZN(n754) );
  NAND2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U819 ( .A(KEYINPUT104), .B(n744), .Z(n747) );
  XOR2_X1 U820 ( .A(KEYINPUT89), .B(G1986), .Z(n745) );
  XNOR2_X1 U821 ( .A(G290), .B(n745), .ZN(n999) );
  NAND2_X1 U822 ( .A1(n999), .A2(n758), .ZN(n746) );
  NAND2_X1 U823 ( .A1(n747), .A2(n746), .ZN(n761) );
  NOR2_X1 U824 ( .A1(G1996), .A2(n862), .ZN(n932) );
  AND2_X1 U825 ( .A1(n953), .A2(n890), .ZN(n920) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n748) );
  XOR2_X1 U827 ( .A(n748), .B(KEYINPUT105), .Z(n749) );
  NOR2_X1 U828 ( .A1(n920), .A2(n749), .ZN(n750) );
  NOR2_X1 U829 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U830 ( .A1(n932), .A2(n752), .ZN(n753) );
  XNOR2_X1 U831 ( .A(n753), .B(KEYINPUT39), .ZN(n755) );
  NAND2_X1 U832 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U833 ( .A1(n756), .A2(n875), .ZN(n937) );
  NAND2_X1 U834 ( .A1(n757), .A2(n937), .ZN(n759) );
  NAND2_X1 U835 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U837 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G82), .ZN(G220) );
  INV_X1 U840 ( .A(G108), .ZN(G238) );
  NAND2_X1 U841 ( .A1(G7), .A2(G661), .ZN(n763) );
  XNOR2_X1 U842 ( .A(n763), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U843 ( .A(G223), .ZN(n828) );
  NAND2_X1 U844 ( .A1(n828), .A2(G567), .ZN(n764) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(n764), .Z(G234) );
  XNOR2_X1 U846 ( .A(G860), .B(KEYINPUT73), .ZN(n771) );
  INV_X1 U847 ( .A(n771), .ZN(n765) );
  NAND2_X1 U848 ( .A1(n1012), .A2(n765), .ZN(G153) );
  INV_X1 U849 ( .A(n992), .ZN(n900) );
  NOR2_X1 U850 ( .A1(G868), .A2(n900), .ZN(n767) );
  INV_X1 U851 ( .A(G868), .ZN(n809) );
  NOR2_X1 U852 ( .A1(n809), .A2(G301), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U854 ( .A(KEYINPUT76), .B(n768), .ZN(G284) );
  NAND2_X1 U855 ( .A1(G868), .A2(G286), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G299), .A2(n809), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(G297) );
  NAND2_X1 U858 ( .A1(n771), .A2(G559), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n772), .A2(n992), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G559), .A2(n809), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n992), .A2(n774), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n1012), .A2(n809), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U865 ( .A(KEYINPUT79), .B(n777), .ZN(G282) );
  NAND2_X1 U866 ( .A1(n881), .A2(G123), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(KEYINPUT18), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n884), .A2(G99), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n880), .A2(G111), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G135), .A2(n711), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n919) );
  XNOR2_X1 U874 ( .A(n919), .B(G2096), .ZN(n786) );
  INV_X1 U875 ( .A(G2100), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(G156) );
  NAND2_X1 U877 ( .A1(G559), .A2(n992), .ZN(n787) );
  XOR2_X1 U878 ( .A(n787), .B(n1012), .Z(n807) );
  NOR2_X1 U879 ( .A1(G860), .A2(n807), .ZN(n800) );
  NAND2_X1 U880 ( .A1(G55), .A2(n788), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G67), .A2(n789), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G93), .A2(n792), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G80), .A2(n793), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U886 ( .A(KEYINPUT81), .B(n796), .Z(n797) );
  OR2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n810) );
  XOR2_X1 U888 ( .A(n810), .B(KEYINPUT80), .Z(n799) );
  XNOR2_X1 U889 ( .A(n800), .B(n799), .ZN(G145) );
  XOR2_X1 U890 ( .A(n810), .B(G305), .Z(n801) );
  XNOR2_X1 U891 ( .A(n801), .B(G166), .ZN(n802) );
  XNOR2_X1 U892 ( .A(KEYINPUT19), .B(n802), .ZN(n805) );
  XNOR2_X1 U893 ( .A(G288), .B(n803), .ZN(n804) );
  XNOR2_X1 U894 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n806), .B(G290), .ZN(n896) );
  XNOR2_X1 U896 ( .A(n896), .B(n807), .ZN(n808) );
  NOR2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n812) );
  NOR2_X1 U898 ( .A1(G868), .A2(n810), .ZN(n811) );
  NOR2_X1 U899 ( .A1(n812), .A2(n811), .ZN(G295) );
  XOR2_X1 U900 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n816) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n813) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U903 ( .A1(n814), .A2(G2090), .ZN(n815) );
  XNOR2_X1 U904 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U905 ( .A1(G2072), .A2(n817), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U907 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NAND2_X1 U908 ( .A1(G120), .A2(G69), .ZN(n818) );
  XOR2_X1 U909 ( .A(KEYINPUT85), .B(n818), .Z(n819) );
  NOR2_X1 U910 ( .A1(G238), .A2(n819), .ZN(n820) );
  NAND2_X1 U911 ( .A1(G57), .A2(n820), .ZN(n832) );
  NAND2_X1 U912 ( .A1(n832), .A2(G567), .ZN(n826) );
  NOR2_X1 U913 ( .A1(G219), .A2(G220), .ZN(n821) );
  XNOR2_X1 U914 ( .A(KEYINPUT22), .B(n821), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n822), .A2(G96), .ZN(n823) );
  NOR2_X1 U916 ( .A1(G218), .A2(n823), .ZN(n824) );
  XOR2_X1 U917 ( .A(KEYINPUT84), .B(n824), .Z(n833) );
  NAND2_X1 U918 ( .A1(n833), .A2(G2106), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n834) );
  NAND2_X1 U920 ( .A1(G483), .A2(G661), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n834), .A2(n827), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U925 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U927 ( .A1(n831), .A2(n830), .ZN(G188) );
  XNOR2_X1 U928 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n833), .A2(n832), .ZN(G325) );
  XOR2_X1 U930 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(n834), .ZN(G319) );
  XNOR2_X1 U935 ( .A(G1976), .B(KEYINPUT41), .ZN(n844) );
  XOR2_X1 U936 ( .A(G1971), .B(G1956), .Z(n836) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1961), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U939 ( .A(G1991), .B(G1996), .Z(n838) );
  XNOR2_X1 U940 ( .A(G1981), .B(G1966), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U942 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U943 ( .A(G2474), .B(KEYINPUT110), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(G229) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2084), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2072), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n847), .B(G2100), .Z(n849) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U953 ( .A(G2678), .B(KEYINPUT109), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n853), .B(n852), .Z(G227) );
  NAND2_X1 U956 ( .A1(n881), .A2(G124), .ZN(n854) );
  XOR2_X1 U957 ( .A(KEYINPUT111), .B(n854), .Z(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G100), .A2(n884), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U961 ( .A1(n880), .A2(G112), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G136), .A2(n711), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U964 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U965 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n864) );
  XOR2_X1 U966 ( .A(n862), .B(KEYINPUT48), .Z(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U968 ( .A(G164), .B(n865), .ZN(n879) );
  NAND2_X1 U969 ( .A1(n880), .A2(G115), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n866), .B(KEYINPUT114), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G127), .A2(n881), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n869), .B(KEYINPUT47), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G103), .A2(n884), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G139), .A2(n711), .ZN(n872) );
  XNOR2_X1 U977 ( .A(KEYINPUT113), .B(n872), .ZN(n873) );
  NOR2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n927) );
  XNOR2_X1 U979 ( .A(n927), .B(n919), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n875), .B(G162), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n894) );
  NAND2_X1 U983 ( .A1(G118), .A2(n880), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G130), .A2(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G106), .A2(n884), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G142), .A2(n711), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n891) );
  XOR2_X1 U991 ( .A(n891), .B(n890), .Z(n892) );
  XNOR2_X1 U992 ( .A(G160), .B(n892), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U994 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U995 ( .A(G286), .B(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(G171), .B(n1012), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(n900), .B(n899), .Z(n901) );
  NOR2_X1 U999 ( .A1(G37), .A2(n901), .ZN(n902) );
  XOR2_X1 U1000 ( .A(KEYINPUT115), .B(n902), .Z(G397) );
  XOR2_X1 U1001 ( .A(KEYINPUT106), .B(G2446), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G2438), .B(G2427), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(n905), .B(G2451), .Z(n907) );
  XNOR2_X1 U1005 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1007 ( .A(G2430), .B(G2443), .Z(n909) );
  XNOR2_X1 U1008 ( .A(G2435), .B(G2454), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1010 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1011 ( .A1(G14), .A2(n912), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G57), .ZN(G237) );
  INV_X1 U1020 ( .A(n918), .ZN(G401) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n940) );
  XOR2_X1 U1026 ( .A(G2072), .B(n927), .Z(n929) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1029 ( .A(KEYINPUT50), .B(n930), .Z(n936) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT116), .B(n934), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n944), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1041 ( .A(G2090), .B(G35), .Z(n961) );
  XNOR2_X1 U1042 ( .A(KEYINPUT117), .B(G2067), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(G26), .ZN(n952) );
  XOR2_X1 U1044 ( .A(G32), .B(G1996), .Z(n946) );
  NAND2_X1 U1045 ( .A1(n946), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G27), .B(n947), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n948), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n957) );
  XOR2_X1 U1050 ( .A(G2072), .B(G33), .Z(n955) );
  XNOR2_X1 U1051 ( .A(n953), .B(G25), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(n958), .B(KEYINPUT53), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(n959), .B(KEYINPUT119), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G34), .B(G2084), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n962), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1060 ( .A(KEYINPUT55), .B(n965), .Z(n966) );
  NOR2_X1 U1061 ( .A1(G29), .A2(n966), .ZN(n1026) );
  XNOR2_X1 U1062 ( .A(G20), .B(n967), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G6), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1067 ( .A(KEYINPUT59), .B(G1348), .Z(n972) );
  XNOR2_X1 U1068 ( .A(G4), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1070 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n975) );
  XNOR2_X1 U1071 ( .A(n976), .B(n975), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(n977), .B(G5), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G21), .B(G1966), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G1976), .B(G23), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1079 ( .A(G1986), .B(KEYINPUT126), .Z(n984) );
  XNOR2_X1 U1080 ( .A(G24), .B(n984), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n987), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1084 ( .A(KEYINPUT61), .B(n990), .Z(n991) );
  NOR2_X1 U1085 ( .A1(G16), .A2(n991), .ZN(n1023) );
  XOR2_X1 U1086 ( .A(KEYINPUT56), .B(G16), .Z(n1020) );
  XNOR2_X1 U1087 ( .A(n992), .B(G1348), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(n993), .B(KEYINPUT121), .ZN(n1018) );
  XOR2_X1 U1089 ( .A(n994), .B(KEYINPUT122), .Z(n995) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1091 ( .A(KEYINPUT123), .B(n997), .Z(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G171), .B(G1961), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(G1971), .A2(G303), .ZN(n1000) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1096 ( .A(G1956), .B(G299), .ZN(n1002) );
  NOR2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G168), .ZN(n1007) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1008), .B(KEYINPUT57), .ZN(n1009) );
  XOR2_X1 U1102 ( .A(KEYINPUT120), .B(n1009), .Z(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(G1341), .B(n1012), .Z(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(KEYINPUT124), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(G11), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1027), .Z(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

