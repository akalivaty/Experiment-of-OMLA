//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT75), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT2), .B1(new_n204), .B2(new_n206), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n212), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT75), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OR3_X1    g018(.A1(new_n205), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n204), .A2(KEYINPUT76), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT77), .B(G148gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n203), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n212), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G211gat), .A2(G218gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT71), .ZN(new_n230));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT71), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n227), .A2(new_n232), .A3(new_n228), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G211gat), .ZN(new_n235));
  INV_X1    g034(.A(G218gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(new_n227), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n239), .A2(new_n230), .A3(new_n231), .A4(new_n233), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT29), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n226), .B(KEYINPUT81), .C1(new_n243), .C2(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(G228gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n242), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n215), .A2(new_n218), .B1(new_n223), .B2(new_n224), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT29), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n244), .B(new_n246), .C1(new_n247), .C2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n226), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT81), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT82), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n248), .A2(new_n249), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n247), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n245), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n254), .A4(new_n244), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n245), .B(KEYINPUT80), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n237), .A2(new_n227), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT29), .B1(new_n234), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n268), .B2(new_n234), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n249), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n226), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n266), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n264), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G78gat), .B(G106gat), .ZN(new_n276));
  INV_X1    g075(.A(G50gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n278), .B(new_n279), .Z(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT83), .B(G22gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n280), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n274), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n282), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n283), .B1(new_n264), .B2(new_n274), .ZN(new_n287));
  AOI211_X1 g086(.A(new_n280), .B(new_n273), .C1(new_n256), .C2(new_n263), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G127gat), .B(G134gat), .ZN(new_n291));
  INV_X1    g090(.A(G113gat), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT68), .B(G120gat), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G113gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n295), .A2(new_n297), .A3(KEYINPUT70), .A4(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n291), .A3(new_n294), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT68), .B(G120gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(new_n292), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT1), .B1(new_n292), .B2(new_n293), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n292), .B2(new_n293), .ZN(new_n307));
  INV_X1    g106(.A(new_n291), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n312), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G183gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT27), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT27), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G183gat), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT66), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT66), .B1(new_n321), .B2(new_n323), .ZN(new_n325));
  INV_X1    g124(.A(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n321), .A2(new_n323), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT28), .B1(new_n329), .B2(new_n326), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n311), .B(new_n319), .C1(new_n328), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n333), .A2(new_n312), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n326), .ZN(new_n336));
  NAND3_X1  g135(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(KEYINPUT65), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n338), .A2(KEYINPUT65), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n334), .B(new_n335), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n320), .A2(new_n326), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n336), .B(new_n337), .C1(new_n342), .C2(KEYINPUT24), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  AND4_X1   g143(.A1(new_n344), .A2(new_n335), .A3(new_n312), .A4(new_n333), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n341), .A2(KEYINPUT25), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n310), .A2(new_n331), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n346), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n299), .A2(new_n304), .B1(new_n308), .B2(new_n307), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G227gat), .ZN(new_n351));
  INV_X1    g150(.A(G233gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n353), .B(KEYINPUT64), .Z(new_n354));
  NAND3_X1  g153(.A1(new_n347), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G15gat), .B(G43gat), .Z(new_n359));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n350), .ZN(new_n363));
  INV_X1    g162(.A(new_n353), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n354), .A2(KEYINPUT34), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n365), .A2(KEYINPUT34), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n361), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n355), .B(KEYINPUT32), .C1(new_n357), .C2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n369), .B2(new_n362), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n290), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n305), .A2(new_n248), .A3(new_n309), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n349), .A2(new_n248), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(KEYINPUT4), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n349), .A2(new_n383), .A3(new_n248), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n226), .A2(new_n386), .A3(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT78), .B1(new_n248), .B2(new_n249), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n257), .A4(new_n310), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n375), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n385), .A2(new_n389), .A3(KEYINPUT5), .A4(new_n375), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399));
  INV_X1    g198(.A(new_n397), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n391), .A2(new_n400), .A3(new_n392), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n391), .A2(KEYINPUT6), .A3(new_n400), .A4(new_n392), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n331), .B2(new_n346), .ZN(new_n405));
  AND2_X1   g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n348), .A2(new_n406), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n260), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT73), .ZN(new_n411));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n348), .A2(new_n406), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n247), .C1(new_n406), .C2(new_n405), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n409), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n413), .B(KEYINPUT74), .Z(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n409), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT30), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n409), .A2(new_n415), .ZN(new_n421));
  INV_X1    g220(.A(new_n413), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n404), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n202), .B1(new_n374), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n402), .B2(new_n403), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n428), .A2(KEYINPUT35), .A3(new_n290), .A4(new_n373), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n409), .A2(new_n415), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT38), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n409), .B2(new_n415), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n416), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n422), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT38), .B1(new_n438), .B2(new_n435), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n402), .A2(new_n437), .A3(new_n403), .A4(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n375), .B1(new_n385), .B2(new_n389), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n400), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n310), .A2(new_n226), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n375), .A3(new_n377), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT39), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI221_X1 g248(.A(new_n443), .B1(KEYINPUT85), .B2(KEYINPUT40), .C1(new_n441), .C2(new_n446), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n424), .A2(new_n449), .A3(new_n401), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n440), .A2(new_n451), .A3(new_n290), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT86), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n440), .A2(new_n451), .A3(new_n290), .A4(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n371), .B2(new_n372), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n362), .A2(new_n369), .ZN(new_n459));
  INV_X1    g258(.A(new_n367), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT36), .A3(new_n370), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n428), .B2(new_n290), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n463), .B(KEYINPUT84), .C1(new_n428), .C2(new_n290), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n430), .B1(new_n456), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n471));
  INV_X1    g270(.A(G8gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473));
  INV_X1    g272(.A(G1gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT16), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n473), .A2(G1gat), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n471), .B(new_n472), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n473), .A2(G1gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g280(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n478), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n478), .B2(new_n483), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT17), .ZN(new_n488));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT15), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  INV_X1    g291(.A(G43gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(G50gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n277), .A2(G43gat), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT87), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT14), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n491), .A2(new_n496), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n491), .A2(new_n503), .A3(new_n496), .A4(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(KEYINPUT15), .A3(new_n489), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n488), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n510), .ZN(new_n512));
  AOI211_X1 g311(.A(KEYINPUT17), .B(new_n512), .C1(new_n506), .C2(new_n507), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n470), .B(new_n487), .C1(new_n511), .C2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT87), .B1(new_n494), .B2(new_n495), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n509), .B1(new_n515), .B2(KEYINPUT15), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT88), .B1(new_n516), .B2(new_n496), .ZN(new_n517));
  INV_X1    g316(.A(new_n507), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n478), .A2(new_n483), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n512), .B1(new_n506), .B2(new_n507), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n488), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n470), .B1(new_n527), .B2(new_n487), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n529), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n487), .B1(new_n511), .B2(new_n513), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT91), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(new_n530), .A3(new_n522), .A4(new_n514), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n530), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n520), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(new_n522), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n535), .B2(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G197gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT11), .B(G169gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT12), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n538), .A2(new_n552), .A3(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n469), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G57gat), .B(G64gat), .Z(new_n556));
  NAND2_X1  g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G71gat), .B(G78gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G127gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n520), .B1(new_n562), .B2(new_n563), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  INV_X1    g371(.A(G155gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n569), .A2(new_n570), .A3(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT41), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT95), .B(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT7), .ZN(new_n593));
  INV_X1    g392(.A(G99gat), .ZN(new_n594));
  INV_X1    g393(.A(G106gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT8), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G99gat), .B(G106gat), .Z(new_n598));
  OR2_X1    g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n524), .B2(new_n526), .ZN(new_n603));
  OAI22_X1  g402(.A1(new_n525), .A2(new_n601), .B1(new_n583), .B2(new_n582), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n588), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n601), .B1(new_n511), .B2(new_n513), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  INV_X1    g406(.A(new_n588), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n587), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n604), .B1(new_n527), .B2(new_n601), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n586), .B1(new_n613), .B2(new_n608), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n606), .A2(new_n607), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(KEYINPUT96), .A3(new_n588), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT96), .B1(new_n615), .B2(new_n588), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n609), .A2(new_n587), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(KEYINPUT97), .A3(new_n616), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n610), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT98), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n601), .A2(new_n562), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n560), .B(new_n561), .Z(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n599), .A3(new_n600), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n626), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n629), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n626), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  OR2_X1    g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n631), .A2(new_n632), .ZN(new_n640));
  INV_X1    g439(.A(new_n626), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n634), .A2(new_n626), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n638), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n580), .A2(new_n624), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n555), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n404), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n474), .ZN(G1324gat));
  OAI21_X1  g455(.A(KEYINPUT101), .B1(new_n649), .B2(new_n425), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n555), .A2(new_n658), .A3(new_n424), .A4(new_n648), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(G8gat), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n555), .A2(new_n648), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND4_X1  g461(.A1(new_n661), .A2(KEYINPUT42), .A3(new_n424), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n657), .B2(new_n659), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n660), .B(new_n663), .C1(new_n665), .C2(new_n666), .ZN(G1325gat));
  INV_X1    g466(.A(new_n463), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT103), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n649), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n661), .A2(new_n373), .ZN(new_n672));
  INV_X1    g471(.A(G15gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n671), .B1(new_n675), .B2(new_n677), .ZN(G1326gat));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  INV_X1    g478(.A(new_n290), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n661), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT104), .B1(new_n649), .B2(new_n290), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n681), .B2(new_n682), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(G1327gat));
  NOR2_X1   g485(.A1(new_n580), .A2(new_n645), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n624), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n555), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n497), .A3(new_n653), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n624), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n469), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n610), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT97), .B1(new_n622), .B2(new_n616), .ZN(new_n698));
  AND4_X1   g497(.A1(KEYINPUT97), .A2(new_n612), .A3(new_n614), .A4(new_n616), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n464), .B1(new_n453), .B2(new_n455), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n427), .A2(new_n429), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n694), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n538), .A2(new_n552), .A3(new_n544), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n552), .B1(new_n538), .B2(new_n544), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n688), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(new_n653), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G29gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n691), .A2(new_n692), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n693), .A2(new_n711), .A3(new_n712), .ZN(G1328gat));
  NOR2_X1   g512(.A1(new_n425), .A2(G36gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n555), .A2(new_n689), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT46), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n696), .A2(new_n704), .A3(new_n424), .A4(new_n709), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G36gat), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n555), .A2(new_n719), .A3(new_n689), .A4(new_n714), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n716), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT105), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n716), .A2(new_n718), .A3(new_n723), .A4(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1329gat));
  NAND4_X1  g524(.A1(new_n696), .A2(new_n704), .A3(new_n668), .A4(new_n709), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G43gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n690), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n373), .A2(new_n493), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT47), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OAI221_X1 g532(.A(new_n727), .B1(new_n731), .B2(KEYINPUT47), .C1(new_n728), .C2(new_n729), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1330gat));
  NAND3_X1  g534(.A1(new_n690), .A2(new_n277), .A3(new_n680), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n696), .A2(new_n704), .A3(new_n680), .A4(new_n709), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n277), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n705), .A2(KEYINPUT107), .A3(new_n680), .A4(new_n709), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(KEYINPUT48), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n739), .A2(KEYINPUT48), .B1(new_n743), .B2(new_n744), .ZN(G1331gat));
  OAI21_X1  g544(.A(new_n430), .B1(new_n456), .B2(new_n464), .ZN(new_n746));
  INV_X1    g545(.A(new_n580), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n554), .A2(new_n747), .A3(new_n700), .A4(new_n646), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n653), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n424), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT49), .B(G64gat), .Z(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n746), .A2(new_n373), .A3(new_n748), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n757));
  AOI21_X1  g556(.A(G71gat), .B1(new_n756), .B2(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n749), .A2(G71gat), .A3(new_n668), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n749), .A2(new_n680), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g563(.A(KEYINPUT109), .B1(new_n554), .B2(new_n580), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n708), .A2(new_n766), .A3(new_n747), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n646), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n705), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n654), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n767), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n700), .A4(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n700), .B(new_n771), .C1(new_n701), .C2(new_n702), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(KEYINPUT110), .A3(new_n775), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n653), .A2(new_n589), .A3(new_n645), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n770), .A2(new_n589), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  NAND3_X1  g580(.A1(new_n645), .A2(new_n590), .A3(new_n424), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT112), .Z(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n777), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n777), .A2(new_n787), .A3(new_n778), .A4(new_n784), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n696), .A2(new_n704), .A3(new_n424), .A4(new_n768), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(new_n789), .B2(G92gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n789), .A2(KEYINPUT111), .A3(G92gat), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT111), .B1(new_n789), .B2(G92gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n783), .B1(new_n772), .B2(new_n776), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n769), .B2(new_n463), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n373), .A2(new_n645), .A3(new_n594), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n779), .B2(new_n799), .ZN(G1338gat));
  NAND3_X1  g599(.A1(new_n705), .A2(new_n680), .A3(new_n768), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n290), .A2(new_n646), .A3(G106gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n779), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n772), .B2(new_n776), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n801), .B2(G106gat), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n804), .A2(new_n807), .B1(new_n809), .B2(new_n803), .ZN(G1339gat));
  NAND3_X1  g609(.A1(new_n522), .A2(new_n542), .A3(new_n541), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT114), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n522), .A2(new_n542), .A3(new_n813), .A4(new_n541), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n534), .A2(new_n522), .A3(new_n514), .ZN(new_n816));
  INV_X1    g615(.A(new_n530), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n549), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n514), .A2(new_n522), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n530), .B1(new_n822), .B2(new_n534), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n821), .B(new_n549), .C1(new_n823), .C2(new_n815), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n553), .A2(new_n825), .A3(new_n645), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n553), .A2(new_n825), .A3(KEYINPUT117), .A4(new_n645), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n631), .A2(new_n632), .A3(new_n626), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n638), .B1(new_n633), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n836), .A2(new_n644), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n706), .B2(new_n707), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n828), .A2(new_n829), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n624), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n700), .A2(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n553), .A2(new_n825), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT116), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n553), .A2(new_n825), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n644), .A3(new_n837), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n619), .A2(new_n623), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n697), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n580), .B1(new_n841), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n647), .A2(new_n554), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR4_X1   g653(.A1(new_n854), .A2(new_n424), .A3(new_n374), .A4(new_n654), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n554), .ZN(new_n856));
  AND2_X1   g655(.A1(KEYINPUT118), .A2(G113gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(KEYINPUT118), .A2(G113gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  INV_X1    g659(.A(new_n855), .ZN(new_n861));
  OAI21_X1  g660(.A(G120gat), .B1(new_n861), .B2(new_n646), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n645), .A2(new_n302), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT119), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n861), .B2(new_n864), .ZN(G1341gat));
  NAND2_X1  g664(.A1(new_n855), .A2(new_n580), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(G127gat), .ZN(G1342gat));
  OAI21_X1  g666(.A(G134gat), .B1(new_n861), .B2(new_n624), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n852), .A2(new_n853), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n654), .A2(new_n374), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n624), .A2(G134gat), .A3(new_n424), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n868), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  AOI21_X1  g674(.A(new_n846), .B1(new_n551), .B2(new_n553), .ZN(new_n876));
  INV_X1    g675(.A(new_n826), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n624), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n853), .B1(new_n879), .B2(new_n747), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n290), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n882), .B(new_n680), .C1(new_n852), .C2(new_n853), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n654), .A2(new_n424), .A3(new_n668), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n881), .A2(new_n883), .A3(new_n554), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G141gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n680), .B1(new_n852), .B2(new_n853), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n654), .A2(new_n668), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n554), .A2(new_n203), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT120), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n888), .A2(new_n425), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n886), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1344gat));
  NOR3_X1   g696(.A1(new_n887), .A2(new_n668), .A3(new_n654), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n425), .ZN(new_n899));
  INV_X1    g698(.A(new_n222), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n645), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n848), .A2(KEYINPUT122), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n842), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n905), .A3(new_n845), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n878), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n747), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n853), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n290), .A2(KEYINPUT57), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n887), .A2(KEYINPUT57), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n645), .A3(new_n884), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n902), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n646), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n222), .A2(new_n902), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n901), .B1(new_n915), .B2(new_n919), .ZN(G1345gat));
  NAND3_X1  g719(.A1(new_n899), .A2(new_n573), .A3(new_n580), .ZN(new_n921));
  OAI21_X1  g720(.A(G155gat), .B1(new_n916), .B2(new_n747), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n916), .B2(new_n624), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n624), .A2(G162gat), .A3(new_n424), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n898), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1347gat));
  NAND2_X1  g726(.A1(new_n654), .A2(new_n424), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(new_n374), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n854), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n554), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n645), .ZN(new_n933));
  XOR2_X1   g732(.A(KEYINPUT123), .B(G176gat), .Z(new_n934));
  XNOR2_X1  g733(.A(new_n933), .B(new_n934), .ZN(G1349gat));
  INV_X1    g734(.A(new_n929), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n869), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n320), .B1(new_n937), .B2(new_n747), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n930), .B(new_n580), .C1(new_n325), .C2(new_n324), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1350gat));
  OAI22_X1  g742(.A1(new_n937), .A2(new_n624), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(G1351gat));
  NOR4_X1   g745(.A1(new_n653), .A2(new_n425), .A3(new_n290), .A4(new_n668), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n869), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n869), .A2(new_n947), .A3(KEYINPUT124), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n554), .A3(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n654), .A2(new_n424), .A3(new_n463), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n913), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n708), .A2(new_n953), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n952), .A2(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  NAND2_X1  g757(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n911), .A2(new_n912), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n645), .A4(new_n955), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n913), .A2(KEYINPUT126), .A3(new_n645), .A4(new_n955), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(G204gat), .A3(new_n964), .ZN(new_n965));
  AOI211_X1 g764(.A(G204gat), .B(new_n646), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n869), .A2(new_n947), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n965), .A2(new_n969), .ZN(G1353gat));
  NAND4_X1  g769(.A1(new_n959), .A2(new_n960), .A3(new_n580), .A4(new_n955), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n950), .A2(new_n951), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n580), .A2(new_n235), .ZN(new_n975));
  OAI22_X1  g774(.A1(new_n972), .A2(new_n973), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  NAND3_X1  g775(.A1(new_n950), .A2(new_n700), .A3(new_n951), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n700), .A2(G218gat), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  AOI22_X1  g778(.A1(new_n977), .A2(new_n236), .B1(new_n956), .B2(new_n979), .ZN(G1355gat));
endmodule


