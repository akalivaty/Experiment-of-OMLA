//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G137), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n469), .B1(new_n474), .B2(KEYINPUT68), .ZN(new_n475));
  INV_X1    g050(.A(new_n473), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G137), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n478), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT69), .Z(G160));
  NOR2_X1   g057(.A1(new_n470), .A2(new_n471), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n483), .A2(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n464), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n488), .A2(G136), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n487), .A2(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n465), .B2(new_n466), .ZN(new_n495));
  NAND2_X1  g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n484), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n465), .B2(new_n466), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n484), .C1(new_n470), .C2(new_n471), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n498), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(G50), .A2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n518), .B(new_n509), .C1(new_n514), .C2(new_n515), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n517), .A2(new_n519), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n524), .A2(KEYINPUT6), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT72), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n528), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n522), .A2(new_n509), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n537), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n536), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n535), .A2(G52), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n524), .ZN(new_n546));
  INV_X1    g121(.A(new_n540), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n547), .A2(G81), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n532), .A2(G43), .A3(G543), .A4(new_n534), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n512), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND4_X1  g139(.A1(new_n532), .A2(G53), .A3(G543), .A4(new_n534), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT74), .B1(new_n540), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n522), .A2(new_n509), .A3(new_n570), .A4(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n522), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n524), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n512), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n579), .A2(KEYINPUT75), .A3(G651), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n576), .A2(new_n580), .B1(new_n566), .B2(new_n565), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n573), .A2(new_n581), .ZN(G299));
  OR2_X1    g157(.A1(new_n536), .A2(new_n542), .ZN(G286));
  NAND2_X1  g158(.A1(new_n547), .A2(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  OAI221_X1 g165(.A(new_n584), .B1(new_n585), .B2(new_n586), .C1(new_n589), .C2(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n524), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n540), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  AND2_X1   g174(.A1(G72), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n522), .B2(G60), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n524), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n602), .A2(new_n603), .B1(new_n585), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n547), .A2(G85), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n512), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n608), .B2(new_n600), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n606), .B1(new_n609), .B2(KEYINPUT77), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n602), .A2(new_n603), .B1(G85), .B2(new_n547), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(KEYINPUT77), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n535), .A2(G47), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT78), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(G290));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n540), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n522), .A2(new_n509), .A3(KEYINPUT10), .A4(G92), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n520), .B2(new_n521), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT79), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(new_n624), .C1(new_n512), .C2(new_n622), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n626), .A2(G651), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n532), .A2(G54), .A3(G543), .A4(new_n534), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n621), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G171), .B2(new_n632), .ZN(G284));
  OAI21_X1  g209(.A(new_n633), .B1(G171), .B2(new_n632), .ZN(G321));
  NAND2_X1  g210(.A1(G299), .A2(new_n632), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n632), .B2(G168), .ZN(G297));
  OAI21_X1  g212(.A(new_n636), .B1(new_n632), .B2(G168), .ZN(G280));
  INV_X1    g213(.A(new_n631), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n643), .A2(new_n644), .B1(new_n632), .B2(new_n557), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n488), .A2(G2104), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  INV_X1    g225(.A(G2100), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  AOI22_X1  g228(.A1(G123), .A2(new_n485), .B1(new_n488), .B2(G135), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n656));
  INV_X1    g231(.A(G111), .ZN(new_n657));
  AOI22_X1  g232(.A1(new_n655), .A2(new_n656), .B1(new_n657), .B2(G2105), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n656), .B2(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n652), .A2(new_n653), .A3(new_n662), .ZN(G156));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2427), .B(G2430), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT14), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT82), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n665), .B2(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2451), .B(G2454), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT16), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1341), .B(G1348), .ZN(new_n678));
  OAI21_X1  g253(.A(KEYINPUT83), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n674), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n682));
  INV_X1    g257(.A(new_n678), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G14), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n677), .B2(new_n678), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(G401));
  XOR2_X1   g263(.A(G2084), .B(G2090), .Z(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT84), .Z(new_n691));
  NOR2_X1   g266(.A1(G2072), .A2(G2078), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n442), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n689), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n693), .B(KEYINPUT17), .Z(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n691), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n689), .A3(new_n690), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT18), .Z(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n691), .A3(new_n689), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(new_n661), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G2100), .ZN(G227));
  XNOR2_X1  g278(.A(G1971), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT19), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n706));
  XOR2_X1   g281(.A(G1956), .B(G2474), .Z(new_n707));
  XOR2_X1   g282(.A(G1961), .B(G1966), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n705), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n706), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT20), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n707), .A2(new_n708), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(new_n709), .ZN(new_n715));
  MUX2_X1   g290(.A(new_n714), .B(new_n715), .S(new_n705), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n717), .B(G1986), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(new_n720), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(G1991), .B(G1996), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT86), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1981), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n722), .A2(new_n724), .A3(new_n728), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(G229));
  NAND3_X1  g307(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  INV_X1    g309(.A(new_n488), .ZN(new_n735));
  INV_X1    g310(.A(G139), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT95), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n484), .B2(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G33), .B(new_n740), .S(G29), .Z(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(G2072), .ZN(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G32), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n484), .A2(G105), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT96), .Z(new_n747));
  INV_X1    g322(.A(new_n485), .ZN(new_n748));
  INV_X1    g323(.A(G129), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  INV_X1    g327(.A(G141), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n735), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n745), .B1(new_n755), .B2(new_n744), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT98), .B(G28), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n744), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n762), .B1(new_n764), .B2(KEYINPUT99), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(KEYINPUT99), .B2(new_n764), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT31), .B(G11), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n660), .B2(new_n744), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n759), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n756), .B2(new_n758), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n742), .A2(new_n743), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n744), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT94), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(new_n484), .B2(G116), .ZN(new_n775));
  INV_X1    g350(.A(G104), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n484), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  AOI22_X1  g353(.A1(G128), .A2(new_n485), .B1(new_n488), .B2(G140), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(new_n744), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(G164), .A2(G29), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G27), .B2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G16), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G5), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G171), .B2(new_n789), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1961), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n785), .A2(new_n786), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n789), .A2(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n558), .B2(new_n789), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1341), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n788), .A2(new_n792), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n789), .A2(G4), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n639), .B2(new_n789), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1348), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n744), .A2(G35), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G162), .B2(new_n744), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT29), .Z(new_n803));
  INV_X1    g378(.A(G2090), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n789), .A2(G20), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G299), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1956), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n771), .A2(new_n797), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G34), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(KEYINPUT24), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(KEYINPUT24), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n744), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G160), .B2(new_n744), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2084), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n789), .A2(G21), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G168), .B2(new_n789), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  INV_X1    g395(.A(G1966), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n803), .B2(new_n804), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n811), .A2(new_n817), .A3(new_n823), .ZN(new_n824));
  MUX2_X1   g399(.A(G23), .B(G288), .S(G16), .Z(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(KEYINPUT91), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(KEYINPUT91), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT33), .B(G1976), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n826), .B2(new_n827), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n789), .A2(G22), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G166), .B2(new_n789), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(G1971), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n789), .A2(G6), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n597), .B2(new_n789), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT32), .B(G1981), .Z(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT90), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G1971), .B2(new_n832), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n829), .A2(new_n830), .A3(new_n833), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(G290), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G16), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G16), .B2(G24), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(new_n718), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n718), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n744), .A2(G25), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n484), .B2(G107), .ZN(new_n850));
  INV_X1    g425(.A(G95), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(new_n484), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT87), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n488), .A2(G131), .ZN(new_n854));
  INV_X1    g429(.A(G119), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n748), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n849), .B1(new_n857), .B2(new_n744), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT35), .B(G1991), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT88), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n858), .B(new_n860), .Z(new_n861));
  NOR3_X1   g436(.A1(new_n847), .A2(new_n848), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n842), .A2(new_n843), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n824), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT92), .B(KEYINPUT36), .Z(new_n866));
  AND2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(G311));
  OR2_X1    g443(.A1(new_n865), .A2(new_n867), .ZN(G150));
  NAND4_X1  g444(.A1(new_n532), .A2(G55), .A3(G543), .A4(new_n534), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n522), .A2(new_n509), .A3(G93), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n547), .A2(G81), .B1(new_n555), .B2(G651), .ZN(new_n873));
  INV_X1    g448(.A(G67), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n520), .B2(new_n521), .ZN(new_n875));
  NAND2_X1  g450(.A1(G80), .A2(G543), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT101), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(new_n876), .C1(new_n512), .C2(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(G651), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n872), .A2(new_n552), .A3(new_n873), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n878), .A2(G651), .A3(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n870), .A2(new_n871), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n557), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT38), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n639), .A2(G559), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n890));
  INV_X1    g465(.A(G860), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n883), .A2(new_n884), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(new_n891), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(G145));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n740), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n780), .B(new_n507), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n750), .B2(new_n754), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n780), .B(G164), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n755), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(G130), .A2(new_n485), .B1(new_n488), .B2(G142), .ZN(new_n905));
  OAI21_X1  g480(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n906));
  INV_X1    g481(.A(G118), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n906), .A2(KEYINPUT103), .B1(new_n907), .B2(G2105), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(KEYINPUT103), .B2(new_n906), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n649), .B(new_n910), .Z(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n899), .A2(new_n901), .A3(new_n903), .A4(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n740), .A2(new_n898), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(new_n857), .Z(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n913), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(G160), .B(G162), .Z(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(new_n660), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n920), .A3(new_n919), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n573), .A2(new_n581), .A3(new_n631), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n631), .B1(new_n573), .B2(new_n581), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G299), .A2(new_n639), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n573), .A2(new_n631), .A3(new_n581), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n935), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n642), .B(new_n886), .ZN(new_n941));
  MUX2_X1   g516(.A(new_n939), .B(new_n940), .S(new_n941), .Z(new_n942));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(G166), .B(G288), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n611), .A2(new_n615), .A3(G305), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G305), .B1(new_n611), .B2(new_n615), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  XNOR2_X1  g527(.A(G288), .B(G303), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n948), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n943), .B2(new_n944), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n942), .A2(new_n945), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n946), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n946), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(G868), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(G868), .B2(new_n894), .ZN(G295));
  OAI21_X1  g536(.A(new_n960), .B1(G868), .B2(new_n894), .ZN(G331));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  OAI21_X1  g539(.A(G286), .B1(G171), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n544), .A2(new_n964), .A3(new_n546), .A4(new_n548), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n882), .A2(new_n885), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n882), .B2(new_n885), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n886), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G168), .B1(G301), .B2(KEYINPUT106), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n882), .A2(new_n885), .A3(new_n966), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n969), .A2(new_n974), .A3(new_n940), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n969), .A2(new_n974), .B1(new_n938), .B2(new_n933), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n951), .A2(new_n954), .ZN(new_n978));
  AOI21_X1  g553(.A(G37), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n937), .B1(new_n931), .B2(new_n932), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n934), .A2(new_n930), .A3(new_n935), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n974), .B2(new_n969), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n955), .B1(new_n983), .B2(new_n975), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n963), .B1(new_n985), .B2(KEYINPUT43), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n955), .B1(new_n975), .B2(new_n976), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n969), .A2(new_n974), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n939), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n969), .A2(new_n974), .A3(new_n940), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n978), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n927), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n986), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n984), .A2(new_n994), .A3(new_n927), .A4(new_n991), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n995), .A2(KEYINPUT107), .B1(new_n992), .B2(KEYINPUT43), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n979), .A2(new_n997), .A3(new_n994), .A4(new_n984), .ZN(new_n998));
  AOI211_X1 g573(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(KEYINPUT107), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1003), .B2(new_n963), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n993), .B1(new_n999), .B2(new_n1004), .ZN(G397));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT109), .B(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(G164), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n479), .B1(new_n478), .B2(G2105), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n472), .A2(new_n473), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(KEYINPUT68), .A3(new_n484), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1010), .A2(G40), .A3(new_n1012), .A4(new_n469), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n780), .B(G2067), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n755), .B(G1996), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT110), .Z(new_n1019));
  XNOR2_X1  g594(.A(new_n857), .B(new_n860), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n844), .A2(new_n718), .A3(new_n1014), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n782), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n857), .A2(new_n860), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1021), .A2(new_n1023), .B1(new_n1026), .B2(new_n1014), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1015), .B1(new_n1016), .B2(new_n755), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT126), .Z(new_n1029));
  INV_X1    g604(.A(G1996), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1014), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT46), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT127), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1029), .A2(KEYINPUT47), .A3(new_n1032), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1027), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1036), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n481), .A3(G40), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  INV_X1    g620(.A(G1384), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1045), .B(KEYINPUT45), .C1(new_n507), .C2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n494), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n470), .B2(new_n471), .ZN(new_n1050));
  AOI21_X1  g625(.A(G2105), .B1(new_n1050), .B2(new_n496), .ZN(new_n1051));
  OAI21_X1  g626(.A(G126), .B1(new_n470), .B2(new_n471), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n484), .B1(new_n1052), .B2(new_n501), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1384), .B1(new_n1054), .B2(new_n506), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1045), .B1(new_n1055), .B2(KEYINPUT45), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1971), .B1(new_n1048), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n507), .B2(new_n1046), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(new_n1013), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n507), .A2(new_n1058), .A3(new_n1046), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT112), .B(G2090), .Z(new_n1062));
  AND3_X1   g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1042), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1008), .B1(new_n1054), .B2(new_n506), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1013), .B1(new_n1065), .B2(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n507), .A2(new_n1046), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(KEYINPUT111), .A3(new_n1006), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1056), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1971), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(KEYINPUT50), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1013), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1061), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1062), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(KEYINPUT113), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G166), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT55), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1064), .A2(G8), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(new_n1078), .B(KEYINPUT55), .Z(new_n1081));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1061), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n507), .A2(KEYINPUT116), .A3(new_n1058), .A4(new_n1046), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1013), .B(new_n1059), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1085), .A2(new_n1062), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1081), .B1(new_n1086), .B2(new_n1077), .ZN(new_n1087));
  OR3_X1    g662(.A1(new_n593), .A2(new_n596), .A3(G1981), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n1089));
  OAI21_X1  g664(.A(G1981), .B1(new_n593), .B2(new_n596), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  NAND3_X1  g667(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1073), .A2(new_n1055), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G8), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1067), .A2(new_n1013), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n1077), .ZN(new_n1100));
  INV_X1    g675(.A(G1976), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT52), .B1(G288), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1100), .B(new_n1102), .C1(new_n1101), .C2(G288), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G288), .A2(new_n1101), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT52), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1098), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1067), .A2(new_n1006), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1046), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1073), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n821), .ZN(new_n1111));
  INV_X1    g686(.A(G2084), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1060), .A2(new_n1112), .A3(new_n1061), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1077), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(G286), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1080), .A2(new_n1087), .A3(new_n1107), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1064), .A2(G8), .A3(new_n1076), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1081), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1115), .A2(new_n1118), .A3(G286), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1121), .A2(new_n1080), .A3(new_n1107), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1080), .A2(new_n1087), .A3(new_n1107), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1013), .B1(new_n1006), .B2(new_n1067), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1966), .B1(new_n1126), .B2(new_n1109), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1112), .A2(new_n1072), .A3(new_n1073), .A4(new_n1061), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT122), .B(G8), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G286), .A2(G8), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1114), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1135), .B(G8), .C1(new_n1136), .C2(G286), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(G8), .A3(G286), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT62), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(G1961), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(G2078), .ZN(new_n1143));
  AND4_X1   g718(.A1(new_n1073), .A2(new_n1108), .A3(new_n1143), .A4(new_n1109), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1056), .A2(new_n1066), .A3(new_n786), .A4(new_n1068), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1141), .B(new_n1144), .C1(new_n1142), .C2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT123), .B1(new_n1146), .B2(G301), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1141), .B1(new_n1145), .B2(new_n1142), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1143), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(new_n1110), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(G171), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1129), .B(new_n1130), .C1(new_n1114), .C2(new_n1132), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(new_n1138), .A4(new_n1137), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1125), .A2(new_n1140), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1080), .ZN(new_n1158));
  NOR2_X1   g733(.A1(G288), .A2(G1976), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT115), .Z(new_n1160));
  NOR2_X1   g735(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1088), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1158), .A2(new_n1107), .B1(new_n1100), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1124), .A2(new_n1157), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g741(.A1(G299), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n573), .A2(new_n581), .A3(KEYINPUT57), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT56), .B(G2072), .ZN(new_n1170));
  AND4_X1   g745(.A1(new_n1056), .A2(new_n1066), .A3(new_n1068), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1172));
  AOI21_X1  g747(.A(G1956), .B1(new_n1172), .B2(new_n1060), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1169), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1056), .A2(new_n1066), .A3(new_n1068), .A4(new_n1170), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1175), .B(new_n1176), .C1(new_n1085), .C2(G1956), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT119), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1178), .A2(KEYINPUT119), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1174), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1056), .A2(new_n1066), .A3(new_n1030), .A4(new_n1068), .ZN(new_n1185));
  XOR2_X1   g760(.A(KEYINPUT58), .B(G1341), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n1096), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n557), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n558), .ZN(new_n1192));
  NOR2_X1   g767(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1189), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1184), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1165), .B1(new_n1183), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1194), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1188), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1199), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1200), .A2(new_n1201), .A3(KEYINPUT120), .A4(new_n1184), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT117), .ZN(new_n1203));
  AOI21_X1  g778(.A(G1348), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1096), .A2(G2067), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1099), .A2(new_n782), .ZN(new_n1207));
  OAI211_X1 g782(.A(KEYINPUT117), .B(new_n1207), .C1(new_n1074), .C2(G1348), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT60), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1206), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT121), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1212), .A2(new_n1213), .A3(new_n639), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1213), .B1(new_n1212), .B2(new_n639), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1210), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1212), .A2(new_n639), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(KEYINPUT121), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1219), .A2(KEYINPUT60), .A3(new_n1209), .A4(new_n1214), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1197), .A2(new_n1202), .A3(new_n1217), .A4(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1174), .B1(new_n1209), .B2(new_n631), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1177), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1154), .A2(new_n1138), .A3(new_n1137), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1125), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1013), .B(KEYINPUT124), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1227), .A2(new_n1043), .A3(new_n1009), .A4(new_n1143), .ZN(new_n1228));
  AND2_X1   g803(.A1(new_n1148), .A2(new_n1228), .ZN(new_n1229));
  OR2_X1    g804(.A1(new_n1229), .A2(KEYINPUT125), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(KEYINPUT125), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1230), .A2(G171), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT54), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1233), .B1(new_n1150), .B2(G301), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g810(.A(KEYINPUT54), .B1(new_n1229), .B2(G301), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1236), .A2(new_n1152), .A3(new_n1147), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1226), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1164), .B1(new_n1224), .B2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g814(.A(G290), .B(new_n718), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1021), .B1(new_n1015), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g816(.A(new_n1041), .B1(new_n1239), .B2(new_n1241), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g817(.A1(G227), .A2(new_n460), .ZN(new_n1244));
  NAND3_X1  g818(.A1(new_n730), .A2(new_n731), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g819(.A(new_n1245), .B1(new_n685), .B2(new_n687), .ZN(new_n1246));
  AND3_X1   g820(.A1(new_n1246), .A2(new_n928), .A3(new_n1003), .ZN(G308));
  NAND3_X1  g821(.A1(new_n1246), .A2(new_n928), .A3(new_n1003), .ZN(G225));
endmodule


