//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n201), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G107), .C2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n202), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n209), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  NOR2_X1   g0031(.A1(G58), .A2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n234), .A2(new_n207), .A3(new_n235), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n228), .A2(new_n231), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT66), .B(G250), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n215), .ZN(new_n245));
  XOR2_X1   g0045(.A(G264), .B(G270), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  NOR2_X1   g0048(.A1(new_n201), .A2(new_n202), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n203), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT67), .ZN(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(G107), .B(G116), .Z(new_n255));
  XNOR2_X1  g0055(.A(G87), .B(G97), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  NAND2_X1  g0058(.A1(new_n225), .A2(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n259), .B1(G226), .B2(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G97), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n262), .B2(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n275), .B2(G238), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT13), .B1(new_n270), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n267), .ZN(new_n279));
  INV_X1    g0079(.A(new_n269), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(new_n265), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(new_n276), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n278), .A2(KEYINPUT73), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT73), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(KEYINPUT13), .C1(new_n270), .C2(new_n277), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G169), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n289), .A3(G169), .A4(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT74), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n278), .A2(new_n291), .A3(new_n283), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n281), .A2(KEYINPUT74), .A3(new_n282), .A4(new_n276), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G179), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n201), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n207), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n297), .B1(new_n298), .B2(new_n202), .C1(new_n300), .C2(new_n220), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n235), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(KEYINPUT11), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n201), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n206), .A2(G20), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT68), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n307), .A2(new_n303), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G68), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n305), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n304), .A2(KEYINPUT11), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n296), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n284), .A2(G200), .A3(new_n286), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n316), .A3(new_n315), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n292), .B2(new_n293), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n326));
  INV_X1    g0126(.A(G223), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n221), .A2(G1698), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n260), .C2(new_n261), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n280), .ZN(new_n334));
  INV_X1    g0134(.A(new_n273), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n269), .A2(G232), .A3(new_n271), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(G179), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n269), .B1(new_n331), .B2(new_n332), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n342), .A2(new_n273), .A3(new_n336), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n260), .A2(new_n261), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT7), .B1(new_n349), .B2(new_n207), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NOR4_X1   g0151(.A1(new_n260), .A2(new_n261), .A3(new_n351), .A4(G20), .ZN(new_n352));
  OAI21_X1  g0152(.A(G68), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G159), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n300), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(G58), .A2(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n356), .B2(new_n232), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT76), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(KEYINPUT76), .B(G20), .C1(new_n356), .C2(new_n232), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n348), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI211_X1 g0164(.A(KEYINPUT77), .B(KEYINPUT16), .C1(new_n353), .C2(new_n361), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n353), .A2(new_n361), .A3(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n303), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT8), .B(G58), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n306), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n313), .B2(new_n369), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(KEYINPUT18), .B(new_n347), .C1(new_n368), .C2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n364), .A2(new_n365), .ZN(new_n377));
  INV_X1    g0177(.A(new_n303), .ZN(new_n378));
  INV_X1    g0178(.A(new_n355), .ZN(new_n379));
  XNOR2_X1  g0179(.A(G58), .B(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT76), .B1(new_n380), .B2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(new_n360), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OR2_X1    g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n207), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n351), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n385), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n201), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n390), .B2(KEYINPUT16), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n372), .B1(new_n377), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n347), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n376), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n363), .B1(new_n383), .B2(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT77), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n362), .A2(new_n348), .A3(new_n363), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n371), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n399), .A2(KEYINPUT79), .A3(KEYINPUT18), .A4(new_n347), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n375), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n273), .B1(new_n333), .B2(new_n280), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT78), .B1(new_n403), .B2(new_n337), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n342), .A2(new_n340), .A3(new_n336), .A4(new_n273), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n343), .A2(new_n321), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n398), .A3(new_n371), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n408), .A2(new_n398), .A3(KEYINPUT17), .A4(new_n371), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n411), .A2(KEYINPUT80), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT80), .B1(new_n411), .B2(new_n412), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n401), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n384), .A2(new_n385), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G238), .A2(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n225), .C2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n280), .C1(G107), .C2(new_n416), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n335), .C1(new_n222), .C2(new_n274), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(G179), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n313), .A2(G77), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT15), .B(G87), .Z(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n298), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n369), .A2(new_n300), .B1(new_n207), .B2(new_n202), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n303), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n307), .A2(new_n202), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n420), .A2(new_n346), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n421), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n325), .A2(new_n326), .A3(new_n415), .A4(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G20), .B1(new_n233), .B2(G50), .ZN(new_n434));
  INV_X1    g0234(.A(G150), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(new_n435), .B2(new_n300), .C1(new_n298), .C2(new_n369), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n303), .B1(new_n220), .B2(new_n307), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n311), .A2(G50), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT69), .ZN(new_n439));
  INV_X1    g0239(.A(new_n312), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT9), .ZN(new_n442));
  AND2_X1   g0242(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n328), .A2(G222), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n416), .B(new_n444), .C1(new_n327), .C2(new_n328), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(new_n280), .C1(G77), .C2(new_n416), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n335), .C1(new_n221), .C2(new_n274), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n443), .B1(new_n447), .B2(G200), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n442), .B(new_n448), .C1(new_n321), .C2(new_n447), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n450));
  XOR2_X1   g0250(.A(new_n449), .B(new_n450), .Z(new_n451));
  OR2_X1    g0251(.A1(new_n447), .A2(G179), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n447), .A2(new_n346), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n441), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n420), .A2(new_n321), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT70), .ZN(new_n456));
  INV_X1    g0256(.A(new_n429), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT70), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n420), .B2(G200), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n456), .B(new_n457), .C1(new_n455), .C2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n451), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n433), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT82), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G33), .A3(G283), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT83), .ZN(new_n469));
  AND2_X1   g0269(.A1(G250), .A2(G1698), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n416), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n469), .B(new_n470), .C1(new_n260), .C2(new_n261), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n468), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G244), .B(new_n328), .C1(new_n260), .C2(new_n261), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n416), .A2(KEYINPUT4), .A3(G244), .A4(new_n328), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n280), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G45), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1), .ZN(new_n482));
  AND2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n485), .A2(new_n269), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G257), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n482), .B(G274), .C1(new_n484), .C2(new_n483), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n480), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n346), .ZN(new_n490));
  OAI21_X1  g0290(.A(G107), .B1(new_n350), .B2(new_n352), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT81), .B(G107), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OR2_X1    g0293(.A1(KEYINPUT6), .A2(G97), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n495), .A3(new_n494), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(G20), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n299), .A2(G77), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n491), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n303), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n306), .A2(G97), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n206), .A2(G33), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n306), .A2(new_n505), .A3(new_n235), .A4(new_n302), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(new_n214), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G179), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n480), .A2(new_n510), .A3(new_n487), .A4(new_n488), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n490), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT85), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT85), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n490), .A2(new_n509), .A3(new_n514), .A4(new_n511), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n480), .A2(G190), .A3(new_n487), .A4(new_n488), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n507), .B1(new_n501), .B2(new_n303), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n504), .ZN(new_n518));
  INV_X1    g0318(.A(new_n468), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n470), .B1(new_n260), .B2(new_n261), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT83), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n521), .B2(new_n472), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n477), .A3(new_n478), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(new_n280), .B1(G257), .B2(new_n486), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n402), .B1(new_n524), .B2(new_n488), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT84), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n489), .A2(G200), .ZN(new_n527));
  AOI211_X1 g0327(.A(new_n503), .B(new_n507), .C1(new_n501), .C2(new_n303), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n516), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n513), .A2(new_n515), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT88), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n213), .B1(new_n481), .B2(G1), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n206), .A2(G45), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n269), .B(new_n533), .C1(G274), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT86), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n328), .A2(G238), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G244), .A2(G1698), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n384), .A2(new_n385), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G33), .ZN(new_n541));
  INV_X1    g0341(.A(G116), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n537), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n210), .A2(G1698), .ZN(new_n545));
  AND2_X1   g0345(.A1(G244), .A2(G1698), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n545), .A2(new_n546), .B1(new_n260), .B2(new_n261), .ZN(new_n547));
  INV_X1    g0347(.A(new_n543), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(KEYINPUT86), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n536), .B1(new_n550), .B2(new_n280), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT87), .B1(new_n551), .B2(G190), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n539), .B1(new_n210), .B2(G1698), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n537), .B(new_n543), .C1(new_n416), .C2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT86), .B1(new_n547), .B2(new_n548), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n280), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(KEYINPUT87), .A3(G190), .A4(new_n535), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n532), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(G20), .B1(new_n384), .B2(new_n385), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G68), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n212), .ZN(new_n564));
  INV_X1    g0364(.A(new_n264), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(G20), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n264), .B2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n303), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n424), .A2(new_n307), .ZN(new_n570));
  INV_X1    g0370(.A(new_n506), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G87), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n551), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(G200), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n556), .A2(G190), .A3(new_n535), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(KEYINPUT88), .A3(new_n557), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n559), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n551), .A2(new_n510), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n569), .B(new_n570), .C1(new_n424), .C2(new_n506), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(G169), .C2(new_n551), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT22), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n560), .A2(new_n585), .A3(G87), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n207), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n207), .A2(G107), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT23), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n543), .A2(new_n207), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(KEYINPUT24), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n586), .A2(new_n588), .B1(new_n207), .B2(new_n543), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n591), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n303), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n486), .A2(G264), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n384), .A2(new_n385), .B1(new_n215), .B2(G1698), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n213), .A2(new_n328), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n600), .A2(new_n601), .B1(G33), .B2(G294), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n599), .B(new_n488), .C1(new_n269), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  INV_X1    g0404(.A(new_n603), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G190), .ZN(new_n606));
  INV_X1    g0406(.A(G107), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT25), .B1(new_n307), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n307), .A2(KEYINPUT25), .A3(new_n607), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n609), .A2(new_n610), .B1(G107), .B2(new_n571), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n598), .A2(new_n604), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n306), .A2(G116), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n506), .A2(new_n542), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n302), .A2(new_n235), .B1(G20), .B2(new_n542), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n207), .B1(new_n214), .B2(G33), .ZN(new_n616));
  OAI211_X1 g0416(.A(KEYINPUT20), .B(new_n615), .C1(new_n519), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT20), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n616), .B1(new_n465), .B2(new_n467), .ZN(new_n619));
  INV_X1    g0419(.A(new_n615), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n613), .B(new_n614), .C1(new_n617), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n328), .A2(G257), .ZN(new_n623));
  NAND2_X1  g0423(.A1(G264), .A2(G1698), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n623), .B(new_n624), .C1(new_n260), .C2(new_n261), .ZN(new_n625));
  INV_X1    g0425(.A(G303), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n384), .A2(new_n626), .A3(new_n385), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n280), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n485), .A2(G270), .A3(new_n269), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(G179), .A4(new_n488), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n488), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(KEYINPUT21), .A3(G169), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n622), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(G169), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n613), .B1(new_n617), .B2(new_n621), .ZN(new_n635));
  INV_X1    g0435(.A(new_n614), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT89), .B1(new_n637), .B2(KEYINPUT21), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT89), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n639), .B(new_n640), .C1(new_n622), .C2(new_n634), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n633), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n603), .A2(new_n346), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n605), .A2(new_n510), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n593), .A2(KEYINPUT24), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n596), .A2(new_n595), .A3(new_n591), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n378), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n611), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n643), .B(new_n644), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n631), .A2(G200), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n622), .B(new_n650), .C1(new_n321), .C2(new_n631), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n612), .A2(new_n642), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n463), .A2(new_n531), .A3(new_n584), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n454), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n394), .A2(new_n373), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n323), .A2(new_n432), .B1(new_n317), .B2(new_n296), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n413), .A2(new_n414), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n654), .B1(new_n658), .B2(new_n451), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n580), .A2(new_n513), .A3(new_n515), .A4(new_n583), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n578), .A2(new_n557), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n535), .B(KEYINPUT90), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n556), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G200), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT91), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n402), .B1(new_n556), .B2(new_n663), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT91), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n573), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n662), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n346), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n581), .A3(new_n582), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n670), .A2(new_n612), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n513), .A2(new_n515), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n526), .A2(new_n530), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n642), .A2(new_n649), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n672), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n512), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n661), .A2(new_n677), .A3(new_n681), .A4(new_n672), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n659), .B1(new_n462), .B2(new_n683), .ZN(G369));
  INV_X1    g0484(.A(G13), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G20), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n235), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT92), .ZN(new_n689));
  INV_X1    g0489(.A(G213), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n687), .B2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(KEYINPUT92), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G343), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT93), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n622), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(new_n642), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n651), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n695), .A2(new_n649), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n647), .A2(new_n648), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n612), .B1(new_n696), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n702), .B1(new_n704), .B2(new_n649), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n642), .A2(new_n695), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT94), .Z(new_n708));
  AOI21_X1  g0508(.A(new_n702), .B1(new_n708), .B2(new_n705), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n229), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G1), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n563), .A2(new_n212), .A3(new_n542), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(new_n234), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n652), .A2(new_n531), .A3(new_n584), .A4(new_n696), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n603), .A2(new_n630), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n524), .A3(new_n551), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n719), .A2(new_n524), .A3(KEYINPUT30), .A4(new_n551), .ZN(new_n723));
  AOI21_X1  g0523(.A(G179), .B1(new_n556), .B2(new_n663), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n489), .A2(new_n603), .A3(new_n631), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n695), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT31), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n729), .A3(new_n695), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n700), .B1(new_n718), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n682), .A2(new_n696), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n677), .A2(new_n672), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT26), .B1(new_n678), .B2(new_n512), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT29), .B(new_n696), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n732), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n717), .B1(new_n740), .B2(G1), .ZN(G364));
  INV_X1    g0541(.A(new_n701), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n714), .B1(G45), .B2(new_n686), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n699), .A2(new_n700), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n744), .B1(new_n699), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n235), .B1(G20), .B2(new_n346), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n207), .B1(new_n752), .B2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n214), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(new_n321), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G179), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n402), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n207), .A2(G190), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G179), .A3(new_n402), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n758), .A2(new_n220), .B1(new_n760), .B2(new_n202), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n756), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(G58), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n754), .B1(new_n763), .B2(KEYINPUT95), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(KEYINPUT95), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n402), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n759), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(G107), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n755), .A2(new_n766), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n212), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n759), .A2(G179), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n349), .B(new_n771), .C1(G68), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n759), .A2(new_n752), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n354), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  AND4_X1   g0577(.A1(new_n764), .A2(new_n769), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G294), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n753), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n760), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G311), .ZN(new_n782));
  INV_X1    g0582(.A(new_n762), .ZN(new_n783));
  INV_X1    g0583(.A(G322), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n349), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT96), .B(G326), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n780), .B(new_n785), .C1(new_n757), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  INV_X1    g0588(.A(new_n775), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n773), .A2(new_n788), .B1(new_n789), .B2(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n787), .B(new_n790), .C1(new_n791), .C2(new_n767), .ZN(new_n792));
  INV_X1    g0592(.A(new_n770), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(G303), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n751), .B1(new_n778), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n711), .A2(new_n349), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G355), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n254), .A2(new_n481), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n711), .A2(new_n416), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n234), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n797), .B1(G116), .B2(new_n229), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n749), .A2(new_n751), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n750), .A2(new_n795), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n746), .A2(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n696), .A2(new_n432), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n460), .B1(new_n696), .B2(new_n457), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n431), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n733), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n718), .A2(new_n731), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G330), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n810), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n744), .ZN(new_n814));
  INV_X1    g0614(.A(new_n809), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n747), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n751), .A2(new_n747), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n202), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n768), .A2(G68), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n224), .B2(new_n753), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n416), .B1(new_n775), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n762), .A2(G143), .B1(new_n773), .B2(G150), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n758), .C1(new_n354), .C2(new_n760), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n820), .B(new_n822), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n827), .B1(new_n826), .B2(new_n825), .C1(new_n220), .C2(new_n770), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G107), .A2(new_n793), .B1(new_n789), .B2(G311), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n829), .B1(new_n542), .B2(new_n760), .C1(new_n626), .C2(new_n758), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n754), .B(new_n830), .C1(G294), .C2(new_n762), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n212), .B2(new_n767), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n349), .B1(new_n835), .B2(new_n791), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n828), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n751), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n816), .A2(new_n743), .A3(new_n818), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n814), .A2(new_n839), .ZN(G384));
  NAND2_X1  g0640(.A1(new_n695), .A2(new_n317), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n296), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n324), .B2(new_n842), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n844), .A2(new_n811), .A3(new_n809), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n372), .B1(new_n391), .B2(new_n395), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n848), .A2(new_n693), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n415), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT100), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n415), .A2(KEYINPUT100), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n399), .A2(new_n347), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n399), .A2(new_n693), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n409), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n347), .A2(new_n693), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n848), .A2(new_n859), .B1(new_n408), .B2(new_n392), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n858), .B1(new_n860), .B2(new_n857), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n415), .A2(KEYINPUT100), .A3(new_n849), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT100), .B1(new_n415), .B2(new_n849), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT38), .B(new_n861), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n846), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n411), .A2(new_n412), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n655), .ZN(new_n871));
  INV_X1    g0671(.A(new_n856), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n855), .A2(new_n856), .A3(new_n409), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n871), .A2(new_n872), .B1(new_n874), .B2(new_n858), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT101), .B1(new_n875), .B2(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT101), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n874), .A2(new_n858), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n856), .B1(new_n870), .B2(new_n655), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n865), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(KEYINPUT40), .A3(new_n846), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n869), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT104), .Z(new_n886));
  NAND2_X1  g0686(.A1(new_n463), .A2(new_n811), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(G330), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n433), .A2(new_n461), .A3(new_n735), .A4(new_n739), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n659), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT102), .Z(new_n892));
  XNOR2_X1  g0692(.A(new_n889), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n878), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n883), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n318), .A2(new_n695), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n806), .B1(new_n733), .B2(new_n815), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n844), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT98), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(KEYINPUT98), .A3(new_n844), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n904), .B(new_n905), .C1(new_n866), .C2(new_n862), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n655), .A2(new_n693), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n893), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n206), .B2(new_n686), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n497), .A2(new_n498), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT35), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n207), .B(new_n235), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(G116), .C1(new_n914), .C2(new_n913), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT36), .ZN(new_n917));
  OAI21_X1  g0717(.A(G77), .B1(new_n224), .B2(new_n201), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n234), .A2(new_n918), .B1(G50), .B2(new_n201), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(G1), .A3(new_n685), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n912), .A2(new_n917), .A3(new_n920), .ZN(G367));
  AOI21_X1  g0721(.A(new_n206), .B1(new_n686), .B2(G45), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n531), .B1(new_n528), .B2(new_n696), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n696), .A2(new_n512), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n709), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT44), .Z(new_n928));
  INV_X1    g0728(.A(new_n706), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n709), .A2(new_n926), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT45), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n708), .B(new_n705), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n701), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n740), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n740), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n712), .B(KEYINPUT41), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n923), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n926), .A2(new_n708), .A3(new_n705), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT42), .Z(new_n943));
  INV_X1    g0743(.A(new_n926), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n674), .B1(new_n944), .B2(new_n649), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n696), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n695), .A2(new_n573), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n672), .A3(new_n670), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n672), .B2(new_n947), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n943), .A2(new_n946), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n706), .A2(new_n944), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n941), .A2(KEYINPUT105), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT105), .B1(new_n941), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n770), .A2(new_n224), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n767), .A2(new_n202), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n753), .A2(new_n201), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n757), .A2(G143), .B1(G137), .B2(new_n789), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n349), .B1(new_n781), .B2(G50), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n435), .B2(new_n783), .C1(new_n354), .C2(new_n835), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n783), .A2(new_n626), .B1(new_n753), .B2(new_n607), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G311), .B2(new_n757), .ZN(new_n967));
  INV_X1    g0767(.A(new_n835), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(G294), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n416), .B1(new_n781), .B2(G283), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G97), .A2(new_n768), .B1(new_n789), .B2(G317), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n967), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n770), .A2(new_n542), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT46), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n965), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n751), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n247), .A2(new_n799), .B1(new_n711), .B2(new_n423), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n744), .B1(new_n802), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT106), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT107), .Z(new_n982));
  INV_X1    g0782(.A(new_n749), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n949), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT108), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n957), .A2(new_n986), .ZN(G387));
  NOR2_X1   g0787(.A1(new_n705), .A2(new_n983), .ZN(new_n988));
  INV_X1    g0788(.A(new_n799), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n243), .B2(G45), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n715), .B2(new_n796), .ZN(new_n991));
  INV_X1    g0791(.A(new_n369), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n220), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT50), .ZN(new_n994));
  NOR4_X1   g0794(.A1(new_n994), .A2(G45), .A3(new_n249), .A4(new_n715), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n991), .A2(new_n995), .B1(G107), .B2(new_n229), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n802), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n743), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n424), .A2(new_n753), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G68), .B2(new_n781), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n354), .B2(new_n758), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n783), .A2(new_n220), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n770), .A2(new_n202), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n775), .A2(new_n435), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n768), .A2(G97), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n773), .A2(new_n992), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1005), .A2(new_n416), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n968), .A2(G311), .B1(G317), .B2(new_n762), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n626), .B2(new_n760), .C1(new_n784), .C2(new_n758), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n791), .B2(new_n753), .C1(new_n779), .C2(new_n770), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT49), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n789), .A2(new_n786), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n768), .A2(G116), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1014), .A2(new_n349), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1008), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n988), .B(new_n998), .C1(new_n1019), .C2(new_n751), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n923), .B2(new_n935), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n712), .B1(new_n935), .B2(new_n740), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1021), .B1(new_n937), .B2(new_n1022), .ZN(G393));
  NAND2_X1  g0823(.A1(new_n932), .A2(new_n933), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n936), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(new_n712), .A3(new_n938), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n932), .A2(new_n923), .A3(new_n933), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n416), .B1(new_n760), .B2(new_n369), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n753), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(G77), .B2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G87), .A2(new_n768), .B1(new_n789), .B2(G143), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n201), .C2(new_n770), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G150), .A2(new_n757), .B1(new_n762), .B2(G159), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT51), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(G50), .C2(new_n968), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n753), .A2(new_n542), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G311), .A2(new_n762), .B1(new_n757), .B2(G317), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  NAND2_X1  g0838(.A1(new_n968), .A2(G303), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G107), .A2(new_n768), .B1(new_n789), .B2(G322), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1038), .A2(new_n349), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1036), .B(new_n1041), .C1(G283), .C2(new_n793), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n781), .A2(G294), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT109), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n751), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n944), .A2(new_n749), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n802), .B1(new_n214), .B2(new_n229), .C1(new_n989), .C2(new_n257), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n743), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1026), .A2(new_n1027), .A3(new_n1049), .ZN(G390));
  INV_X1    g0850(.A(KEYINPUT112), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n844), .A2(new_n732), .A3(new_n809), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n899), .B1(new_n865), .B2(new_n882), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n808), .A2(new_n431), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n696), .B(new_n1054), .C1(new_n736), .C2(new_n738), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n806), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT110), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT110), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1058), .A3(new_n806), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n844), .A3(new_n1059), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1053), .A2(new_n1060), .A3(KEYINPUT111), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT111), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n899), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n896), .A2(new_n898), .B1(new_n1064), .B2(new_n902), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1051), .B(new_n1052), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1051), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n811), .A2(G330), .A3(new_n809), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n843), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n320), .A2(new_n322), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n317), .B2(new_n296), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1069), .B1(new_n1071), .B2(new_n841), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n896), .A2(new_n898), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n902), .A2(new_n1064), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(KEYINPUT112), .C1(new_n1062), .C2(new_n1061), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1067), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n901), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT113), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(new_n1073), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1068), .A2(new_n1080), .A3(new_n1072), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1079), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1055), .A2(new_n1058), .A3(new_n806), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1058), .B1(new_n1055), .B2(new_n806), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1052), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n815), .B1(new_n812), .B2(KEYINPUT114), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n732), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n844), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1088), .A2(new_n1092), .A3(KEYINPUT115), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT115), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1073), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n732), .A2(new_n1090), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n809), .B1(new_n732), .B2(new_n1090), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1072), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1094), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1085), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n433), .A2(G330), .A3(new_n461), .A4(new_n811), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n890), .A2(new_n1101), .A3(new_n659), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1100), .A2(KEYINPUT116), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT116), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT115), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1107), .A2(new_n1098), .A3(new_n1094), .A4(new_n1052), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1084), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1105), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1104), .A2(new_n1110), .A3(KEYINPUT117), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT117), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1066), .B(new_n1078), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1078), .A2(new_n1066), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n712), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1074), .A2(new_n747), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n771), .B1(new_n968), .B2(G107), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n781), .A2(G97), .B1(new_n1029), .B2(G77), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n819), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n775), .A2(new_n779), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n783), .A2(new_n542), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n349), .B1(new_n758), .B2(new_n791), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n349), .B1(new_n789), .B2(G125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n835), .B2(new_n824), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G128), .A2(new_n757), .B1(new_n762), .B2(G132), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n768), .A2(G50), .ZN(new_n1129));
  OR3_X1    g0929(.A1(new_n770), .A2(KEYINPUT53), .A3(new_n435), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT53), .B1(new_n770), .B2(new_n435), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n753), .A2(new_n354), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT54), .B(G143), .Z(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n760), .ZN(new_n1136));
  NOR4_X1   g0936(.A1(new_n1127), .A2(new_n1132), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n751), .B1(new_n1125), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1118), .A2(new_n743), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n369), .B2(new_n817), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1114), .B2(new_n923), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1117), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT118), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT118), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1117), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(G378));
  AOI21_X1  g0946(.A(new_n845), .B1(new_n895), .B2(new_n865), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n868), .ZN(new_n1148));
  OAI211_X1 g0948(.A(G330), .B(new_n884), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT119), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT119), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n869), .A2(new_n1151), .A3(G330), .A4(new_n884), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n451), .A2(new_n454), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n441), .A2(new_n693), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1150), .A2(new_n1152), .A3(new_n1158), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n909), .A2(KEYINPUT120), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1157), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1160), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n923), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n747), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n220), .B1(new_n260), .B2(G41), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n757), .A2(G125), .B1(new_n793), .B2(new_n1134), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n762), .A2(G128), .B1(G150), .B2(new_n1029), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n821), .B2(new_n772), .C1(new_n824), .C2(new_n760), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n768), .A2(G159), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G41), .B1(new_n789), .B2(G124), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(new_n541), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1167), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n423), .A2(new_n781), .B1(new_n768), .B2(G58), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n791), .B2(new_n775), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n783), .A2(new_n607), .ZN(new_n1180));
  INV_X1    g0980(.A(G41), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n772), .B2(new_n214), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1179), .A2(new_n960), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1003), .A2(new_n416), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n542), .C2(new_n758), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT58), .Z(new_n1186));
  OAI21_X1  g0986(.A(new_n751), .B1(new_n1177), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n817), .A2(new_n220), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1166), .A2(new_n743), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1165), .A2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1078), .A2(new_n1066), .B1(new_n1110), .B2(new_n1104), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1191), .A2(new_n1102), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n713), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1116), .A2(new_n1103), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT121), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n910), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1159), .A2(new_n1198), .A3(new_n910), .A4(new_n1161), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1195), .A2(new_n1202), .A3(KEYINPUT57), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1190), .B1(new_n1194), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n1109), .A2(new_n1102), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n940), .B(new_n1206), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT122), .Z(new_n1208));
  AOI22_X1  g1008(.A1(new_n762), .A2(G283), .B1(new_n781), .B2(G107), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n779), .B2(new_n758), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n770), .A2(new_n214), .B1(new_n775), .B2(new_n626), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1210), .A2(new_n999), .A3(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n959), .A2(new_n416), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT123), .Z(new_n1214));
  OAI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(new_n542), .C2(new_n835), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n349), .B1(new_n793), .B2(G159), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n224), .B2(new_n767), .C1(new_n435), .C2(new_n760), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G50), .B2(new_n1029), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n762), .A2(G137), .B1(G128), .B2(new_n789), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n821), .C2(new_n758), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n835), .A2(new_n1135), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT124), .Z(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n751), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n743), .B(new_n1224), .C1(new_n844), .C2(new_n748), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n201), .B2(new_n817), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1100), .B2(new_n923), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1208), .A2(new_n1227), .ZN(G381));
  NOR2_X1   g1028(.A1(G381), .A2(G384), .ZN(new_n1229));
  INV_X1    g1029(.A(G390), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n957), .A2(new_n986), .A3(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1231), .A2(G396), .A3(G393), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1142), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1229), .A2(new_n1232), .A3(new_n1233), .A4(new_n1204), .ZN(G407));
  INV_X1    g1034(.A(G343), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1204), .A2(new_n1233), .ZN(new_n1237));
  OAI21_X1  g1037(.A(G213), .B1(new_n1236), .B2(new_n1237), .ZN(G409));
  INV_X1    g1038(.A(KEYINPUT60), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1206), .B1(new_n1115), .B2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1240), .B(new_n712), .C1(new_n1239), .C2(new_n1206), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1227), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n814), .A3(new_n839), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(G384), .A3(new_n1227), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n690), .A2(G343), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G2897), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1243), .A2(new_n1244), .A3(new_n1247), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1102), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1193), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1203), .A2(new_n712), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1190), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1117), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1144), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1254), .B(new_n1255), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1195), .A2(new_n940), .A3(new_n1164), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1202), .A2(new_n923), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1189), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1233), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1246), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1245), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G387), .A2(G390), .ZN(new_n1270));
  XOR2_X1   g1070(.A(G393), .B(G396), .Z(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1231), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1270), .B2(new_n1231), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1246), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1245), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1266), .A2(new_n1269), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1250), .A2(new_n1265), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G378), .A2(new_n1204), .B1(new_n1233), .B2(new_n1261), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1283), .A2(new_n1246), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1285), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1277), .B2(new_n1245), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1282), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(KEYINPUT126), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1275), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1273), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(KEYINPUT127), .B(new_n1279), .C1(new_n1291), .C2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1267), .A2(new_n1285), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1277), .A2(new_n1245), .A3(new_n1287), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1290), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1296), .B1(new_n1301), .B2(new_n1266), .ZN(new_n1302));
  AND4_X1   g1102(.A1(new_n1266), .A2(new_n1269), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1298), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1297), .A2(new_n1304), .ZN(G405));
  OAI21_X1  g1105(.A(new_n1258), .B1(new_n1142), .B2(new_n1204), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1284), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1276), .ZN(G402));
endmodule


