

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n737), .B(n736), .ZN(n741) );
  NOR2_X1 U550 ( .A1(G543), .A2(G651), .ZN(n641) );
  NOR2_X1 U551 ( .A1(n526), .A2(n525), .ZN(G160) );
  NAND2_X1 U552 ( .A1(n1012), .A2(G29), .ZN(n515) );
  AND2_X1 U553 ( .A1(n699), .A2(G1996), .ZN(n674) );
  AND2_X1 U554 ( .A1(n725), .A2(n724), .ZN(n726) );
  INV_X1 U555 ( .A(KEYINPUT99), .ZN(n736) );
  INV_X1 U556 ( .A(n699), .ZN(n717) );
  XOR2_X1 U557 ( .A(KEYINPUT1), .B(n535), .Z(n638) );
  INV_X1 U558 ( .A(KEYINPUT83), .ZN(n533) );
  XNOR2_X1 U559 ( .A(n534), .B(n533), .ZN(G164) );
  AND2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U561 ( .A1(G113), .A2(n874), .ZN(n517) );
  INV_X1 U562 ( .A(G2105), .ZN(n521) );
  NOR2_X2 U563 ( .A1(G2104), .A2(n521), .ZN(n872) );
  NAND2_X1 U564 ( .A1(G125), .A2(n872), .ZN(n516) );
  NAND2_X1 U565 ( .A1(n517), .A2(n516), .ZN(n526) );
  XNOR2_X1 U566 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n519) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XNOR2_X2 U568 ( .A(n519), .B(n518), .ZN(n881) );
  NAND2_X1 U569 ( .A1(G137), .A2(n881), .ZN(n520) );
  XNOR2_X1 U570 ( .A(n520), .B(KEYINPUT66), .ZN(n524) );
  AND2_X1 U571 ( .A1(n521), .A2(G2104), .ZN(n878) );
  NAND2_X1 U572 ( .A1(G101), .A2(n878), .ZN(n522) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U575 ( .A1(G138), .A2(n881), .ZN(n528) );
  NAND2_X1 U576 ( .A1(G102), .A2(n878), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U578 ( .A1(G114), .A2(n874), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G126), .A2(n872), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n534) );
  AND2_X1 U582 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U583 ( .A(G132), .ZN(G219) );
  INV_X1 U584 ( .A(G82), .ZN(G220) );
  INV_X1 U585 ( .A(G69), .ZN(G235) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NOR2_X2 U587 ( .A1(G651), .A2(n622), .ZN(n637) );
  NAND2_X1 U588 ( .A1(G52), .A2(n637), .ZN(n537) );
  INV_X1 U589 ( .A(G651), .ZN(n538) );
  NOR2_X1 U590 ( .A1(G543), .A2(n538), .ZN(n535) );
  NAND2_X1 U591 ( .A1(G64), .A2(n638), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G90), .A2(n641), .ZN(n540) );
  NOR2_X1 U594 ( .A1(n622), .A2(n538), .ZN(n635) );
  NAND2_X1 U595 ( .A1(G77), .A2(n635), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U597 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U598 ( .A1(n543), .A2(n542), .ZN(G171) );
  NAND2_X1 U599 ( .A1(n641), .A2(G89), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n544), .B(KEYINPUT4), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G76), .A2(n635), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U603 ( .A(n547), .B(KEYINPUT5), .ZN(n552) );
  NAND2_X1 U604 ( .A1(G51), .A2(n637), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G63), .A2(n638), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n550), .Z(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n553), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(n554) );
  XNOR2_X1 U611 ( .A(KEYINPUT74), .B(n554), .ZN(G286) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n555), .B(KEYINPUT10), .ZN(n556) );
  XNOR2_X1 U614 ( .A(KEYINPUT68), .B(n556), .ZN(G223) );
  INV_X1 U615 ( .A(G223), .ZN(n819) );
  NAND2_X1 U616 ( .A1(n819), .A2(G567), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  NAND2_X1 U618 ( .A1(G56), .A2(n638), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n558), .B(KEYINPUT14), .ZN(n569) );
  NAND2_X1 U620 ( .A1(n637), .A2(G43), .ZN(n559) );
  XNOR2_X1 U621 ( .A(KEYINPUT71), .B(n559), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n635), .A2(G68), .ZN(n560) );
  XNOR2_X1 U623 ( .A(KEYINPUT69), .B(n560), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n641), .A2(G81), .ZN(n561) );
  XOR2_X1 U625 ( .A(n561), .B(KEYINPUT12), .Z(n562) );
  NOR2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT70), .B(n564), .Z(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT13), .B(n565), .Z(n566) );
  NOR2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n948) );
  INV_X1 U631 ( .A(G860), .ZN(n606) );
  OR2_X1 U632 ( .A1(n948), .A2(n606), .ZN(G153) );
  INV_X1 U633 ( .A(G171), .ZN(G301) );
  NAND2_X1 U634 ( .A1(G868), .A2(G301), .ZN(n580) );
  NAND2_X1 U635 ( .A1(G92), .A2(n641), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G66), .A2(n638), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n637), .A2(G54), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT72), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G79), .A2(n635), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT73), .B(n575), .Z(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT15), .B(n578), .Z(n890) );
  INV_X1 U645 ( .A(n890), .ZN(n953) );
  INV_X1 U646 ( .A(G868), .ZN(n655) );
  NAND2_X1 U647 ( .A1(n953), .A2(n655), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(G284) );
  NAND2_X1 U649 ( .A1(G53), .A2(n637), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G65), .A2(n638), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G91), .A2(n641), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G78), .A2(n635), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n939) );
  INV_X1 U656 ( .A(n939), .ZN(G299) );
  NAND2_X1 U657 ( .A1(G868), .A2(G286), .ZN(n588) );
  NAND2_X1 U658 ( .A1(G299), .A2(n655), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G297) );
  NAND2_X1 U660 ( .A1(n606), .A2(G559), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n589), .A2(n890), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U663 ( .A1(G868), .A2(n948), .ZN(n591) );
  XOR2_X1 U664 ( .A(KEYINPUT75), .B(n591), .Z(n594) );
  NAND2_X1 U665 ( .A1(G868), .A2(n890), .ZN(n592) );
  NOR2_X1 U666 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G99), .A2(n878), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G135), .A2(n881), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G111), .A2(n874), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n872), .A2(G123), .ZN(n597) );
  XOR2_X1 U673 ( .A(KEYINPUT18), .B(n597), .Z(n598) );
  NOR2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT76), .ZN(n989) );
  XNOR2_X1 U677 ( .A(G2096), .B(n989), .ZN(n603) );
  NOR2_X1 U678 ( .A1(G2100), .A2(n603), .ZN(n604) );
  XNOR2_X1 U679 ( .A(KEYINPUT77), .B(n604), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G559), .A2(n890), .ZN(n605) );
  XOR2_X1 U681 ( .A(n948), .B(n605), .Z(n652) );
  NAND2_X1 U682 ( .A1(n606), .A2(n652), .ZN(n614) );
  NAND2_X1 U683 ( .A1(G93), .A2(n641), .ZN(n608) );
  NAND2_X1 U684 ( .A1(G80), .A2(n635), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n637), .A2(G55), .ZN(n609) );
  XOR2_X1 U687 ( .A(KEYINPUT78), .B(n609), .Z(n610) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n638), .A2(G67), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n654) );
  XNOR2_X1 U691 ( .A(n614), .B(n654), .ZN(G145) );
  NAND2_X1 U692 ( .A1(G85), .A2(n641), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G47), .A2(n637), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G72), .A2(n635), .ZN(n617) );
  XNOR2_X1 U696 ( .A(KEYINPUT67), .B(n617), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n638), .A2(G60), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(G290) );
  NAND2_X1 U700 ( .A1(G49), .A2(n637), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G87), .A2(n622), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n638), .A2(n625), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n626) );
  XOR2_X1 U705 ( .A(KEYINPUT79), .B(n626), .Z(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G88), .A2(n641), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G75), .A2(n635), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G50), .A2(n637), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G62), .A2(n638), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(G166) );
  NAND2_X1 U714 ( .A1(n635), .A2(G73), .ZN(n636) );
  XNOR2_X1 U715 ( .A(KEYINPUT2), .B(n636), .ZN(n646) );
  NAND2_X1 U716 ( .A1(G48), .A2(n637), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G61), .A2(n638), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G86), .A2(n641), .ZN(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT80), .B(n642), .Z(n643) );
  NOR2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(G305) );
  XNOR2_X1 U723 ( .A(n939), .B(KEYINPUT19), .ZN(n648) );
  XNOR2_X1 U724 ( .A(G288), .B(G166), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U726 ( .A(n649), .B(G305), .Z(n650) );
  XNOR2_X1 U727 ( .A(G290), .B(n650), .ZN(n651) );
  XOR2_X1 U728 ( .A(n654), .B(n651), .Z(n891) );
  XNOR2_X1 U729 ( .A(n652), .B(n891), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n653), .A2(G868), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2078), .A2(G2084), .ZN(n658) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U735 ( .A1(G2090), .A2(n659), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(KEYINPUT21), .Z(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U738 ( .A1(G2072), .A2(n662), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U740 ( .A1(G120), .A2(G57), .ZN(n663) );
  NOR2_X1 U741 ( .A1(G235), .A2(n663), .ZN(n664) );
  XNOR2_X1 U742 ( .A(KEYINPUT82), .B(n664), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n665), .A2(G108), .ZN(n823) );
  NAND2_X1 U744 ( .A1(n823), .A2(G567), .ZN(n670) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U746 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U747 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U748 ( .A1(G96), .A2(n668), .ZN(n824) );
  NAND2_X1 U749 ( .A1(n824), .A2(G2106), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n670), .A2(n669), .ZN(n825) );
  NAND2_X1 U751 ( .A1(G661), .A2(G483), .ZN(n671) );
  NOR2_X1 U752 ( .A1(n825), .A2(n671), .ZN(n822) );
  NAND2_X1 U753 ( .A1(n822), .A2(G36), .ZN(G176) );
  INV_X1 U754 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U755 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n818) );
  NOR2_X1 U756 ( .A1(G164), .A2(G1384), .ZN(n673) );
  INV_X1 U757 ( .A(KEYINPUT64), .ZN(n672) );
  XNOR2_X1 U758 ( .A(n673), .B(n672), .ZN(n748) );
  NAND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n749) );
  NOR2_X4 U760 ( .A1(n748), .A2(n749), .ZN(n699) );
  XOR2_X1 U761 ( .A(n674), .B(KEYINPUT26), .Z(n676) );
  NAND2_X1 U762 ( .A1(n717), .A2(G1341), .ZN(n675) );
  NAND2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U764 ( .A1(n948), .A2(n677), .ZN(n683) );
  NAND2_X1 U765 ( .A1(n683), .A2(n890), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n717), .A2(G1348), .ZN(n678) );
  XNOR2_X1 U767 ( .A(n678), .B(KEYINPUT96), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n699), .A2(G2067), .ZN(n679) );
  NAND2_X1 U769 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n685) );
  OR2_X1 U771 ( .A1(n890), .A2(n683), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n699), .A2(G2072), .ZN(n686) );
  XNOR2_X1 U774 ( .A(KEYINPUT27), .B(n686), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT93), .B(G1956), .ZN(n917) );
  NOR2_X1 U776 ( .A1(n699), .A2(n917), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT94), .ZN(n688) );
  NOR2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U779 ( .A1(n939), .A2(n692), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n696) );
  NOR2_X1 U781 ( .A1(n939), .A2(n692), .ZN(n694) );
  XNOR2_X1 U782 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n693) );
  XNOR2_X1 U783 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U785 ( .A(KEYINPUT29), .B(n697), .ZN(n704) );
  XNOR2_X1 U786 ( .A(KEYINPUT25), .B(G2078), .ZN(n968) );
  NAND2_X1 U787 ( .A1(n699), .A2(n968), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n698), .B(KEYINPUT91), .ZN(n701) );
  NOR2_X1 U789 ( .A1(n699), .A2(G1961), .ZN(n700) );
  NOR2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n709) );
  NOR2_X1 U791 ( .A1(n709), .A2(G301), .ZN(n702) );
  XNOR2_X1 U792 ( .A(n702), .B(KEYINPUT92), .ZN(n703) );
  NOR2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n714) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n717), .ZN(n729) );
  INV_X1 U795 ( .A(n729), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n705), .A2(G8), .ZN(n706) );
  NAND2_X1 U797 ( .A1(G8), .A2(n717), .ZN(n771) );
  NOR2_X1 U798 ( .A1(G1966), .A2(n771), .ZN(n728) );
  OR2_X1 U799 ( .A1(n706), .A2(n728), .ZN(n707) );
  XNOR2_X1 U800 ( .A(KEYINPUT30), .B(n707), .ZN(n708) );
  NOR2_X1 U801 ( .A1(G168), .A2(n708), .ZN(n711) );
  AND2_X1 U802 ( .A1(G301), .A2(n709), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U804 ( .A(n712), .B(KEYINPUT31), .ZN(n713) );
  NOR2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n727) );
  INV_X1 U806 ( .A(n727), .ZN(n716) );
  AND2_X1 U807 ( .A1(G286), .A2(G8), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n725) );
  INV_X1 U809 ( .A(G8), .ZN(n723) );
  NOR2_X1 U810 ( .A1(G1971), .A2(n771), .ZN(n719) );
  NOR2_X1 U811 ( .A1(G2090), .A2(n717), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n720), .A2(G303), .ZN(n721) );
  XNOR2_X1 U814 ( .A(n721), .B(KEYINPUT98), .ZN(n722) );
  OR2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U816 ( .A(n726), .B(KEYINPUT32), .ZN(n734) );
  NOR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U818 ( .A1(G8), .A2(n729), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U820 ( .A(n732), .B(KEYINPUT97), .Z(n733) );
  NAND2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n770) );
  NOR2_X1 U822 ( .A1(G1976), .A2(G288), .ZN(n743) );
  NOR2_X1 U823 ( .A1(G1971), .A2(G303), .ZN(n735) );
  NOR2_X1 U824 ( .A1(n743), .A2(n735), .ZN(n944) );
  NAND2_X1 U825 ( .A1(n770), .A2(n944), .ZN(n737) );
  NAND2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n938) );
  INV_X1 U827 ( .A(n938), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n738), .A2(KEYINPUT33), .ZN(n739) );
  INV_X1 U829 ( .A(n771), .ZN(n742) );
  AND2_X1 U830 ( .A1(n739), .A2(n742), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  NAND2_X1 U834 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U835 ( .A(n747), .B(KEYINPUT100), .ZN(n763) );
  XOR2_X1 U836 ( .A(G1981), .B(G305), .Z(n956) );
  INV_X1 U837 ( .A(n748), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n813) );
  NAND2_X1 U839 ( .A1(G140), .A2(n881), .ZN(n752) );
  NAND2_X1 U840 ( .A1(G104), .A2(n878), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U842 ( .A(KEYINPUT34), .B(n753), .ZN(n759) );
  NAND2_X1 U843 ( .A1(G116), .A2(n874), .ZN(n755) );
  NAND2_X1 U844 ( .A1(G128), .A2(n872), .ZN(n754) );
  NAND2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U846 ( .A(KEYINPUT35), .B(n756), .Z(n757) );
  XNOR2_X1 U847 ( .A(KEYINPUT84), .B(n757), .ZN(n758) );
  NOR2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U849 ( .A(n760), .B(KEYINPUT36), .Z(n761) );
  XNOR2_X1 U850 ( .A(KEYINPUT85), .B(n761), .ZN(n887) );
  XNOR2_X1 U851 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NOR2_X1 U852 ( .A1(n887), .A2(n811), .ZN(n995) );
  NAND2_X1 U853 ( .A1(n813), .A2(n995), .ZN(n809) );
  AND2_X1 U854 ( .A1(n956), .A2(n809), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n779) );
  INV_X1 U856 ( .A(n809), .ZN(n777) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U858 ( .A(n764), .B(KEYINPUT90), .Z(n765) );
  XNOR2_X1 U859 ( .A(KEYINPUT24), .B(n765), .ZN(n766) );
  OR2_X1 U860 ( .A1(n771), .A2(n766), .ZN(n775) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n767) );
  XOR2_X1 U862 ( .A(KEYINPUT101), .B(n767), .Z(n768) );
  NAND2_X1 U863 ( .A1(G8), .A2(n768), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U866 ( .A(n773), .B(KEYINPUT102), .ZN(n774) );
  AND2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  OR2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n801) );
  XOR2_X1 U870 ( .A(G1986), .B(G290), .Z(n940) );
  NAND2_X1 U871 ( .A1(G131), .A2(n881), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G107), .A2(n874), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G95), .A2(n878), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G119), .A2(n872), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n864) );
  INV_X1 U878 ( .A(G1991), .ZN(n802) );
  NOR2_X1 U879 ( .A1(n864), .A2(n802), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G117), .A2(n874), .ZN(n787) );
  NAND2_X1 U881 ( .A1(G129), .A2(n872), .ZN(n786) );
  NAND2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U883 ( .A(KEYINPUT86), .B(n788), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n881), .A2(G141), .ZN(n789) );
  XOR2_X1 U885 ( .A(KEYINPUT88), .B(n789), .Z(n790) );
  NOR2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n795) );
  XOR2_X1 U887 ( .A(KEYINPUT87), .B(KEYINPUT38), .Z(n793) );
  NAND2_X1 U888 ( .A1(G105), .A2(n878), .ZN(n792) );
  XNOR2_X1 U889 ( .A(n793), .B(n792), .ZN(n794) );
  NAND2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U891 ( .A(n796), .B(KEYINPUT89), .Z(n862) );
  AND2_X1 U892 ( .A1(n862), .A2(G1996), .ZN(n797) );
  NOR2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n997) );
  NAND2_X1 U894 ( .A1(n940), .A2(n997), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n799), .A2(n813), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n816) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n862), .ZN(n999) );
  INV_X1 U898 ( .A(n997), .ZN(n806) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n803) );
  AND2_X1 U900 ( .A1(n802), .A2(n864), .ZN(n992) );
  NOR2_X1 U901 ( .A1(n803), .A2(n992), .ZN(n804) );
  XOR2_X1 U902 ( .A(KEYINPUT103), .B(n804), .Z(n805) );
  NOR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n999), .A2(n807), .ZN(n808) );
  XNOR2_X1 U905 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n887), .A2(n811), .ZN(n996) );
  NAND2_X1 U908 ( .A1(n812), .A2(n996), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n818), .B(n817), .ZN(G329) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U914 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(G188) );
  XNOR2_X1 U917 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XOR2_X1 U918 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G57), .ZN(G237) );
  NOR2_X1 U922 ( .A1(n824), .A2(n823), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n825), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2096), .B(G2678), .Z(n827) );
  XNOR2_X1 U926 ( .A(G2090), .B(KEYINPUT43), .ZN(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U928 ( .A(n828), .B(KEYINPUT42), .Z(n830) );
  XNOR2_X1 U929 ( .A(G2072), .B(G2067), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U931 ( .A(KEYINPUT106), .B(G2100), .Z(n832) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2084), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1991), .B(G1956), .Z(n836) );
  XNOR2_X1 U936 ( .A(G1981), .B(G1966), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U938 ( .A(G1986), .B(G1961), .Z(n838) );
  XNOR2_X1 U939 ( .A(G1976), .B(G1971), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U941 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U942 ( .A(G2474), .B(KEYINPUT107), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U944 ( .A(KEYINPUT41), .B(n843), .ZN(n844) );
  XOR2_X1 U945 ( .A(n844), .B(G1996), .Z(G229) );
  NAND2_X1 U946 ( .A1(n872), .A2(G124), .ZN(n846) );
  XNOR2_X1 U947 ( .A(KEYINPUT44), .B(KEYINPUT108), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G136), .A2(n881), .ZN(n848) );
  NAND2_X1 U950 ( .A1(G112), .A2(n874), .ZN(n847) );
  NAND2_X1 U951 ( .A1(n848), .A2(n847), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G100), .A2(n878), .ZN(n849) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(n849), .ZN(n850) );
  NOR2_X1 U954 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U955 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(KEYINPUT110), .B(n854), .Z(G162) );
  NAND2_X1 U957 ( .A1(G118), .A2(n874), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G130), .A2(n872), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G142), .A2(n881), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G106), .A2(n878), .ZN(n857) );
  NAND2_X1 U962 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U963 ( .A(n859), .B(KEYINPUT45), .Z(n860) );
  NOR2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n871) );
  XOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n866) );
  XNOR2_X1 U967 ( .A(n864), .B(KEYINPUT113), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U969 ( .A(n867), .B(n989), .Z(n869) );
  XNOR2_X1 U970 ( .A(G164), .B(G160), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n886) );
  NAND2_X1 U973 ( .A1(n872), .A2(G127), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(KEYINPUT112), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G115), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT47), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G103), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G139), .A2(n881), .ZN(n882) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n882), .ZN(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n1001) );
  XNOR2_X1 U983 ( .A(G162), .B(n1001), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U985 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U986 ( .A1(G37), .A2(n889), .ZN(G395) );
  XNOR2_X1 U987 ( .A(n890), .B(G286), .ZN(n894) );
  XNOR2_X1 U988 ( .A(G171), .B(n891), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n892), .B(n948), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U992 ( .A(G2451), .B(G2430), .Z(n897) );
  XNOR2_X1 U993 ( .A(G2438), .B(G2443), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n903) );
  XOR2_X1 U995 ( .A(G2435), .B(G2454), .Z(n899) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U998 ( .A(G2446), .B(G2427), .Z(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n903), .B(n902), .Z(n904) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n904), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n910), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(n910), .ZN(G401) );
  XNOR2_X1 U1010 ( .A(KEYINPUT123), .B(G1981), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n911), .B(G6), .ZN(n916) );
  XOR2_X1 U1012 ( .A(G1348), .B(KEYINPUT59), .Z(n912) );
  XNOR2_X1 U1013 ( .A(G4), .B(n912), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(G19), .B(G1341), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n920) );
  XOR2_X1 U1017 ( .A(KEYINPUT122), .B(n917), .Z(n918) );
  XNOR2_X1 U1018 ( .A(G20), .B(n918), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(KEYINPUT60), .B(n921), .ZN(n931) );
  XNOR2_X1 U1021 ( .A(G1966), .B(KEYINPUT124), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(G21), .ZN(n929) );
  XNOR2_X1 U1023 ( .A(G1976), .B(G23), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G1971), .B(G22), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n926) );
  XOR2_X1 U1026 ( .A(G1986), .B(G24), .Z(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT58), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(G5), .B(G1961), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT61), .B(n934), .Z(n935) );
  NOR2_X1 U1034 ( .A1(G16), .A2(n935), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(KEYINPUT125), .B(n936), .ZN(n964) );
  XNOR2_X1 U1036 ( .A(KEYINPUT56), .B(G16), .ZN(n962) );
  NAND2_X1 U1037 ( .A1(G1971), .A2(G303), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n939), .B(G1956), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT121), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G1961), .B(KEYINPUT120), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(n947), .B(G301), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G1341), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G1348), .B(n953), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n958), .B(KEYINPUT57), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(n965), .B(KEYINPUT126), .ZN(n1015) );
  XOR2_X1 U1058 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n988) );
  INV_X1 U1059 ( .A(G29), .ZN(n986) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(G34), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(G2084), .B(n967), .ZN(n984) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G35), .ZN(n982) );
  XOR2_X1 U1064 ( .A(n968), .B(G27), .Z(n970) );
  XNOR2_X1 U1065 ( .A(G1996), .B(G32), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(KEYINPUT118), .B(n971), .ZN(n977) );
  XOR2_X1 U1068 ( .A(G2072), .B(G33), .Z(n972) );
  NAND2_X1 U1069 ( .A1(n972), .A2(G28), .ZN(n975) );
  XOR2_X1 U1070 ( .A(G25), .B(G1991), .Z(n973) );
  XNOR2_X1 U1071 ( .A(KEYINPUT117), .B(n973), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(G26), .B(G2067), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n980), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n988), .B(n987), .ZN(n1013) );
  XNOR2_X1 U1081 ( .A(G160), .B(G2084), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT115), .B(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1010) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1008) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(KEYINPUT51), .B(n1000), .Z(n1006) );
  XOR2_X1 U1090 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1013), .A2(n515), .ZN(n1014) );
  NOR2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(G11), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(n1017), .B(KEYINPUT62), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1018), .ZN(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

