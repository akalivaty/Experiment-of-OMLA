

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n527), .A2(n526), .ZN(n529) );
  INV_X1 U558 ( .A(n700), .ZN(n725) );
  AND2_X1 U559 ( .A1(n698), .A2(n790), .ZN(n699) );
  XNOR2_X1 U560 ( .A(n697), .B(KEYINPUT93), .ZN(n790) );
  NOR2_X4 U561 ( .A1(G2104), .A2(n535), .ZN(n613) );
  BUF_X1 U562 ( .A(n896), .Z(n524) );
  XNOR2_X1 U563 ( .A(n529), .B(n528), .ZN(n896) );
  AND2_X1 U564 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U565 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U566 ( .A(n713), .B(KEYINPUT27), .ZN(n714) );
  NAND2_X1 U567 ( .A1(n696), .A2(G160), .ZN(n700) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n652) );
  AND2_X2 U569 ( .A1(n535), .A2(G2104), .ZN(n899) );
  INV_X1 U570 ( .A(G2105), .ZN(n527) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NOR2_X1 U572 ( .A1(n775), .A2(n768), .ZN(n525) );
  INV_X1 U573 ( .A(KEYINPUT30), .ZN(n703) );
  INV_X1 U574 ( .A(KEYINPUT29), .ZN(n738) );
  XNOR2_X1 U575 ( .A(n739), .B(n738), .ZN(n742) );
  INV_X1 U576 ( .A(KEYINPUT103), .ZN(n771) );
  NOR2_X1 U577 ( .A1(G164), .A2(G1384), .ZN(n816) );
  INV_X1 U578 ( .A(G2104), .ZN(n526) );
  XNOR2_X1 U579 ( .A(n577), .B(KEYINPUT13), .ZN(n578) );
  INV_X1 U580 ( .A(KEYINPUT17), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n579), .B(n578), .ZN(n582) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(n540), .ZN(n648) );
  NOR2_X1 U583 ( .A1(G651), .A2(n661), .ZN(n655) );
  NAND2_X1 U584 ( .A1(n584), .A2(n583), .ZN(n1036) );
  NAND2_X1 U585 ( .A1(G137), .A2(n896), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n530), .B(KEYINPUT65), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G113), .A2(n892), .ZN(n532) );
  INV_X1 U588 ( .A(G2105), .ZN(n535) );
  NAND2_X1 U589 ( .A1(G125), .A2(n613), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G101), .A2(n899), .ZN(n536) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(n536), .Z(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X2 U595 ( .A(n539), .B(KEYINPUT64), .Z(G160) );
  INV_X1 U596 ( .A(G651), .ZN(n547) );
  XOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .Z(n661) );
  OR2_X1 U598 ( .A1(n547), .A2(n661), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n648), .A2(G76), .ZN(n541) );
  XNOR2_X1 U600 ( .A(KEYINPUT78), .B(n541), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT4), .B(KEYINPUT77), .Z(n543) );
  NAND2_X1 U602 ( .A1(G89), .A2(n652), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U605 ( .A(n546), .B(KEYINPUT5), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G51), .A2(n655), .ZN(n550) );
  NOR2_X1 U607 ( .A1(G543), .A2(n547), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT1), .B(n548), .Z(n659) );
  NAND2_X1 U609 ( .A1(G63), .A2(n659), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U613 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U614 ( .A1(n652), .A2(G90), .ZN(n555) );
  XOR2_X1 U615 ( .A(KEYINPUT69), .B(n555), .Z(n557) );
  NAND2_X1 U616 ( .A1(n648), .A2(G77), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n558), .B(KEYINPUT9), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G64), .A2(n659), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n655), .A2(G52), .ZN(n561) );
  XOR2_X1 U622 ( .A(KEYINPUT68), .B(n561), .Z(n562) );
  NOR2_X1 U623 ( .A1(n563), .A2(n562), .ZN(G171) );
  INV_X1 U624 ( .A(G171), .ZN(G301) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U626 ( .A(G120), .ZN(G236) );
  INV_X1 U627 ( .A(G69), .ZN(G235) );
  INV_X1 U628 ( .A(G108), .ZN(G238) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  NAND2_X1 U631 ( .A1(G138), .A2(n896), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G102), .A2(n899), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G114), .A2(n892), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G126), .A2(n613), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U637 ( .A(KEYINPUT89), .B(n568), .Z(n569) );
  NOR2_X1 U638 ( .A1(n570), .A2(n569), .ZN(G164) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n573) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n571) );
  XOR2_X1 U642 ( .A(n571), .B(KEYINPUT10), .Z(n844) );
  NAND2_X1 U643 ( .A1(G567), .A2(n844), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n573), .B(n572), .ZN(G234) );
  NAND2_X1 U645 ( .A1(n652), .A2(G81), .ZN(n574) );
  XNOR2_X1 U646 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U647 ( .A1(G68), .A2(n648), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n579) );
  XNOR2_X1 U649 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n659), .A2(G56), .ZN(n580) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n580), .Z(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n655), .A2(G43), .ZN(n583) );
  INV_X1 U654 ( .A(G860), .ZN(n607) );
  OR2_X1 U655 ( .A1(n1036), .A2(n607), .ZN(G153) );
  NAND2_X1 U656 ( .A1(G79), .A2(n648), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G92), .A2(n652), .ZN(n586) );
  NAND2_X1 U658 ( .A1(G66), .A2(n659), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G54), .A2(n655), .ZN(n587) );
  XNOR2_X1 U661 ( .A(KEYINPUT75), .B(n587), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U664 ( .A(n592), .B(KEYINPUT15), .Z(n1016) );
  INV_X1 U665 ( .A(G868), .ZN(n604) );
  NAND2_X1 U666 ( .A1(n1016), .A2(n604), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT76), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U670 ( .A1(n652), .A2(G91), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n596), .B(KEYINPUT70), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G78), .A2(n648), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U674 ( .A(KEYINPUT71), .B(n599), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n655), .A2(G53), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G65), .A2(n659), .ZN(n600) );
  AND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(G299) );
  NOR2_X1 U679 ( .A1(G286), .A2(n604), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n607), .A2(G559), .ZN(n608) );
  INV_X1 U683 ( .A(n1016), .ZN(n915) );
  NAND2_X1 U684 ( .A1(n608), .A2(n915), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n1036), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G868), .A2(n915), .ZN(n610) );
  NOR2_X1 U688 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G123), .A2(n613), .ZN(n614) );
  XOR2_X1 U691 ( .A(KEYINPUT18), .B(n614), .Z(n615) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT79), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G111), .A2(n892), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G135), .A2(n524), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G99), .A2(n899), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n950) );
  XNOR2_X1 U699 ( .A(n950), .B(G2096), .ZN(n622) );
  INV_X1 U700 ( .A(G2100), .ZN(n853) );
  NAND2_X1 U701 ( .A1(n622), .A2(n853), .ZN(G156) );
  NAND2_X1 U702 ( .A1(n915), .A2(G559), .ZN(n671) );
  XNOR2_X1 U703 ( .A(n1036), .B(n671), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n623), .A2(G860), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G55), .A2(n655), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G67), .A2(n659), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G93), .A2(n652), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G80), .A2(n648), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n674) );
  XNOR2_X1 U712 ( .A(n630), .B(n674), .ZN(G145) );
  NAND2_X1 U713 ( .A1(G60), .A2(n659), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G72), .A2(n648), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n652), .A2(G85), .ZN(n633) );
  XOR2_X1 U717 ( .A(KEYINPUT66), .B(n633), .Z(n634) );
  NOR2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n655), .A2(G47), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(G290) );
  NAND2_X1 U721 ( .A1(G50), .A2(n655), .ZN(n638) );
  XNOR2_X1 U722 ( .A(n638), .B(KEYINPUT82), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G62), .A2(n659), .ZN(n639) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n639), .Z(n640) );
  NAND2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G88), .A2(n652), .ZN(n643) );
  NAND2_X1 U727 ( .A1(G75), .A2(n648), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(G166) );
  INV_X1 U730 ( .A(G166), .ZN(G303) );
  NAND2_X1 U731 ( .A1(G48), .A2(n655), .ZN(n647) );
  NAND2_X1 U732 ( .A1(G61), .A2(n659), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U734 ( .A1(G73), .A2(n648), .ZN(n649) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(n649), .Z(n650) );
  NOR2_X1 U736 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n652), .A2(G86), .ZN(n653) );
  NAND2_X1 U738 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U739 ( .A1(G49), .A2(n655), .ZN(n657) );
  NAND2_X1 U740 ( .A1(G74), .A2(G651), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n660), .B(KEYINPUT80), .ZN(n663) );
  NAND2_X1 U744 ( .A1(G87), .A2(n661), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n663), .A2(n662), .ZN(G288) );
  XNOR2_X1 U746 ( .A(KEYINPUT83), .B(n1036), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n664), .B(G290), .ZN(n665) );
  XOR2_X1 U748 ( .A(n665), .B(KEYINPUT19), .Z(n667) );
  XOR2_X1 U749 ( .A(G303), .B(n674), .Z(n666) );
  XNOR2_X1 U750 ( .A(n667), .B(n666), .ZN(n670) );
  XOR2_X1 U751 ( .A(G299), .B(G305), .Z(n668) );
  XNOR2_X1 U752 ( .A(n668), .B(G288), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n670), .B(n669), .ZN(n916) );
  XNOR2_X1 U754 ( .A(n916), .B(n671), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n672), .A2(G868), .ZN(n673) );
  XOR2_X1 U756 ( .A(KEYINPUT84), .B(n673), .Z(n676) );
  NOR2_X1 U757 ( .A1(n674), .A2(G868), .ZN(n675) );
  NOR2_X1 U758 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U759 ( .A(KEYINPUT85), .B(n677), .ZN(G295) );
  XOR2_X1 U760 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n679) );
  NAND2_X1 U761 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XNOR2_X1 U762 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U769 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G96), .A2(n685), .ZN(n849) );
  NAND2_X1 U771 ( .A1(n849), .A2(G2106), .ZN(n691) );
  NOR2_X1 U772 ( .A1(G235), .A2(G236), .ZN(n686) );
  XNOR2_X1 U773 ( .A(n686), .B(KEYINPUT87), .ZN(n687) );
  NOR2_X1 U774 ( .A1(G238), .A2(n687), .ZN(n688) );
  NAND2_X1 U775 ( .A1(G57), .A2(n688), .ZN(n848) );
  NAND2_X1 U776 ( .A1(G567), .A2(n848), .ZN(n689) );
  XNOR2_X1 U777 ( .A(KEYINPUT88), .B(n689), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n850) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n850), .A2(n692), .ZN(n847) );
  NAND2_X1 U781 ( .A1(n847), .A2(G36), .ZN(G176) );
  INV_X1 U782 ( .A(G1966), .ZN(n698) );
  INV_X1 U783 ( .A(G40), .ZN(n695) );
  INV_X1 U784 ( .A(n816), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n700), .A2(G8), .ZN(n697) );
  XNOR2_X1 U787 ( .A(KEYINPUT94), .B(n699), .ZN(n746) );
  INV_X1 U788 ( .A(G8), .ZN(n701) );
  INV_X1 U789 ( .A(n725), .ZN(n750) );
  NOR2_X1 U790 ( .A1(G2084), .A2(n750), .ZN(n747) );
  OR2_X1 U791 ( .A1(n701), .A2(n747), .ZN(n702) );
  NOR2_X1 U792 ( .A1(n746), .A2(n702), .ZN(n704) );
  XNOR2_X1 U793 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U794 ( .A1(n705), .A2(G168), .ZN(n710) );
  XOR2_X1 U795 ( .A(KEYINPUT25), .B(G2078), .Z(n970) );
  NOR2_X1 U796 ( .A1(n970), .A2(n750), .ZN(n707) );
  XOR2_X1 U797 ( .A(G1961), .B(KEYINPUT95), .Z(n991) );
  NOR2_X1 U798 ( .A1(n725), .A2(n991), .ZN(n706) );
  NOR2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n740) );
  NAND2_X1 U800 ( .A1(n740), .A2(G301), .ZN(n708) );
  XOR2_X1 U801 ( .A(KEYINPUT100), .B(n708), .Z(n709) );
  NOR2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U803 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n711) );
  XNOR2_X1 U804 ( .A(n712), .B(n711), .ZN(n755) );
  INV_X1 U805 ( .A(G299), .ZN(n733) );
  NAND2_X1 U806 ( .A1(G2072), .A2(n725), .ZN(n713) );
  XNOR2_X1 U807 ( .A(n714), .B(KEYINPUT96), .ZN(n716) );
  INV_X1 U808 ( .A(G1956), .ZN(n1022) );
  NOR2_X1 U809 ( .A1(n725), .A2(n1022), .ZN(n715) );
  NOR2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n732) );
  NOR2_X1 U811 ( .A1(n733), .A2(n732), .ZN(n718) );
  XNOR2_X1 U812 ( .A(KEYINPUT28), .B(KEYINPUT97), .ZN(n717) );
  XNOR2_X1 U813 ( .A(n718), .B(n717), .ZN(n737) );
  XNOR2_X1 U814 ( .A(KEYINPUT98), .B(G1996), .ZN(n963) );
  NAND2_X1 U815 ( .A1(n963), .A2(n725), .ZN(n719) );
  XNOR2_X1 U816 ( .A(n719), .B(KEYINPUT26), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n750), .A2(G1341), .ZN(n720) );
  NAND2_X1 U818 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U819 ( .A1(n1036), .A2(n722), .ZN(n723) );
  OR2_X1 U820 ( .A1(n915), .A2(n723), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n915), .A2(n723), .ZN(n729) );
  AND2_X1 U822 ( .A1(n750), .A2(G1348), .ZN(n724) );
  XNOR2_X1 U823 ( .A(n724), .B(KEYINPUT99), .ZN(n727) );
  NAND2_X1 U824 ( .A1(n725), .A2(G2067), .ZN(n726) );
  NAND2_X1 U825 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U826 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n735) );
  NAND2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n739) );
  OR2_X1 U831 ( .A1(n740), .A2(G301), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n754) );
  NAND2_X1 U833 ( .A1(n755), .A2(n754), .ZN(n744) );
  INV_X1 U834 ( .A(KEYINPUT102), .ZN(n743) );
  XNOR2_X1 U835 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n749) );
  NAND2_X1 U837 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n764) );
  INV_X1 U839 ( .A(n790), .ZN(n775) );
  NOR2_X1 U840 ( .A1(G1971), .A2(n775), .ZN(n752) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n750), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n753), .A2(G303), .ZN(n757) );
  AND2_X1 U844 ( .A1(n754), .A2(n757), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n761) );
  INV_X1 U846 ( .A(n757), .ZN(n758) );
  OR2_X1 U847 ( .A1(n758), .A2(G286), .ZN(n759) );
  AND2_X1 U848 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U850 ( .A(n762), .B(KEYINPUT32), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n781) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n773) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n773), .A2(n765), .ZN(n1021) );
  INV_X1 U855 ( .A(KEYINPUT33), .ZN(n766) );
  AND2_X1 U856 ( .A1(n1021), .A2(n766), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n781), .A2(n767), .ZN(n770) );
  NAND2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n1020) );
  INV_X1 U859 ( .A(n1020), .ZN(n768) );
  OR2_X1 U860 ( .A1(KEYINPUT33), .A2(n525), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n772) );
  XNOR2_X1 U862 ( .A(n772), .B(n771), .ZN(n778) );
  NAND2_X1 U863 ( .A1(KEYINPUT33), .A2(n773), .ZN(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U865 ( .A(KEYINPUT104), .B(n776), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT105), .ZN(n780) );
  XNOR2_X1 U867 ( .A(G1981), .B(G305), .ZN(n1031) );
  NOR2_X1 U868 ( .A1(n780), .A2(n1031), .ZN(n787) );
  INV_X1 U869 ( .A(n781), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G166), .A2(G8), .ZN(n782) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n782), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n790), .A2(n785), .ZN(n786) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n788), .B(KEYINPUT106), .ZN(n831) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(KEYINPUT24), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n829) );
  NAND2_X1 U879 ( .A1(G105), .A2(n899), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n792), .B(KEYINPUT38), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n892), .A2(G117), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G129), .A2(n613), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G141), .A2(n524), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n888) );
  NOR2_X1 U887 ( .A1(G1996), .A2(n888), .ZN(n939) );
  XOR2_X1 U888 ( .A(KEYINPUT91), .B(G1991), .Z(n964) );
  NAND2_X1 U889 ( .A1(G95), .A2(n899), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n799), .B(KEYINPUT90), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n892), .A2(G107), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G119), .A2(n613), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G131), .A2(n524), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n906) );
  NOR2_X1 U897 ( .A1(n964), .A2(n906), .ZN(n951) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n806) );
  XOR2_X1 U899 ( .A(n806), .B(KEYINPUT107), .Z(n807) );
  NOR2_X1 U900 ( .A1(n951), .A2(n807), .ZN(n811) );
  AND2_X1 U901 ( .A1(n906), .A2(n964), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(KEYINPUT92), .ZN(n810) );
  AND2_X1 U903 ( .A1(G1996), .A2(n888), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n833) );
  INV_X1 U905 ( .A(n833), .ZN(n954) );
  NOR2_X1 U906 ( .A1(n811), .A2(n954), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n939), .A2(n812), .ZN(n813) );
  XNOR2_X1 U908 ( .A(n813), .B(KEYINPUT108), .ZN(n814) );
  XNOR2_X1 U909 ( .A(n814), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G40), .A2(G160), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n838) );
  NAND2_X1 U912 ( .A1(n817), .A2(n838), .ZN(n828) );
  XOR2_X1 U913 ( .A(G2067), .B(KEYINPUT37), .Z(n837) );
  NAND2_X1 U914 ( .A1(G140), .A2(n524), .ZN(n819) );
  NAND2_X1 U915 ( .A1(G104), .A2(n899), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U917 ( .A(KEYINPUT34), .B(n820), .ZN(n825) );
  NAND2_X1 U918 ( .A1(G116), .A2(n892), .ZN(n822) );
  NAND2_X1 U919 ( .A1(G128), .A2(n613), .ZN(n821) );
  NAND2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U921 ( .A(KEYINPUT35), .B(n823), .Z(n824) );
  NOR2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U923 ( .A(KEYINPUT36), .B(n826), .Z(n912) );
  NOR2_X1 U924 ( .A1(n837), .A2(n912), .ZN(n942) );
  NAND2_X1 U925 ( .A1(n942), .A2(n838), .ZN(n827) );
  AND2_X1 U926 ( .A1(n828), .A2(n827), .ZN(n832) );
  AND2_X1 U927 ( .A1(n829), .A2(n832), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n842) );
  INV_X1 U929 ( .A(n832), .ZN(n836) );
  XOR2_X1 U930 ( .A(G1986), .B(G290), .Z(n1015) );
  NAND2_X1 U931 ( .A1(n1015), .A2(n833), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n834), .A2(n838), .ZN(n835) );
  OR2_X1 U933 ( .A1(n836), .A2(n835), .ZN(n840) );
  AND2_X1 U934 ( .A1(n837), .A2(n912), .ZN(n937) );
  NAND2_X1 U935 ( .A1(n937), .A2(n838), .ZN(n839) );
  AND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n843), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n844), .ZN(G217) );
  INV_X1 U939 ( .A(n844), .ZN(G223) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U941 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U945 ( .A(G96), .ZN(G221) );
  NOR2_X1 U946 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  INV_X1 U948 ( .A(n850), .ZN(G319) );
  XOR2_X1 U949 ( .A(KEYINPUT109), .B(G2084), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n856) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2072), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(G2096), .B(G2678), .Z(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n860), .B(n859), .Z(G227) );
  XOR2_X1 U959 ( .A(KEYINPUT111), .B(G1991), .Z(n862) );
  XNOR2_X1 U960 ( .A(G1981), .B(G1996), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n863), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U963 ( .A(G1961), .B(G1986), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U965 ( .A(G1976), .B(G1971), .Z(n867) );
  XOR2_X1 U966 ( .A(G1966), .B(n1022), .Z(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U969 ( .A(KEYINPUT110), .B(G2474), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U971 ( .A1(G124), .A2(n613), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT112), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G112), .A2(n892), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G136), .A2(n524), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G100), .A2(n899), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(G162) );
  XOR2_X1 U980 ( .A(G164), .B(G162), .Z(n880) );
  XNOR2_X1 U981 ( .A(G160), .B(n880), .ZN(n891) );
  NAND2_X1 U982 ( .A1(G118), .A2(n892), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G130), .A2(n613), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G142), .A2(n524), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G106), .A2(n899), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U988 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U991 ( .A(n891), .B(n890), .Z(n911) );
  XOR2_X1 U992 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n904) );
  NAND2_X1 U993 ( .A1(G115), .A2(n892), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G127), .A2(n613), .ZN(n893) );
  NAND2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n895), .B(KEYINPUT47), .ZN(n898) );
  NAND2_X1 U997 ( .A1(G139), .A2(n524), .ZN(n897) );
  NAND2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n902) );
  NAND2_X1 U999 ( .A1(n899), .A2(G103), .ZN(n900) );
  XOR2_X1 U1000 ( .A(KEYINPUT114), .B(n900), .Z(n901) );
  NOR2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n946) );
  XNOR2_X1 U1002 ( .A(n946), .B(KEYINPUT115), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(n905), .B(KEYINPUT46), .Z(n908) );
  XOR2_X1 U1005 ( .A(n906), .B(KEYINPUT113), .Z(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n950), .B(n909), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G395) );
  XOR2_X1 U1011 ( .A(G286), .B(n915), .Z(n917) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1013 ( .A(n918), .B(G301), .Z(n919) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n919), .ZN(G397) );
  XOR2_X1 U1015 ( .A(G2451), .B(G2430), .Z(n921) );
  XNOR2_X1 U1016 ( .A(G2438), .B(G2443), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n927) );
  XOR2_X1 U1018 ( .A(G2435), .B(G2454), .Z(n923) );
  XNOR2_X1 U1019 ( .A(G1348), .B(G1341), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n925) );
  XOR2_X1 U1021 ( .A(G2446), .B(G2427), .Z(n924) );
  XNOR2_X1 U1022 ( .A(n925), .B(n924), .ZN(n926) );
  XOR2_X1 U1023 ( .A(n927), .B(n926), .Z(n928) );
  NAND2_X1 U1024 ( .A1(G14), .A2(n928), .ZN(n935) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n935), .ZN(n932) );
  NOR2_X1 U1026 ( .A1(G227), .A2(G229), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT49), .B(n929), .Z(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(KEYINPUT117), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(G57), .ZN(G237) );
  INV_X1 U1034 ( .A(n935), .ZN(G401) );
  XOR2_X1 U1035 ( .A(G2084), .B(G160), .Z(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n944) );
  XOR2_X1 U1037 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(n940), .B(KEYINPUT51), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n958) );
  XNOR2_X1 U1042 ( .A(G164), .B(G2078), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT119), .ZN(n948) );
  XOR2_X1 U1044 ( .A(G2072), .B(n946), .Z(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(KEYINPUT50), .B(n949), .ZN(n956) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1048 ( .A(KEYINPUT118), .B(n952), .Z(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(KEYINPUT52), .B(n959), .ZN(n960) );
  INV_X1 U1053 ( .A(KEYINPUT55), .ZN(n983) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n983), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n961), .A2(G29), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT120), .B(n962), .ZN(n1013) );
  XNOR2_X1 U1057 ( .A(n963), .B(G32), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G25), .B(n964), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n975) );
  XNOR2_X1 U1060 ( .A(G2067), .B(G26), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(G28), .A2(n969), .ZN(n973) );
  XOR2_X1 U1064 ( .A(G27), .B(n970), .Z(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT121), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT53), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G2084), .B(G34), .Z(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT54), .B(n977), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G35), .B(G2090), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n983), .B(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(G29), .A2(n984), .ZN(n1011) );
  XNOR2_X1 U1076 ( .A(G1986), .B(G24), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G1976), .B(G23), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(KEYINPUT127), .B(n987), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n990), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G21), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G5), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1006) );
  XOR2_X1 U1087 ( .A(G20), .B(G1956), .Z(n999) );
  XNOR2_X1 U1088 ( .A(G1981), .B(G6), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(KEYINPUT59), .B(G1348), .Z(n1000) );
  XNOR2_X1 U1093 ( .A(G4), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1096 ( .A(KEYINPUT126), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1007), .ZN(n1008) );
  INV_X1 U1099 ( .A(G16), .ZN(n1039) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1039), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(G11), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1044) );
  NAND2_X1 U1104 ( .A1(G1971), .A2(G303), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1028) );
  XOR2_X1 U1106 ( .A(G1348), .B(n1016), .Z(n1018) );
  XOR2_X1 U1107 ( .A(G301), .B(G1961), .Z(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(KEYINPUT123), .B(n1019), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(n1022), .B(G299), .Z(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(KEYINPUT124), .B(n1029), .ZN(n1035) );
  XOR2_X1 U1116 ( .A(G168), .B(G1966), .Z(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1118 ( .A(KEYINPUT57), .B(n1032), .Z(n1033) );
  XNOR2_X1 U1119 ( .A(KEYINPUT122), .B(n1033), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1038) );
  XNOR2_X1 U1121 ( .A(G1341), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1041) );
  XNOR2_X1 U1123 ( .A(n1039), .B(KEYINPUT56), .ZN(n1040) );
  NOR2_X1 U1124 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XOR2_X1 U1125 ( .A(KEYINPUT125), .B(n1042), .Z(n1043) );
  NOR2_X1 U1126 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XOR2_X1 U1127 ( .A(n1045), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1128 ( .A(G150), .ZN(G311) );
endmodule

