//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G120gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT71), .B(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G134gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT72), .B1(new_n217), .B2(new_n212), .ZN(new_n218));
  INV_X1    g017(.A(G127gat), .ZN(new_n219));
  INV_X1    g018(.A(G134gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT72), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n216), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n213), .A2(new_n215), .B1(new_n224), .B2(new_n211), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT84), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT83), .A2(G155gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n226), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G148gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT82), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G148gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n241), .A3(G141gat), .ZN(new_n242));
  INV_X1    g041(.A(G141gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G148gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n237), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n231), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT83), .A2(G155gat), .ZN(new_n247));
  OAI21_X1  g046(.A(G162gat), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT84), .A3(KEYINPUT2), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT80), .B1(new_n235), .B2(new_n236), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n235), .B2(new_n233), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n238), .A2(G141gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n244), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n235), .A2(new_n254), .A3(new_n233), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n251), .B(new_n253), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n225), .A2(new_n250), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT4), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(KEYINPUT87), .A3(KEYINPUT4), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n225), .A2(new_n250), .A3(new_n267), .A4(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT86), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n260), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g070(.A(new_n225), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n250), .A2(new_n273), .A3(new_n260), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT85), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n271), .A2(new_n277), .A3(new_n272), .A4(new_n274), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n266), .A2(new_n269), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n264), .A2(KEYINPUT86), .A3(new_n268), .A4(new_n265), .ZN(new_n281));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n279), .A2(new_n280), .A3(new_n281), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n276), .A2(new_n278), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n261), .A2(KEYINPUT87), .A3(KEYINPUT4), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT87), .B1(new_n261), .B2(KEYINPUT4), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n269), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n286), .A2(new_n281), .A3(new_n289), .A4(new_n284), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT88), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n262), .A2(new_n268), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n282), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n272), .A2(new_n270), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n261), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n297), .B2(new_n283), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n206), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n206), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(new_n294), .B2(new_n298), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT89), .B1(new_n292), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n202), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n290), .A2(KEYINPUT88), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT88), .ZN(new_n306));
  OAI211_X1 g105(.A(KEYINPUT89), .B(new_n302), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n202), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n299), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n301), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n312), .B(new_n313), .Z(new_n314));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n317));
  OAI21_X1  g116(.A(G211gat), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G211gat), .ZN(new_n321));
  INV_X1    g120(.A(G211gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G218gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n318), .A2(new_n319), .B1(new_n324), .B2(KEYINPUT78), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT76), .B(G197gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G204gat), .ZN(new_n327));
  OR2_X1    g126(.A1(KEYINPUT76), .A2(G197gat), .ZN(new_n328));
  INV_X1    g127(.A(G204gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT76), .A2(G197gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n324), .A2(KEYINPUT78), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n325), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n325), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n315), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n332), .ZN(new_n337));
  INV_X1    g136(.A(new_n333), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n325), .A2(new_n332), .A3(new_n333), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n344), .A2(new_n345), .A3(G183gat), .A4(G190gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(G169gat), .B2(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT25), .ZN(new_n354));
  INV_X1    g153(.A(G183gat), .ZN(new_n355));
  INV_X1    g154(.A(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n344), .A2(new_n345), .B1(G183gat), .B2(G190gat), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n352), .A2(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G169gat), .ZN(new_n363));
  INV_X1    g162(.A(G176gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(new_n347), .ZN(new_n366));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(new_n348), .A3(new_n349), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT65), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(G183gat), .B2(G190gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT24), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n369), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OAI22_X1  g175(.A1(new_n362), .A2(new_n366), .B1(new_n376), .B2(KEYINPUT25), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT70), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n349), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n363), .A3(new_n364), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT69), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT69), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n374), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n379), .A2(new_n349), .ZN(new_n389));
  NOR4_X1   g188(.A1(KEYINPUT69), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n384), .B1(new_n367), .B2(new_n381), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(KEYINPUT70), .A3(new_n374), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT28), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT27), .B(G183gat), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n356), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n355), .A2(KEYINPUT27), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G183gat), .ZN(new_n399));
  AND4_X1   g198(.A1(new_n394), .A2(new_n397), .A3(new_n399), .A4(new_n356), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n388), .A2(new_n393), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n377), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n343), .B1(new_n404), .B2(KEYINPUT29), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n343), .B1(new_n377), .B2(new_n402), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n342), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n403), .A2(new_n409), .B1(G226gat), .B2(G233gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n334), .A2(new_n335), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n410), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n314), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n410), .A2(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(new_n411), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n314), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n341), .B(new_n336), .C1(new_n410), .C2(new_n406), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n413), .A2(new_n419), .A3(KEYINPUT30), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n314), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n304), .A2(new_n311), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n339), .A2(new_n409), .A3(new_n340), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n273), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(new_n270), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT90), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n274), .A2(new_n409), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n342), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n342), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n429), .A2(new_n270), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n411), .B1(new_n409), .B2(new_n274), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n427), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G22gat), .ZN(new_n440));
  INV_X1    g239(.A(G22gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G78gat), .B(G106gat), .Z(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n441), .B1(new_n435), .B2(new_n438), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n440), .A2(new_n448), .A3(new_n442), .A4(new_n446), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n403), .A2(new_n225), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n377), .A2(new_n402), .A3(new_n272), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n457), .B(KEYINPUT64), .Z(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(KEYINPUT34), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT74), .B(new_n461), .C1(new_n454), .C2(new_n455), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT73), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n377), .A2(new_n402), .A3(new_n272), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n272), .B1(new_n377), .B2(new_n402), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n455), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n457), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT34), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT33), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(G15gat), .B(G43gat), .Z(new_n476));
  XNOR2_X1  g275(.A(G71gat), .B(G99gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n472), .B(KEYINPUT32), .C1(new_n474), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT75), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n463), .A2(new_n479), .A3(new_n470), .A4(new_n481), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n482), .A3(KEYINPUT75), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n452), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT35), .B1(new_n425), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n293), .A2(new_n282), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n276), .B2(new_n278), .ZN(new_n492));
  INV_X1    g291(.A(new_n298), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n206), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n291), .B2(new_n285), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n285), .A2(new_n291), .B1(new_n294), .B2(new_n298), .ZN(new_n496));
  OAI22_X1  g295(.A1(KEYINPUT89), .A2(new_n495), .B1(new_n496), .B2(new_n206), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n497), .A2(new_n202), .B1(new_n308), .B2(new_n310), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n450), .A2(new_n451), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n498), .A2(new_n500), .A3(new_n424), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n490), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(KEYINPUT40), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n286), .A2(new_n281), .A3(new_n289), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n283), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n206), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT39), .B1(new_n297), .B2(new_n283), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n507), .B2(new_n283), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n506), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n283), .ZN(new_n514));
  INV_X1    g313(.A(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n506), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n206), .A3(new_n517), .A4(new_n509), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n300), .A2(new_n424), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n499), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n314), .B1(new_n421), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n414), .B2(new_n342), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n411), .B1(new_n410), .B2(new_n406), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT38), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n523), .A2(new_n526), .B1(new_n314), .B2(new_n421), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n421), .A2(new_n522), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n416), .A2(KEYINPUT37), .A3(new_n418), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n417), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n530), .A2(KEYINPUT94), .A3(KEYINPUT38), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT94), .B1(new_n530), .B2(KEYINPUT38), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n521), .B1(new_n498), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n486), .A2(KEYINPUT36), .A3(new_n487), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT36), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n483), .A2(new_n536), .A3(new_n485), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n425), .B2(new_n499), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(new_n539), .B2(KEYINPUT92), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n541), .B(new_n538), .C1(new_n425), .C2(new_n499), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n504), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G197gat), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT11), .B(G169gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT12), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(G1gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT16), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n550), .A2(G1gat), .ZN(new_n554));
  OAI21_X1  g353(.A(G8gat), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n552), .ZN(new_n556));
  INV_X1    g355(.A(G8gat), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n556), .B(new_n557), .C1(G1gat), .C2(new_n550), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n555), .A2(new_n558), .A3(KEYINPUT98), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT98), .B1(new_n555), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  INV_X1    g361(.A(G50gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G43gat), .ZN(new_n564));
  INV_X1    g363(.A(G43gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G50gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT15), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT96), .B(G29gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G36gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(G29gat), .A2(G36gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT14), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n568), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n564), .A2(new_n566), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT15), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n567), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(KEYINPUT97), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n569), .A2(new_n581), .A3(G36gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n562), .B(new_n574), .C1(new_n579), .C2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n573), .A2(new_n568), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(new_n578), .A3(new_n580), .A4(new_n582), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n562), .B1(new_n587), .B2(new_n574), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n561), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n574), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n555), .A2(new_n558), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n589), .A2(KEYINPUT99), .A3(new_n590), .A4(new_n593), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT100), .B(KEYINPUT18), .Z(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n589), .A2(KEYINPUT18), .A3(new_n590), .A4(new_n593), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n590), .B(KEYINPUT13), .Z(new_n601));
  INV_X1    g400(.A(new_n593), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n591), .A2(new_n592), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n549), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI211_X1 g407(.A(KEYINPUT95), .B(new_n548), .C1(new_n599), .C2(new_n605), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n543), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT8), .A2(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT103), .B1(G85gat), .B2(G92gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT7), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n623), .A2(new_n618), .A3(new_n619), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n613), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n618), .A2(new_n619), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n622), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n627), .A2(new_n612), .A3(new_n620), .A4(new_n617), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n628), .A3(KEYINPUT104), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n630), .B(new_n613), .C1(new_n621), .C2(new_n624), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n632), .A2(new_n591), .B1(KEYINPUT41), .B2(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n585), .A2(new_n588), .ZN(new_n635));
  INV_X1    g434(.A(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT105), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n639), .B1(new_n635), .B2(new_n636), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n634), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G190gat), .B(G218gat), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n642), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n647), .B(new_n634), .C1(new_n638), .C2(new_n640), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n646), .B1(new_n643), .B2(new_n648), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n229), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G57gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT101), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G57gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n661), .A3(G64gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n658), .B2(G64gat), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n662), .B(KEYINPUT102), .C1(new_n658), .C2(G64gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(G71gat), .A2(G78gat), .ZN(new_n667));
  OR2_X1    g466(.A1(G71gat), .A2(G78gat), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT9), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n665), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G57gat), .B(G64gat), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n667), .B(new_n668), .C1(new_n672), .C2(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(KEYINPUT21), .ZN(new_n676));
  NAND2_X1  g475(.A1(G231gat), .A2(G233gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(G127gat), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n592), .B1(new_n675), .B2(KEYINPUT21), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(G127gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n679), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n657), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n683), .A3(new_n656), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G230gat), .A2(G233gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n632), .A2(new_n674), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n625), .A2(new_n628), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n671), .A2(new_n692), .A3(new_n673), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT10), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT10), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n636), .A2(new_n695), .A3(new_n674), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n690), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n690), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n691), .A2(new_n698), .A3(new_n693), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(G120gat), .B(G148gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT106), .ZN(new_n702));
  XNOR2_X1  g501(.A(G176gat), .B(G204gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n697), .A2(new_n699), .A3(new_n704), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n652), .A2(new_n689), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n611), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n498), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT107), .B(G1gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1324gat));
  INV_X1    g513(.A(new_n424), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  AND3_X1   g515(.A1(new_n710), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n557), .B1(new_n710), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT42), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT42), .B2(new_n717), .ZN(G1325gat));
  INV_X1    g519(.A(G15gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n710), .A2(new_n721), .A3(new_n502), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n535), .A2(KEYINPUT108), .A3(new_n537), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(new_n535), .B2(new_n537), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n611), .A2(new_n709), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n722), .B1(new_n721), .B2(new_n726), .ZN(G1326gat));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n499), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT43), .B(G22gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n425), .A2(new_n499), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n725), .A2(new_n534), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n504), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n651), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n652), .A2(new_n731), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n731), .A2(new_n735), .B1(new_n543), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n689), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n708), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n606), .A2(new_n607), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n548), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n606), .A2(new_n607), .A3(new_n549), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n711), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n569), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n739), .A2(new_n652), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n543), .A2(new_n610), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n749), .A2(new_n498), .A3(new_n569), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n750), .A2(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(KEYINPUT45), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n747), .A2(new_n751), .A3(new_n752), .ZN(G1328gat));
  NAND2_X1  g552(.A1(new_n745), .A2(new_n715), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G36gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n749), .A2(G36gat), .A3(new_n424), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(G1329gat));
  OR2_X1    g559(.A1(new_n723), .A2(new_n724), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n737), .A2(new_n761), .A3(new_n744), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764));
  INV_X1    g563(.A(new_n749), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n565), .A3(new_n502), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n763), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(G1330gat));
  NAND2_X1  g568(.A1(new_n735), .A2(new_n731), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n543), .A2(new_n736), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n499), .A4(new_n744), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n499), .A4(new_n744), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n774), .A2(new_n775), .A3(G50gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n765), .A2(new_n563), .A3(new_n499), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT48), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(G50gat), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n777), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n776), .A2(new_n778), .B1(new_n780), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g580(.A1(new_n652), .A2(new_n689), .A3(new_n743), .A4(new_n707), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n733), .B2(new_n504), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n711), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n659), .A2(new_n661), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n784), .B(new_n785), .Z(G1332gat));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n715), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT49), .B(G64gat), .Z(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(G1333gat));
  AND2_X1   g589(.A1(new_n783), .A2(new_n502), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(G71gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n783), .A2(G71gat), .A3(new_n761), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n499), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g599(.A1(new_n689), .A2(new_n610), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n734), .A2(new_n651), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n652), .B1(new_n733), .B2(new_n504), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(KEYINPUT51), .A3(new_n801), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n708), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n615), .A3(new_n711), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n689), .A2(new_n610), .A3(new_n708), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n737), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n711), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n615), .ZN(G1336gat));
  NAND2_X1  g611(.A1(new_n804), .A2(new_n806), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n424), .A2(G92gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n707), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n770), .A2(new_n771), .A3(new_n715), .A4(new_n809), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G92gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g618(.A(G99gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n807), .A2(new_n820), .A3(new_n502), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n810), .A2(new_n761), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n820), .ZN(G1338gat));
  NOR2_X1   g622(.A1(new_n452), .A2(G106gat), .ZN(new_n824));
  AND4_X1   g623(.A1(KEYINPUT51), .A2(new_n734), .A3(new_n651), .A4(new_n801), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n805), .B2(new_n801), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n707), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n829), .A3(new_n707), .A4(new_n824), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n770), .A2(new_n771), .A3(new_n499), .A4(new_n809), .ZN(new_n831));
  XOR2_X1   g630(.A(KEYINPUT111), .B(G106gat), .Z(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  XNOR2_X1  g634(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n827), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1339gat));
  NAND3_X1  g637(.A1(new_n599), .A2(new_n605), .A3(new_n549), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n590), .B1(new_n589), .B2(new_n593), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n602), .A2(new_n603), .A3(new_n601), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n547), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n707), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n631), .A2(new_n629), .B1(new_n671), .B2(new_n673), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n671), .A2(new_n692), .A3(new_n673), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n695), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n675), .A2(KEYINPUT10), .A3(new_n632), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n698), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n697), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n698), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n704), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT55), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n706), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n844), .B1(new_n743), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n652), .ZN(new_n860));
  INV_X1    g659(.A(new_n858), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n651), .A2(new_n843), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n689), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n709), .A2(new_n610), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n865), .A2(new_n498), .A3(new_n499), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n424), .A3(new_n502), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n868), .A2(G113gat), .A3(new_n610), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n488), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n424), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n209), .B1(new_n873), .B2(new_n743), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n870), .A2(new_n874), .ZN(G1340gat));
  NAND4_X1  g674(.A1(new_n868), .A2(G120gat), .A3(new_n707), .A4(new_n869), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n207), .B1(new_n873), .B2(new_n708), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1341gat));
  NAND3_X1  g677(.A1(new_n868), .A2(new_n689), .A3(new_n869), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n214), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n738), .A2(new_n214), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n873), .B2(new_n881), .ZN(G1342gat));
  NOR2_X1   g681(.A1(new_n652), .A2(new_n715), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n220), .ZN(new_n884));
  XOR2_X1   g683(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OR3_X1    g685(.A1(new_n871), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n871), .B2(new_n884), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n868), .A2(new_n651), .A3(new_n869), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n220), .ZN(G1343gat));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n499), .C1(new_n863), .C2(new_n864), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n761), .A2(new_n498), .A3(new_n715), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n864), .ZN(new_n895));
  INV_X1    g694(.A(new_n862), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n857), .A2(new_n706), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT55), .B1(new_n854), .B2(KEYINPUT116), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n850), .A2(new_n853), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n610), .B1(new_n901), .B2(KEYINPUT117), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n903), .B(new_n897), .C1(new_n900), .C2(new_n898), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n844), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n896), .B1(new_n905), .B2(new_n652), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n895), .B1(new_n906), .B2(new_n689), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n499), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n894), .B1(KEYINPUT57), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n243), .B1(new_n909), .B2(new_n610), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n865), .A2(new_n452), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n711), .A3(new_n725), .ZN(new_n912));
  NOR4_X1   g711(.A1(new_n912), .A2(G141gat), .A3(new_n743), .A4(new_n715), .ZN(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n910), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n910), .B2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1344gat));
  AND2_X1   g717(.A1(new_n893), .A2(new_n707), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n919), .A2(new_n239), .A3(new_n241), .A4(new_n911), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT57), .B1(new_n907), .B2(new_n499), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n865), .A2(new_n891), .A3(new_n452), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n239), .A2(new_n241), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n921), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n909), .B2(new_n707), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n920), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT119), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n931), .B(new_n920), .C1(new_n925), .C2(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1345gat));
  NAND2_X1  g732(.A1(new_n230), .A2(new_n231), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n912), .A2(new_n715), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n689), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(KEYINPUT120), .A3(new_n689), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n909), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n689), .A2(new_n934), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT121), .Z(new_n943));
  NOR2_X1   g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n940), .A2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n941), .B2(new_n652), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n883), .A2(new_n227), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n912), .B2(new_n947), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n865), .A2(new_n711), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n489), .A2(new_n424), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n951), .A2(G169gat), .A3(new_n743), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n860), .A2(new_n862), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n738), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n895), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n711), .A2(new_n424), .A3(new_n501), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n452), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G169gat), .B1(new_n958), .B2(new_n743), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n953), .A2(new_n959), .ZN(G1348gat));
  OAI21_X1  g759(.A(G176gat), .B1(new_n958), .B2(new_n708), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n707), .A2(new_n364), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n951), .B2(new_n962), .ZN(G1349gat));
  OAI21_X1  g762(.A(G183gat), .B1(new_n958), .B2(new_n738), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n689), .A2(new_n395), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n951), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g766(.A(G190gat), .B1(new_n958), .B2(new_n652), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n651), .A2(new_n356), .ZN(new_n971));
  OAI22_X1  g770(.A1(new_n969), .A2(new_n970), .B1(new_n951), .B2(new_n971), .ZN(G1351gat));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n498), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n761), .A2(new_n424), .A3(new_n452), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n949), .A2(KEYINPUT123), .A3(new_n975), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(new_n610), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(G197gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n725), .A2(new_n498), .A3(new_n715), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT124), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n983), .B1(new_n922), .B2(new_n923), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n610), .A2(G197gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT125), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n981), .B(new_n988), .C1(new_n984), .C2(new_n985), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(G1352gat));
  NAND4_X1  g789(.A1(new_n949), .A2(new_n329), .A3(new_n707), .A4(new_n975), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT62), .Z(new_n992));
  OAI21_X1  g791(.A(G204gat), .B1(new_n984), .B2(new_n708), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1353gat));
  NAND4_X1  g793(.A1(new_n977), .A2(new_n978), .A3(new_n322), .A4(new_n689), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n922), .A2(new_n923), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n982), .A2(new_n738), .ZN(new_n998));
  OAI21_X1  g797(.A(G211gat), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT63), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n999), .A2(KEYINPUT63), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n996), .A2(new_n1000), .A3(new_n1001), .ZN(G1354gat));
  NOR2_X1   g801(.A1(new_n316), .A2(new_n317), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n984), .A2(new_n1003), .A3(new_n652), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n977), .A2(new_n651), .A3(new_n978), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(new_n320), .ZN(new_n1006));
  OR2_X1    g805(.A1(new_n1006), .A2(KEYINPUT127), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(KEYINPUT127), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(G1355gat));
endmodule


