//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n467), .A2(KEYINPUT67), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n467), .B2(new_n469), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n465), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(G136), .B2(new_n466), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(G162));
  NAND3_X1  g062(.A1(new_n473), .A2(G126), .A3(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n480), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n466), .A2(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n466), .A2(new_n494), .A3(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G62), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n504), .B(KEYINPUT73), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n497), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n497), .B2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT70), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n502), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n512), .A2(G543), .A3(new_n513), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n507), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n506), .B1(new_n518), .B2(new_n519), .ZN(G166));
  NAND4_X1  g095(.A1(new_n512), .A2(new_n502), .A3(G89), .A4(new_n513), .ZN(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n502), .A2(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n512), .A2(G51), .A3(G543), .A4(new_n513), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n521), .A2(new_n527), .A3(new_n528), .ZN(G168));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n500), .B2(new_n501), .ZN(new_n531));
  AND2_X1   g106(.A1(G77), .A2(G543), .ZN(new_n532));
  OAI21_X1  g107(.A(G651), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n512), .A2(G52), .A3(G543), .A4(new_n513), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n512), .A2(new_n502), .A3(G90), .A4(new_n513), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G171));
  NAND4_X1  g111(.A1(new_n512), .A2(new_n502), .A3(G81), .A4(new_n513), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n512), .A2(G43), .A3(G543), .A4(new_n513), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n500), .B2(new_n501), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  AND3_X1   g120(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g123(.A(KEYINPUT74), .B(new_n543), .C1(new_n548), .C2(new_n541), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n549), .A3(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n539), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(new_n514), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n548), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n558), .A2(G91), .B1(new_n561), .B2(G651), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n512), .A2(G53), .A3(G543), .A4(new_n513), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n509), .A2(new_n511), .B1(KEYINPUT6), .B2(new_n497), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n565), .A2(new_n566), .A3(G53), .A4(G543), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n564), .A2(KEYINPUT75), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT75), .B1(new_n564), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n562), .B1(new_n568), .B2(new_n569), .ZN(G299));
  NAND3_X1  g145(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G301));
  NAND3_X1  g146(.A1(new_n521), .A2(new_n527), .A3(new_n528), .ZN(G286));
  XNOR2_X1  g147(.A(new_n517), .B(KEYINPUT72), .ZN(new_n573));
  INV_X1    g148(.A(new_n506), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G303));
  NAND3_X1  g150(.A1(new_n565), .A2(G87), .A3(new_n502), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n515), .ZN(G288));
  NAND4_X1  g154(.A1(new_n512), .A2(G48), .A3(G543), .A4(new_n513), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n497), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n558), .A2(G86), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n548), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n514), .B1(new_n515), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n594), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n512), .A2(new_n502), .A3(G92), .A4(new_n513), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n601), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n565), .A2(G92), .A3(new_n603), .A4(new_n502), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n500), .B2(new_n501), .ZN(new_n606));
  AND2_X1   g181(.A1(G79), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n565), .A2(G54), .A3(G543), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n602), .A2(new_n604), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n599), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n599), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  OAI21_X1  g194(.A(G868), .B1(new_n610), .B2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n473), .A2(new_n468), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT79), .B(G2100), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n466), .A2(G135), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT80), .Z(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G2105), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n481), .B2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n627), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT82), .Z(G156));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n642), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(G14), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(G2072), .A2(G2078), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n442), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2084), .B(G2090), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n655), .A2(new_n659), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n658), .A2(KEYINPUT83), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(KEYINPUT83), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n666), .A3(new_n656), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n667), .B(new_n659), .C1(new_n662), .C2(new_n656), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n684), .C1(new_n675), .C2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n686), .ZN(new_n691));
  INV_X1    g266(.A(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g268(.A1(new_n689), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n689), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  OR2_X1    g271(.A1(G6), .A2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(G305), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT32), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G1981), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G288), .B2(new_n698), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT33), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G1976), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(G1976), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n703), .A2(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n698), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n698), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1971), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(KEYINPUT89), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(KEYINPUT89), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n711), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n711), .A2(new_n719), .A3(new_n715), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n698), .A2(G24), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT87), .Z(new_n722));
  INV_X1    g297(.A(new_n597), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n723), .A2(new_n595), .B1(G651), .B2(new_n589), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n722), .B1(new_n724), .B2(new_n698), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1986), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT86), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n466), .A2(G131), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n481), .A2(G119), .ZN(new_n731));
  OR2_X1    g306(.A1(G95), .A2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G107), .C2(new_n480), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n726), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n720), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT36), .B1(new_n718), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n741), .A2(new_n742), .A3(new_n720), .A4(new_n738), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n473), .A2(G127), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n480), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n466), .A2(G139), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT25), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n747), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT91), .ZN(new_n753));
  MUX2_X1   g328(.A(G33), .B(new_n753), .S(G29), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G2072), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT92), .ZN(new_n756));
  NOR2_X1   g331(.A1(G27), .A2(G29), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G164), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n698), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n698), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1961), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n754), .B2(G2072), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n756), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G34), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(new_n727), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G160), .B2(new_n727), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G29), .A2(G35), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G162), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT29), .B(G2090), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n698), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n698), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G1966), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n774), .A2(new_n775), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n778), .A2(G1966), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n776), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n611), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G4), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT90), .B(G1348), .Z(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n698), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n552), .B2(new_n698), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n787), .C1(G1341), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(G28), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n727), .B1(new_n792), .B2(G28), .ZN(new_n794));
  OAI221_X1 g369(.A(new_n791), .B1(new_n793), .B2(new_n794), .C1(new_n634), .C2(new_n727), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n727), .A2(G32), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n481), .A2(G129), .ZN(new_n797));
  NAND3_X1  g372(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT26), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(KEYINPUT26), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n468), .A2(G105), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  AOI211_X1 g378(.A(new_n801), .B(new_n803), .C1(G141), .C2(new_n466), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n796), .B1(new_n804), .B2(new_n727), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT27), .B(G1996), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n795), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n805), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n789), .A2(G1341), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n727), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n466), .A2(G140), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n481), .A2(G128), .ZN(new_n814));
  OR2_X1    g389(.A1(G104), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(new_n727), .ZN(new_n819));
  INV_X1    g394(.A(G2067), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n782), .A2(new_n790), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n698), .A2(G20), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT23), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n615), .B2(new_n698), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1956), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n766), .A2(new_n772), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT96), .B1(new_n744), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n832), .B(new_n829), .C1(new_n740), .C2(new_n743), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(G311));
  NAND2_X1  g409(.A1(new_n744), .A2(new_n830), .ZN(G150));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n618), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n512), .A2(new_n502), .A3(G93), .A4(new_n513), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n512), .A2(G55), .A3(G543), .A4(new_n513), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n500), .B2(new_n501), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n841), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(G67), .B1(new_n546), .B2(new_n547), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n847), .A2(KEYINPUT97), .A3(new_n844), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(G651), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n840), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n551), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n550), .A2(new_n539), .A3(new_n840), .A4(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n837), .B(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n855), .A2(new_n856), .A3(G860), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n850), .A2(G860), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  INV_X1    g435(.A(new_n634), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n478), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G164), .B(new_n818), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n753), .B(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n804), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n804), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n466), .A2(G142), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n481), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n480), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n624), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n734), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT98), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n876), .A2(KEYINPUT98), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n869), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n869), .A2(KEYINPUT99), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n876), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n869), .A2(KEYINPUT99), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n864), .B(new_n879), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n877), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n867), .A3(new_n868), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n886), .B2(new_n863), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g464(.A1(new_n850), .A2(G868), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n724), .A2(G303), .ZN(new_n891));
  NAND2_X1  g466(.A1(G290), .A2(G166), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G288), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT100), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n896));
  NAND2_X1  g471(.A1(G288), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G305), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(G305), .A2(new_n895), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n893), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n891), .A2(new_n892), .A3(new_n901), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT42), .Z(new_n906));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n907));
  NAND2_X1  g482(.A1(G299), .A2(new_n610), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n611), .B(new_n562), .C1(new_n569), .C2(new_n568), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n610), .A2(G559), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n853), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n908), .A2(new_n909), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n916), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n906), .B1(new_n907), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n907), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n920), .B(new_n921), .Z(new_n922));
  AOI21_X1  g497(.A(new_n890), .B1(new_n922), .B2(G868), .ZN(G295));
  AOI21_X1  g498(.A(new_n890), .B1(new_n922), .B2(G868), .ZN(G331));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND2_X1  g500(.A1(G171), .A2(G168), .ZN(new_n926));
  NAND2_X1  g501(.A1(G301), .A2(G286), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n853), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n918), .A2(new_n930), .ZN(new_n931));
  AND4_X1   g506(.A1(new_n550), .A2(new_n539), .A3(new_n840), .A4(new_n849), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n550), .A2(new_n539), .B1(new_n840), .B2(new_n849), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n853), .A2(new_n938), .A3(new_n928), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n929), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT103), .B1(new_n914), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT41), .B1(new_n908), .B2(new_n909), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n853), .A2(new_n938), .A3(new_n928), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n938), .B1(new_n853), .B2(new_n928), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n930), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n936), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n905), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n925), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n936), .B(new_n905), .C1(new_n941), .C2(new_n949), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n936), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n914), .A2(new_n940), .A3(KEYINPUT103), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n948), .B1(new_n944), .B2(new_n947), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n951), .B(new_n955), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n935), .A2(new_n929), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n945), .A2(new_n946), .ZN(new_n961));
  OAI22_X1  g536(.A1(new_n914), .A2(new_n960), .B1(new_n931), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n905), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n958), .A2(new_n963), .A3(KEYINPUT104), .A4(new_n959), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n954), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n971), .B2(new_n905), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT43), .B1(new_n972), .B2(new_n958), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n958), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT44), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT105), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n970), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(G397));
  NOR2_X1   g555(.A1(G164), .A2(G1384), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT107), .B(G40), .Z(new_n986));
  OAI211_X1 g561(.A(new_n476), .B(new_n986), .C1(new_n470), .C2(new_n471), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1986), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n724), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n991), .B2(KEYINPUT108), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(KEYINPUT108), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n724), .A2(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n804), .B(G1996), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n817), .B(new_n820), .ZN(new_n997));
  INV_X1    g572(.A(new_n734), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n736), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n998), .A2(new_n736), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n996), .A2(new_n997), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n992), .A2(new_n995), .B1(new_n988), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT109), .B1(new_n981), .B2(new_n983), .ZN(new_n1003));
  INV_X1    g578(.A(new_n987), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1005), .B(new_n982), .C1(G164), .C2(G1384), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n493), .A2(new_n495), .ZN(new_n1009));
  INV_X1    g584(.A(new_n491), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n981), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1971), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1019), .A3(new_n1012), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1004), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G2090), .ZN(new_n1023));
  OAI21_X1  g598(.A(G8), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(G166), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n987), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1020), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1022), .A2(KEYINPUT116), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1032), .B1(new_n1039), .B2(new_n1018), .ZN(new_n1040));
  INV_X1    g615(.A(G1971), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1017), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1003), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT117), .A3(new_n1038), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(G8), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1031), .B1(new_n1047), .B2(new_n1030), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n1013), .B2(new_n987), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(G288), .B2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n576), .A2(new_n577), .ZN(new_n1054));
  INV_X1    g629(.A(new_n515), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G49), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1054), .A2(new_n1056), .A3(KEYINPUT111), .A4(G1976), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT112), .B(KEYINPUT52), .C1(new_n1050), .C2(new_n1058), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1059), .B(new_n1060), .C1(G1976), .C2(new_n894), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n584), .A2(new_n585), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n580), .B(KEYINPUT76), .ZN(new_n1066));
  OAI21_X1  g641(.A(G1981), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n582), .A2(new_n702), .A3(new_n584), .A4(new_n585), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1050), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(KEYINPUT49), .A3(new_n1068), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT113), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT113), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1063), .B(new_n1064), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1050), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1072), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1073), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(KEYINPUT118), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n981), .A2(new_n983), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n1004), .C1(KEYINPUT45), .C2(new_n981), .ZN(new_n1088));
  INV_X1    g663(.A(G1966), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1033), .A2(new_n771), .A3(new_n1020), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1027), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1092), .A2(G168), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1048), .A2(new_n1086), .A3(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1092), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1023), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1027), .B1(new_n1045), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1029), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1076), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT120), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1100), .A2(new_n1101), .A3(new_n1105), .A4(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1096), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1101), .A2(new_n1031), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n894), .A2(new_n1052), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1083), .B2(new_n1073), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1068), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1050), .B(KEYINPUT114), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1112), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1109), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1048), .A2(new_n1086), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1090), .A2(new_n1091), .A3(G168), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  AND2_X1   g696(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  NOR2_X1   g699(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1120), .A2(G8), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1092), .A2(G286), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1123), .A2(new_n1124), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n760), .A2(KEYINPUT53), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1088), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1022), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(G1961), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1017), .A2(new_n760), .A3(new_n1003), .A4(new_n1043), .ZN(new_n1135));
  AOI211_X1 g710(.A(new_n1131), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(G301), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1129), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1121), .A2(new_n1122), .B1(G286), .B2(new_n1092), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1124), .B1(new_n1139), .B2(new_n1127), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1118), .B1(new_n1119), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1108), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1133), .B1(new_n1135), .B2(new_n1134), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n760), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1017), .A2(new_n477), .A3(new_n985), .A4(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(G301), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1136), .B2(G301), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1148), .A2(new_n1149), .B1(new_n1127), .B2(new_n1139), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1151), .B2(G171), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT124), .B1(new_n1136), .B2(G301), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1131), .ZN(new_n1154));
  AND4_X1   g729(.A1(KEYINPUT124), .A2(new_n1144), .A3(G301), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1152), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1150), .A2(new_n1156), .A3(new_n1086), .A4(new_n1048), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT56), .B(G2072), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1017), .A2(new_n1003), .A3(new_n1043), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n564), .A2(new_n567), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n562), .A2(new_n1160), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n615), .A2(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G1956), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1022), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1159), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1159), .A2(new_n1165), .A3(KEYINPUT121), .A4(new_n1167), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1164), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT61), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(KEYINPUT61), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1168), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT59), .ZN(new_n1178));
  INV_X1    g753(.A(G1996), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1017), .A2(new_n1179), .A3(new_n1003), .A4(new_n1043), .ZN(new_n1180));
  XOR2_X1   g755(.A(KEYINPUT58), .B(G1341), .Z(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n1013), .B2(new_n987), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1178), .B1(new_n1183), .B2(new_n552), .ZN(new_n1184));
  AOI211_X1 g759(.A(KEYINPUT59), .B(new_n551), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1176), .A2(new_n1177), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT122), .B1(new_n1175), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1183), .A2(new_n552), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1183), .A2(new_n1178), .A3(new_n552), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1173), .B2(new_n1164), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1189), .A2(new_n1190), .B1(new_n1192), .B2(new_n1168), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n1194));
  AOI22_X1  g769(.A1(new_n1170), .A2(new_n1171), .B1(new_n1164), .B2(new_n1173), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1193), .B(new_n1194), .C1(KEYINPUT61), .C2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(G1348), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1013), .A2(new_n987), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1022), .A2(new_n1197), .B1(new_n1198), .B2(new_n820), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT60), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(new_n611), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(KEYINPUT60), .B2(new_n1199), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1187), .A2(new_n1196), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1174), .B1(new_n610), .B2(new_n1199), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1172), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1157), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1002), .B1(new_n1143), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n989), .A2(new_n994), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1208), .A2(KEYINPUT48), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1208), .A2(KEYINPUT48), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n1209), .B(new_n1210), .C1(new_n988), .C2(new_n1001), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n988), .A2(new_n1179), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT46), .Z(new_n1213));
  NAND2_X1  g788(.A1(new_n804), .A2(new_n997), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT125), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT47), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n996), .A2(new_n997), .ZN(new_n1219));
  OAI22_X1  g794(.A1(new_n1219), .A2(new_n999), .B1(G2067), .B2(new_n817), .ZN(new_n1220));
  AOI211_X1 g795(.A(new_n1211), .B(new_n1218), .C1(new_n988), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1207), .A2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g797(.A1(G227), .A2(new_n460), .ZN(new_n1224));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n1225));
  XNOR2_X1  g799(.A(new_n1224), .B(new_n1225), .ZN(new_n1226));
  OAI211_X1 g800(.A(new_n1226), .B(new_n653), .C1(new_n694), .C2(new_n695), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n883), .B2(new_n887), .ZN(new_n1228));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1229));
  AND3_X1   g803(.A1(new_n1228), .A2(new_n1229), .A3(new_n968), .ZN(new_n1230));
  AOI21_X1  g804(.A(new_n1229), .B1(new_n1228), .B2(new_n968), .ZN(new_n1231));
  NOR2_X1   g805(.A1(new_n1230), .A2(new_n1231), .ZN(G308));
  NAND2_X1  g806(.A1(new_n1228), .A2(new_n968), .ZN(G225));
endmodule


