//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921;
  NOR3_X1   g000(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n210), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n207), .B(KEYINPUT90), .ZN(new_n216));
  INV_X1    g015(.A(new_n205), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(new_n202), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n211), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT91), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n215), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n212), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(G1gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G1gat), .B2(new_n226), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n229), .B(G8gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n225), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n224), .A2(new_n230), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G197gat), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT11), .B(G169gat), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT12), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n224), .B(new_n230), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n233), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n232), .A2(KEYINPUT18), .A3(new_n233), .A4(new_n234), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n237), .A2(new_n243), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n235), .A2(new_n236), .B1(new_n244), .B2(new_n245), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(KEYINPUT92), .A3(new_n243), .A4(new_n247), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n247), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n250), .A2(new_n252), .B1(new_n253), .B2(new_n242), .ZN(new_n254));
  XOR2_X1   g053(.A(G141gat), .B(G148gat), .Z(new_n255));
  INV_X1    g054(.A(G155gat), .ZN(new_n256));
  INV_X1    g055(.A(G162gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT2), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(KEYINPUT77), .A3(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G155gat), .B(G162gat), .Z(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(KEYINPUT77), .A3(new_n258), .A4(new_n255), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT22), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT75), .B(G218gat), .Z(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G197gat), .B(G204gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT29), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT3), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n264), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(G228gat), .A2(G233gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n273), .A2(new_n274), .ZN(new_n282));
  INV_X1    g081(.A(new_n264), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n278), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT78), .B1(new_n264), .B2(KEYINPUT3), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT29), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n280), .B(new_n281), .C1(new_n282), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n264), .B1(new_n275), .B2(KEYINPUT3), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n287), .B2(new_n282), .ZN(new_n290));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT82), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n290), .A2(KEYINPUT83), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT83), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G22gat), .ZN(new_n296));
  INV_X1    g095(.A(G22gat), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n288), .B(new_n297), .C1(new_n293), .C2(new_n294), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n300), .B1(new_n295), .B2(G22gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G78gat), .B(G106gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT31), .B(G50gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n299), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n296), .A2(new_n300), .A3(new_n298), .A4(new_n304), .ZN(new_n307));
  XOR2_X1   g106(.A(G15gat), .B(G43gat), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT70), .ZN(new_n309));
  XNOR2_X1  g108(.A(G71gat), .B(G99gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G227gat), .A2(G233gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(KEYINPUT1), .ZN(new_n315));
  XOR2_X1   g114(.A(G127gat), .B(G134gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n325), .A2(KEYINPUT67), .B1(new_n323), .B2(new_n320), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n319), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT65), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n332), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n331), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT27), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(G190gat), .B1(new_n344), .B2(new_n338), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n341), .A2(KEYINPUT66), .B1(new_n345), .B2(KEYINPUT28), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n347), .B(new_n331), .C1(new_n335), .C2(new_n340), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n328), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT68), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(new_n328), .C1(new_n346), .C2(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n322), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n318), .A2(KEYINPUT24), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT64), .B(G183gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G190gat), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n359), .A2(new_n361), .B1(new_n337), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n357), .B1(new_n356), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n317), .B1(new_n353), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n317), .ZN(new_n371));
  INV_X1    g170(.A(new_n369), .ZN(new_n372));
  AOI211_X1 g171(.A(new_n371), .B(new_n372), .C1(new_n350), .C2(new_n352), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n313), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n311), .B1(new_n374), .B2(KEYINPUT32), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n376));
  INV_X1    g175(.A(new_n352), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT65), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n339), .B1(new_n338), .B2(new_n332), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n330), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n347), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n341), .A2(KEYINPUT66), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n334), .B1(new_n363), .B2(KEYINPUT27), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n329), .B1(new_n383), .B2(G190gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n351), .B1(new_n385), .B2(new_n328), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n369), .B1(new_n377), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n371), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n353), .A2(new_n317), .A3(new_n369), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n312), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n376), .B1(new_n390), .B2(KEYINPUT33), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n374), .A2(KEYINPUT69), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n312), .A3(new_n389), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT34), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT34), .B1(new_n395), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n374), .B(KEYINPUT32), .C1(new_n392), .C2(new_n311), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n394), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n306), .A2(new_n307), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n400), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT71), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(KEYINPUT71), .A3(new_n400), .ZN(new_n406));
  INV_X1    g205(.A(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n283), .A2(new_n410), .A3(new_n317), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n283), .A2(new_n317), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT4), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n412), .A3(KEYINPUT4), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n285), .A2(new_n286), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n317), .B1(new_n264), .B2(KEYINPUT3), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n416), .A2(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n419), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n415), .A2(new_n411), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n371), .A2(new_n264), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n414), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(new_n422), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n420), .A2(new_n423), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G1gat), .B(G29gat), .Z(new_n432));
  XNOR2_X1  g231(.A(G57gat), .B(G85gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT6), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT6), .B1(new_n431), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n438), .B2(KEYINPUT81), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n438), .A2(KEYINPUT81), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n349), .A2(new_n369), .ZN(new_n444));
  AND2_X1   g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n282), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n372), .B1(new_n350), .B2(new_n352), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n445), .A2(KEYINPUT29), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n451), .A2(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n349), .A2(new_n369), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n448), .A2(new_n445), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n451), .B(KEYINPUT76), .C1(new_n454), .C2(new_n447), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n452), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(KEYINPUT30), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(new_n464), .A3(new_n459), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n443), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT35), .B1(new_n409), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n401), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n399), .B1(new_n400), .B2(new_n394), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n403), .A2(KEYINPUT74), .A3(new_n407), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n306), .A2(new_n307), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n420), .A2(new_n423), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n426), .A2(new_n430), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n436), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n440), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT35), .B1(new_n481), .B2(new_n439), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n466), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n468), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(new_n443), .A3(new_n466), .ZN(new_n485));
  INV_X1    g284(.A(new_n420), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n422), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n414), .A2(new_n421), .A3(new_n428), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT39), .B(new_n489), .C1(new_n420), .C2(new_n421), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(new_n437), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n438), .B1(new_n491), .B2(new_n492), .ZN(new_n494));
  AND4_X1   g293(.A1(new_n465), .A2(new_n463), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT37), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT87), .A3(new_n461), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT37), .B1(new_n452), .B2(new_n455), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT86), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n500), .B(KEYINPUT37), .C1(new_n452), .C2(new_n455), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT87), .B1(new_n496), .B2(new_n461), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT38), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n481), .A2(new_n460), .A3(new_n439), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n498), .B(KEYINPUT86), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n454), .A2(new_n282), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n387), .A2(new_n449), .B1(new_n445), .B2(new_n444), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n282), .ZN(new_n510));
  AOI211_X1 g309(.A(KEYINPUT38), .B(new_n459), .C1(new_n507), .C2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n505), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n495), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n485), .B1(new_n513), .B2(new_n476), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n401), .A2(KEYINPUT36), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n408), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n403), .A2(new_n407), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(new_n469), .A3(new_n401), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n473), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT73), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n408), .A2(new_n522), .A3(new_n515), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n254), .B1(new_n484), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT103), .ZN(new_n527));
  XNOR2_X1  g326(.A(G183gat), .B(G211gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT97), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(new_n256), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n529), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G127gat), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT94), .B(G57gat), .Z(new_n535));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536));
  NAND2_X1  g335(.A1(G71gat), .A2(G78gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n535), .A2(G64gat), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G64gat), .B2(new_n535), .ZN(new_n539));
  OR2_X1    g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(KEYINPUT93), .B2(new_n537), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(KEYINPUT93), .B2(new_n537), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n537), .B1(new_n540), .B2(new_n536), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G57gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G64gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n539), .A2(new_n542), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT21), .ZN(new_n550));
  INV_X1    g349(.A(G231gat), .ZN(new_n551));
  INV_X1    g350(.A(G233gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(G231gat), .B(G233gat), .C1(new_n549), .C2(KEYINPUT21), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n534), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n230), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n549), .B2(KEYINPUT21), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(new_n534), .A3(new_n554), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n556), .B2(new_n560), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n533), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n561), .A3(new_n532), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT8), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n570), .B(new_n572), .C1(G85gat), .C2(G92gat), .ZN(new_n573));
  XOR2_X1   g372(.A(G99gat), .B(G106gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n568), .B1(new_n224), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT98), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n225), .A2(new_n231), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n580), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n577), .A2(new_n585), .A3(new_n578), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n581), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n581), .B2(new_n586), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n567), .A2(new_n589), .A3(KEYINPUT99), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT99), .B1(new_n567), .B2(new_n589), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT102), .Z(new_n595));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n575), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n549), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT100), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n549), .A2(new_n602), .A3(new_n599), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n575), .A2(new_n547), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n549), .B2(new_n575), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n597), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n597), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n595), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n601), .B(new_n603), .C1(KEYINPUT10), .C2(new_n606), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n612), .B2(new_n596), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n614), .A3(new_n594), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n614), .B1(new_n613), .B2(new_n594), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n590), .A2(new_n591), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n526), .A2(new_n527), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n527), .B1(new_n526), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n443), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G1gat), .ZN(G1324gat));
  INV_X1    g427(.A(new_n466), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT16), .B(G8gat), .Z(new_n630));
  OAI211_X1 g429(.A(new_n629), .B(new_n630), .C1(new_n622), .C2(new_n623), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT42), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT105), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n629), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n636));
  AOI22_X1  g435(.A1(new_n635), .A2(G8gat), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(G1325gat));
  OR3_X1    g437(.A1(new_n624), .A2(G15gat), .A3(new_n475), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n521), .A2(new_n523), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n522), .B1(new_n408), .B2(new_n515), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT106), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n517), .A2(new_n643), .A3(new_n521), .A4(new_n523), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(G15gat), .B1(new_n624), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n639), .A2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n624), .A2(new_n477), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  AND4_X1   g450(.A1(new_n526), .A2(new_n567), .A3(new_n589), .A4(new_n619), .ZN(new_n652));
  INV_X1    g451(.A(G29gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n653), .A3(new_n626), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT45), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n484), .A2(new_n525), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(KEYINPUT44), .A3(new_n589), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n250), .A2(new_n252), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n253), .A2(new_n242), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n254), .A2(KEYINPUT107), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n567), .A2(new_n619), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n589), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n642), .A2(new_n514), .A3(new_n644), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(new_n484), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n657), .B(new_n666), .C1(new_n669), .C2(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n443), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n671), .ZN(G1328gat));
  INV_X1    g471(.A(G36gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n652), .A2(new_n673), .A3(new_n629), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT46), .Z(new_n675));
  OAI21_X1  g474(.A(G36gat), .B1(new_n670), .B2(new_n466), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1329gat));
  OAI21_X1  g476(.A(G43gat), .B1(new_n670), .B2(new_n646), .ZN(new_n678));
  INV_X1    g477(.A(G43gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n475), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n652), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684));
  OAI21_X1  g483(.A(G50gat), .B1(new_n670), .B2(new_n477), .ZN(new_n685));
  INV_X1    g484(.A(G50gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n652), .A2(new_n686), .A3(new_n476), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(KEYINPUT108), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n685), .A2(new_n684), .A3(new_n687), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n689), .A2(KEYINPUT48), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(KEYINPUT48), .ZN(new_n693));
  INV_X1    g492(.A(new_n691), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n688), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(G1331gat));
  NAND2_X1  g495(.A1(new_n668), .A2(new_n484), .ZN(new_n697));
  AND4_X1   g496(.A1(new_n591), .A2(new_n664), .A3(new_n590), .A4(new_n618), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n443), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT110), .B(G57gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1332gat));
  XNOR2_X1  g501(.A(new_n466), .B(KEYINPUT111), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  AND2_X1   g505(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n705), .B2(new_n706), .ZN(G1333gat));
  OR3_X1    g508(.A1(new_n699), .A2(G71gat), .A3(new_n475), .ZN(new_n710));
  OAI21_X1  g509(.A(G71gat), .B1(new_n699), .B2(new_n646), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g512(.A1(new_n699), .A2(new_n477), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(G78gat), .Z(G1335gat));
  INV_X1    g514(.A(new_n664), .ZN(new_n716));
  INV_X1    g515(.A(new_n567), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n618), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n657), .B(new_n720), .C1(KEYINPUT44), .C2(new_n669), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n443), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n669), .A2(KEYINPUT51), .A3(new_n718), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT51), .B1(new_n669), .B2(new_n718), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n619), .A2(G85gat), .A3(new_n443), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT112), .Z(new_n728));
  OAI21_X1  g527(.A(new_n722), .B1(new_n726), .B2(new_n728), .ZN(G1336gat));
  OAI21_X1  g528(.A(G92gat), .B1(new_n721), .B2(new_n466), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n697), .A2(new_n589), .A3(new_n718), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n723), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n725), .A2(KEYINPUT113), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n704), .A2(new_n619), .A3(G92gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n730), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT52), .ZN(new_n740));
  OAI21_X1  g539(.A(G92gat), .B1(new_n721), .B2(new_n704), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n741), .B(new_n742), .C1(new_n726), .C2(new_n738), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1337gat));
  OAI21_X1  g543(.A(G99gat), .B1(new_n721), .B2(new_n646), .ZN(new_n745));
  OR3_X1    g544(.A1(new_n475), .A2(new_n619), .A3(G99gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n726), .B2(new_n746), .ZN(G1338gat));
  NOR3_X1   g546(.A1(new_n477), .A2(new_n619), .A3(G106gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n735), .A2(new_n736), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G106gat), .B1(new_n721), .B2(new_n477), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT53), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n748), .B1(new_n724), .B2(new_n725), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n755), .B1(new_n749), .B2(new_n750), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT114), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n594), .B1(new_n608), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n604), .A2(new_n597), .A3(new_n607), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n612), .A2(new_n596), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT54), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n617), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n615), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n763), .A2(KEYINPUT55), .A3(new_n766), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n662), .A2(new_n774), .A3(new_n663), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n232), .A2(new_n234), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(G229gat), .A3(G233gat), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n244), .B2(new_n245), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n241), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n782), .A2(new_n658), .A3(new_n618), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n589), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n782), .A2(new_n658), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n774), .A3(new_n589), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n567), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n621), .A2(new_n664), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n476), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n703), .A2(new_n475), .A3(new_n443), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G113gat), .B1(new_n793), .B2(new_n254), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n443), .B1(new_n789), .B2(new_n790), .ZN(new_n795));
  INV_X1    g594(.A(new_n409), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n796), .A3(new_n704), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n664), .A2(G113gat), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(KEYINPUT116), .Z(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n797), .B2(new_n799), .ZN(G1340gat));
  OAI21_X1  g599(.A(G120gat), .B1(new_n793), .B2(new_n619), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n619), .A2(G120gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT117), .ZN(G1341gat));
  OAI21_X1  g603(.A(G127gat), .B1(new_n793), .B2(new_n567), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n717), .A2(new_n534), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT118), .Z(G1342gat));
  NAND2_X1  g607(.A1(new_n795), .A2(new_n796), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n589), .A2(new_n466), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT119), .Z(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(G134gat), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n809), .A2(KEYINPUT56), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G134gat), .B1(new_n793), .B2(new_n667), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT56), .B1(new_n809), .B2(new_n813), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT120), .ZN(G1343gat));
  AND3_X1   g617(.A1(new_n795), .A2(new_n476), .A3(new_n646), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n704), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n254), .A2(G141gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n645), .A2(new_n443), .A3(new_n703), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n789), .A2(new_n790), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n476), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n476), .A2(KEYINPUT57), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n773), .A2(new_n254), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n667), .B1(new_n831), .B2(new_n783), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n717), .B1(new_n832), .B2(new_n787), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n833), .A2(new_n834), .B1(new_n621), .B2(new_n664), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n830), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n825), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n254), .ZN(new_n839));
  INV_X1    g638(.A(G141gat), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n716), .B(new_n825), .C1(new_n829), .C2(new_n837), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n820), .A2(new_n821), .B1(new_n842), .B2(G141gat), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n824), .A2(new_n841), .B1(new_n843), .B2(new_n823), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n620), .A2(new_n660), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(new_n833), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n846), .B2(new_n476), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n477), .B(new_n826), .C1(new_n789), .C2(new_n790), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n618), .B(new_n825), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G148gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT59), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n618), .B(new_n825), .C1(new_n829), .C2(new_n837), .ZN(new_n852));
  INV_X1    g651(.A(G148gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(KEYINPUT59), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n852), .A2(KEYINPUT123), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT123), .B1(new_n852), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n820), .A2(new_n853), .A3(new_n618), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1345gat));
  NAND3_X1  g658(.A1(new_n820), .A2(new_n256), .A3(new_n717), .ZN(new_n860));
  OAI21_X1  g659(.A(G155gat), .B1(new_n838), .B2(new_n567), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1346gat));
  OAI21_X1  g661(.A(G162gat), .B1(new_n838), .B2(new_n667), .ZN(new_n863));
  INV_X1    g662(.A(new_n811), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n819), .A2(new_n257), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1347gat));
  NOR3_X1   g665(.A1(new_n475), .A2(new_n626), .A3(new_n466), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n791), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(G169gat), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n254), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n626), .B1(new_n789), .B2(new_n790), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n704), .A2(new_n409), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n716), .A3(new_n872), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n868), .A2(new_n870), .B1(new_n873), .B2(new_n869), .ZN(G1348gat));
  INV_X1    g673(.A(G176gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n868), .B2(new_n618), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n871), .A2(new_n872), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(G176gat), .A3(new_n619), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n876), .A2(new_n878), .ZN(G1349gat));
  OAI21_X1  g678(.A(new_n717), .B1(new_n379), .B2(new_n378), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n868), .A2(new_n717), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n363), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT60), .Z(G1350gat));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n589), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n887));
  AND4_X1   g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(G190gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n366), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n886), .A2(new_n889), .B1(new_n885), .B2(new_n887), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n589), .A2(new_n366), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n888), .A2(new_n890), .B1(new_n877), .B2(new_n891), .ZN(G1351gat));
  INV_X1    g691(.A(G197gat), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n645), .A2(new_n626), .A3(new_n466), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n660), .B(new_n894), .C1(new_n847), .C2(new_n848), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(KEYINPUT126), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(KEYINPUT126), .B2(new_n895), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n645), .A2(new_n477), .A3(new_n704), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n871), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n893), .A3(new_n716), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n897), .A2(new_n904), .ZN(G1352gat));
  XOR2_X1   g704(.A(KEYINPUT127), .B(G204gat), .Z(new_n906));
  OR3_X1    g705(.A1(new_n902), .A2(new_n619), .A3(new_n906), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT62), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(KEYINPUT62), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n847), .A2(new_n848), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n618), .A3(new_n894), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n906), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(G1353gat));
  NAND3_X1  g712(.A1(new_n903), .A2(new_n267), .A3(new_n717), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n717), .A3(new_n894), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n915), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT63), .B1(new_n915), .B2(G211gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1354gat));
  AOI21_X1  g717(.A(G218gat), .B1(new_n903), .B2(new_n589), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n910), .A2(new_n894), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n667), .A2(new_n266), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1355gat));
endmodule


