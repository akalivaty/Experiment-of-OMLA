

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U556 ( .A1(G8), .A2(n680), .ZN(n724) );
  INV_X2 U557 ( .A(n662), .ZN(n680) );
  AND2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n600) );
  XNOR2_X1 U559 ( .A(n521), .B(G543), .ZN(n526) );
  BUF_X1 U560 ( .A(n600), .Z(n891) );
  INV_X1 U561 ( .A(KEYINPUT17), .ZN(n539) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n540) );
  INV_X1 U563 ( .A(KEYINPUT28), .ZN(n620) );
  AND2_X1 U564 ( .A1(n541), .A2(G2105), .ZN(n598) );
  XNOR2_X1 U565 ( .A(n628), .B(KEYINPUT13), .ZN(n629) );
  INV_X1 U566 ( .A(KEYINPUT91), .ZN(n601) );
  NAND2_X1 U567 ( .A1(G114), .A2(n600), .ZN(n602) );
  NOR2_X1 U568 ( .A1(G651), .A2(n526), .ZN(n522) );
  NOR2_X2 U569 ( .A1(n545), .A2(n544), .ZN(G160) );
  OR2_X1 U570 ( .A1(n709), .A2(n724), .ZN(n520) );
  XNOR2_X1 U571 ( .A(n622), .B(KEYINPUT26), .ZN(n624) );
  INV_X1 U572 ( .A(KEYINPUT27), .ZN(n613) );
  XNOR2_X1 U573 ( .A(n614), .B(n613), .ZN(n618) );
  INV_X1 U574 ( .A(KEYINPUT100), .ZN(n647) );
  BUF_X1 U575 ( .A(n615), .Z(n665) );
  BUF_X1 U576 ( .A(n612), .Z(n662) );
  AND2_X1 U577 ( .A1(n999), .A2(n520), .ZN(n710) );
  INV_X1 U578 ( .A(KEYINPUT0), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n639), .A2(G68), .ZN(n626) );
  INV_X1 U580 ( .A(G2105), .ZN(n535) );
  XNOR2_X1 U581 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n645) );
  XNOR2_X1 U582 ( .A(n630), .B(n629), .ZN(n633) );
  XNOR2_X1 U583 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U584 ( .A(n540), .B(n539), .ZN(n733) );
  NOR2_X1 U585 ( .A1(n608), .A2(n607), .ZN(n787) );
  XOR2_X1 U586 ( .A(KEYINPUT71), .B(n534), .Z(G299) );
  XOR2_X2 U587 ( .A(KEYINPUT65), .B(n522), .Z(n806) );
  NAND2_X1 U588 ( .A1(n806), .A2(G53), .ZN(n533) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n809) );
  NAND2_X1 U590 ( .A1(G91), .A2(n809), .ZN(n525) );
  INV_X1 U591 ( .A(G651), .ZN(n527) );
  NOR2_X1 U592 ( .A1(G543), .A2(n527), .ZN(n523) );
  XOR2_X2 U593 ( .A(KEYINPUT1), .B(n523), .Z(n805) );
  NAND2_X1 U594 ( .A1(G65), .A2(n805), .ZN(n524) );
  NAND2_X1 U595 ( .A1(n525), .A2(n524), .ZN(n531) );
  OR2_X1 U596 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X2 U597 ( .A(KEYINPUT66), .B(n528), .Z(n639) );
  NAND2_X1 U598 ( .A1(n639), .A2(G78), .ZN(n529) );
  XOR2_X1 U599 ( .A(KEYINPUT70), .B(n529), .Z(n530) );
  NOR2_X1 U600 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U602 ( .A1(n891), .A2(G113), .ZN(n538) );
  AND2_X4 U603 ( .A1(n535), .A2(G2104), .ZN(n895) );
  NAND2_X1 U604 ( .A1(G101), .A2(n895), .ZN(n536) );
  XOR2_X1 U605 ( .A(KEYINPUT23), .B(n536), .Z(n537) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n545) );
  NAND2_X1 U607 ( .A1(G137), .A2(n733), .ZN(n543) );
  INV_X1 U608 ( .A(G2104), .ZN(n541) );
  BUF_X1 U609 ( .A(n598), .Z(n892) );
  NAND2_X1 U610 ( .A1(G125), .A2(n892), .ZN(n542) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  BUF_X1 U612 ( .A(n639), .Z(n590) );
  NAND2_X1 U613 ( .A1(G77), .A2(n590), .ZN(n546) );
  XOR2_X1 U614 ( .A(KEYINPUT69), .B(n546), .Z(n548) );
  NAND2_X1 U615 ( .A1(n809), .A2(G90), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(KEYINPUT9), .ZN(n551) );
  NAND2_X1 U618 ( .A1(G52), .A2(n806), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n805), .A2(G64), .ZN(n552) );
  XOR2_X1 U621 ( .A(KEYINPUT68), .B(n552), .Z(n553) );
  NOR2_X1 U622 ( .A1(n554), .A2(n553), .ZN(G171) );
  NAND2_X1 U623 ( .A1(n809), .A2(G89), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U625 ( .A1(G76), .A2(n590), .ZN(n556) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n558), .B(KEYINPUT5), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n562) );
  NAND2_X1 U629 ( .A1(G63), .A2(n805), .ZN(n560) );
  NAND2_X1 U630 ( .A1(G51), .A2(n806), .ZN(n559) );
  NAND2_X1 U631 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U632 ( .A(n562), .B(n561), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(KEYINPUT7), .B(n565), .ZN(G168) );
  NAND2_X1 U635 ( .A1(G88), .A2(n809), .ZN(n566) );
  XNOR2_X1 U636 ( .A(n566), .B(KEYINPUT87), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G62), .A2(n805), .ZN(n568) );
  NAND2_X1 U638 ( .A1(G50), .A2(n806), .ZN(n567) );
  NAND2_X1 U639 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U640 ( .A(KEYINPUT86), .B(n569), .Z(n571) );
  NAND2_X1 U641 ( .A1(G75), .A2(n590), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U643 ( .A1(n573), .A2(n572), .ZN(G166) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U645 ( .A(G166), .ZN(G303) );
  NAND2_X1 U646 ( .A1(G49), .A2(n806), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n574), .B(KEYINPUT82), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G87), .A2(n526), .ZN(n576) );
  NAND2_X1 U649 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U651 ( .A1(n805), .A2(n577), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U653 ( .A1(G86), .A2(n809), .ZN(n581) );
  NAND2_X1 U654 ( .A1(G61), .A2(n805), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n583) );
  NAND2_X1 U657 ( .A1(G73), .A2(n590), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U659 ( .A(KEYINPUT83), .B(n584), .Z(n585) );
  NOR2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U661 ( .A(KEYINPUT85), .B(n587), .Z(n589) );
  NAND2_X1 U662 ( .A1(n806), .A2(G48), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(G305) );
  NAND2_X1 U664 ( .A1(G72), .A2(n590), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n809), .A2(G85), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U667 ( .A(KEYINPUT67), .B(n593), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G60), .A2(n805), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G47), .A2(n806), .ZN(n594) );
  AND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G290) );
  NAND2_X1 U672 ( .A1(G160), .A2(G40), .ZN(n730) );
  NAND2_X1 U673 ( .A1(G126), .A2(n598), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT90), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n733), .A2(G138), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G102), .A2(n895), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n787), .A2(G1384), .ZN(n610) );
  INV_X1 U680 ( .A(KEYINPUT64), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n610), .B(n609), .ZN(n728) );
  NOR2_X2 U682 ( .A1(n730), .A2(n728), .ZN(n612) );
  INV_X1 U683 ( .A(KEYINPUT97), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n615), .A2(G2072), .ZN(n614) );
  INV_X1 U686 ( .A(n665), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n616), .A2(G1956), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT99), .ZN(n656) );
  INV_X1 U690 ( .A(G299), .ZN(n817) );
  NOR2_X2 U691 ( .A1(n656), .A2(n817), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(n620), .ZN(n660) );
  NAND2_X1 U693 ( .A1(n662), .A2(G1996), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n680), .A2(G1341), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n636) );
  NAND2_X1 U696 ( .A1(n809), .A2(G81), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT12), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n805), .A2(G56), .ZN(n631) );
  XOR2_X1 U701 ( .A(KEYINPUT14), .B(n631), .Z(n632) );
  NOR2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U703 ( .A1(n806), .A2(G43), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n994) );
  NOR2_X1 U705 ( .A1(n636), .A2(n994), .ZN(n649) );
  NAND2_X1 U706 ( .A1(G54), .A2(n806), .ZN(n644) );
  NAND2_X1 U707 ( .A1(G92), .A2(n809), .ZN(n638) );
  NAND2_X1 U708 ( .A1(G66), .A2(n805), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U710 ( .A1(G79), .A2(n639), .ZN(n640) );
  XNOR2_X1 U711 ( .A(KEYINPUT77), .B(n640), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X2 U714 ( .A(n646), .B(n645), .ZN(n993) );
  NOR2_X1 U715 ( .A1(n649), .A2(n993), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(n655) );
  NAND2_X1 U717 ( .A1(n649), .A2(n993), .ZN(n653) );
  NAND2_X1 U718 ( .A1(G2067), .A2(n665), .ZN(n651) );
  NAND2_X1 U719 ( .A1(G1348), .A2(n680), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n817), .A2(n656), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U726 ( .A(n661), .B(KEYINPUT29), .ZN(n669) );
  NOR2_X1 U727 ( .A1(n662), .A2(G1961), .ZN(n663) );
  XOR2_X1 U728 ( .A(KEYINPUT96), .B(n663), .Z(n667) );
  XNOR2_X1 U729 ( .A(G2078), .B(KEYINPUT25), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n664), .B(KEYINPUT98), .ZN(n964) );
  NAND2_X1 U731 ( .A1(n964), .A2(n665), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n674) );
  AND2_X1 U733 ( .A1(G171), .A2(n674), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT101), .ZN(n693) );
  NOR2_X1 U736 ( .A1(G1966), .A2(n724), .ZN(n695) );
  NOR2_X1 U737 ( .A1(G2084), .A2(n680), .ZN(n691) );
  NOR2_X1 U738 ( .A1(n695), .A2(n691), .ZN(n671) );
  NAND2_X1 U739 ( .A1(G8), .A2(n671), .ZN(n672) );
  XNOR2_X1 U740 ( .A(KEYINPUT30), .B(n672), .ZN(n673) );
  NOR2_X1 U741 ( .A1(G168), .A2(n673), .ZN(n676) );
  NOR2_X1 U742 ( .A1(G171), .A2(n674), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U744 ( .A(KEYINPUT31), .B(n677), .Z(n692) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n724), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(KEYINPUT102), .ZN(n679) );
  NOR2_X1 U747 ( .A1(G166), .A2(n679), .ZN(n683) );
  NOR2_X1 U748 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(KEYINPUT103), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n685) );
  AND2_X1 U751 ( .A1(n692), .A2(n685), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n693), .A2(n684), .ZN(n689) );
  INV_X1 U753 ( .A(n685), .ZN(n686) );
  OR2_X1 U754 ( .A1(n686), .A2(G286), .ZN(n687) );
  AND2_X1 U755 ( .A1(n687), .A2(G8), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT32), .ZN(n699) );
  NAND2_X1 U758 ( .A1(G8), .A2(n691), .ZN(n697) );
  AND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n712), .B(KEYINPUT104), .ZN(n702) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n700) );
  NOR2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n987) );
  NOR2_X1 U766 ( .A1(n700), .A2(n987), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U768 ( .A1(G288), .A2(G1976), .ZN(n703) );
  XOR2_X1 U769 ( .A(KEYINPUT105), .B(n703), .Z(n988) );
  NAND2_X1 U770 ( .A1(n704), .A2(n988), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT106), .ZN(n706) );
  NOR2_X1 U772 ( .A1(n724), .A2(n706), .ZN(n707) );
  NOR2_X1 U773 ( .A1(KEYINPUT33), .A2(n707), .ZN(n708) );
  INV_X1 U774 ( .A(n708), .ZN(n711) );
  XOR2_X1 U775 ( .A(G1981), .B(G305), .Z(n999) );
  NAND2_X1 U776 ( .A1(n987), .A2(KEYINPUT33), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n720) );
  XOR2_X1 U778 ( .A(KEYINPUT104), .B(n712), .Z(n715) );
  NAND2_X1 U779 ( .A1(G166), .A2(G8), .ZN(n713) );
  NOR2_X1 U780 ( .A1(G2090), .A2(n713), .ZN(n714) );
  NOR2_X2 U781 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n716), .B(KEYINPUT107), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n717), .A2(n724), .ZN(n718) );
  XNOR2_X1 U784 ( .A(n718), .B(KEYINPUT108), .ZN(n719) );
  NAND2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n726) );
  NOR2_X1 U786 ( .A1(G1981), .A2(G305), .ZN(n721) );
  XNOR2_X1 U787 ( .A(KEYINPUT24), .B(n721), .ZN(n722) );
  XNOR2_X1 U788 ( .A(KEYINPUT95), .B(n722), .ZN(n723) );
  NOR2_X1 U789 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X2 U790 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U791 ( .A(n727), .B(KEYINPUT109), .ZN(n764) );
  XNOR2_X1 U792 ( .A(G1986), .B(G290), .ZN(n996) );
  INV_X1 U793 ( .A(n728), .ZN(n729) );
  NOR2_X1 U794 ( .A1(n730), .A2(n729), .ZN(n774) );
  NAND2_X1 U795 ( .A1(n996), .A2(n774), .ZN(n762) );
  NAND2_X1 U796 ( .A1(n895), .A2(G105), .ZN(n732) );
  XNOR2_X1 U797 ( .A(KEYINPUT38), .B(KEYINPUT94), .ZN(n731) );
  XNOR2_X1 U798 ( .A(n732), .B(n731), .ZN(n740) );
  BUF_X1 U799 ( .A(n733), .Z(n896) );
  NAND2_X1 U800 ( .A1(G141), .A2(n896), .ZN(n735) );
  NAND2_X1 U801 ( .A1(G129), .A2(n892), .ZN(n734) );
  NAND2_X1 U802 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U803 ( .A1(G117), .A2(n891), .ZN(n736) );
  XNOR2_X1 U804 ( .A(KEYINPUT93), .B(n736), .ZN(n737) );
  NOR2_X1 U805 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U806 ( .A1(n740), .A2(n739), .ZN(n873) );
  AND2_X1 U807 ( .A1(n873), .A2(G1996), .ZN(n748) );
  NAND2_X1 U808 ( .A1(G95), .A2(n895), .ZN(n742) );
  NAND2_X1 U809 ( .A1(G131), .A2(n896), .ZN(n741) );
  NAND2_X1 U810 ( .A1(n742), .A2(n741), .ZN(n746) );
  NAND2_X1 U811 ( .A1(G107), .A2(n891), .ZN(n744) );
  NAND2_X1 U812 ( .A1(G119), .A2(n892), .ZN(n743) );
  NAND2_X1 U813 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U814 ( .A1(n746), .A2(n745), .ZN(n904) );
  INV_X1 U815 ( .A(G1991), .ZN(n958) );
  NOR2_X1 U816 ( .A1(n904), .A2(n958), .ZN(n747) );
  NOR2_X1 U817 ( .A1(n748), .A2(n747), .ZN(n937) );
  INV_X1 U818 ( .A(n774), .ZN(n749) );
  NOR2_X1 U819 ( .A1(n937), .A2(n749), .ZN(n767) );
  XNOR2_X1 U820 ( .A(KEYINPUT37), .B(G2067), .ZN(n772) );
  NAND2_X1 U821 ( .A1(G116), .A2(n891), .ZN(n751) );
  NAND2_X1 U822 ( .A1(G128), .A2(n892), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U824 ( .A(n752), .B(KEYINPUT35), .ZN(n757) );
  NAND2_X1 U825 ( .A1(G104), .A2(n895), .ZN(n754) );
  NAND2_X1 U826 ( .A1(G140), .A2(n896), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U828 ( .A(KEYINPUT34), .B(n755), .Z(n756) );
  NAND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U830 ( .A(n758), .B(KEYINPUT36), .Z(n884) );
  OR2_X1 U831 ( .A1(n772), .A2(n884), .ZN(n759) );
  XOR2_X1 U832 ( .A(KEYINPUT92), .B(n759), .Z(n940) );
  NAND2_X1 U833 ( .A1(n774), .A2(n940), .ZN(n770) );
  INV_X1 U834 ( .A(n770), .ZN(n760) );
  NOR2_X1 U835 ( .A1(n767), .A2(n760), .ZN(n761) );
  AND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n777) );
  NOR2_X1 U838 ( .A1(G1996), .A2(n873), .ZN(n945) );
  AND2_X1 U839 ( .A1(n958), .A2(n904), .ZN(n933) );
  NOR2_X1 U840 ( .A1(G1986), .A2(G290), .ZN(n765) );
  NOR2_X1 U841 ( .A1(n933), .A2(n765), .ZN(n766) );
  NOR2_X1 U842 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U843 ( .A1(n945), .A2(n768), .ZN(n769) );
  XNOR2_X1 U844 ( .A(n769), .B(KEYINPUT39), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U846 ( .A1(n884), .A2(n772), .ZN(n943) );
  NAND2_X1 U847 ( .A1(n773), .A2(n943), .ZN(n775) );
  NAND2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U849 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U850 ( .A(n778), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U851 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U852 ( .A1(G111), .A2(n891), .ZN(n780) );
  NAND2_X1 U853 ( .A1(G135), .A2(n896), .ZN(n779) );
  NAND2_X1 U854 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U855 ( .A1(n892), .A2(G123), .ZN(n781) );
  XOR2_X1 U856 ( .A(KEYINPUT18), .B(n781), .Z(n782) );
  NOR2_X1 U857 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U858 ( .A1(n895), .A2(G99), .ZN(n784) );
  NAND2_X1 U859 ( .A1(n785), .A2(n784), .ZN(n934) );
  XNOR2_X1 U860 ( .A(G2096), .B(n934), .ZN(n786) );
  OR2_X1 U861 ( .A1(G2100), .A2(n786), .ZN(G156) );
  INV_X1 U862 ( .A(G82), .ZN(G220) );
  INV_X1 U863 ( .A(G120), .ZN(G236) );
  BUF_X1 U864 ( .A(n787), .Z(G164) );
  NAND2_X1 U865 ( .A1(G7), .A2(G661), .ZN(n788) );
  XNOR2_X1 U866 ( .A(n788), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U867 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n790) );
  INV_X1 U868 ( .A(G223), .ZN(n840) );
  NAND2_X1 U869 ( .A1(G567), .A2(n840), .ZN(n789) );
  XNOR2_X1 U870 ( .A(n790), .B(n789), .ZN(G234) );
  INV_X1 U871 ( .A(G860), .ZN(n804) );
  OR2_X1 U872 ( .A1(n994), .A2(n804), .ZN(G153) );
  INV_X1 U873 ( .A(G171), .ZN(G301) );
  INV_X1 U874 ( .A(G868), .ZN(n798) );
  AND2_X1 U875 ( .A1(n993), .A2(n798), .ZN(n792) );
  NOR2_X1 U876 ( .A1(n798), .A2(G301), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(G284) );
  NOR2_X1 U878 ( .A1(G868), .A2(G299), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n793), .B(KEYINPUT80), .ZN(n795) );
  NOR2_X1 U880 ( .A1(n798), .A2(G286), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(G297) );
  NAND2_X1 U882 ( .A1(n804), .A2(G559), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n796), .A2(n993), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U885 ( .A1(G559), .A2(n798), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n799), .A2(n993), .ZN(n800) );
  XNOR2_X1 U887 ( .A(n800), .B(KEYINPUT81), .ZN(n802) );
  NOR2_X1 U888 ( .A1(n994), .A2(G868), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(G282) );
  NAND2_X1 U890 ( .A1(n993), .A2(G559), .ZN(n803) );
  XOR2_X1 U891 ( .A(n994), .B(n803), .Z(n821) );
  NAND2_X1 U892 ( .A1(n804), .A2(n821), .ZN(n814) );
  NAND2_X1 U893 ( .A1(G67), .A2(n805), .ZN(n808) );
  NAND2_X1 U894 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n808), .A2(n807), .ZN(n813) );
  NAND2_X1 U896 ( .A1(G93), .A2(n809), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G80), .A2(n590), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U899 ( .A1(n813), .A2(n812), .ZN(n823) );
  XOR2_X1 U900 ( .A(n814), .B(n823), .Z(G145) );
  XOR2_X1 U901 ( .A(KEYINPUT19), .B(n823), .Z(n815) );
  XNOR2_X1 U902 ( .A(G288), .B(n815), .ZN(n816) );
  XNOR2_X1 U903 ( .A(n817), .B(n816), .ZN(n819) );
  XNOR2_X1 U904 ( .A(G290), .B(G166), .ZN(n818) );
  XNOR2_X1 U905 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U906 ( .A(n820), .B(G305), .ZN(n908) );
  XNOR2_X1 U907 ( .A(n821), .B(n908), .ZN(n822) );
  NAND2_X1 U908 ( .A1(n822), .A2(G868), .ZN(n825) );
  OR2_X1 U909 ( .A1(G868), .A2(n823), .ZN(n824) );
  NAND2_X1 U910 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(n826), .Z(n827) );
  NAND2_X1 U913 ( .A1(G2090), .A2(n827), .ZN(n828) );
  XNOR2_X1 U914 ( .A(KEYINPUT21), .B(n828), .ZN(n829) );
  NAND2_X1 U915 ( .A1(n829), .A2(G2072), .ZN(G158) );
  XOR2_X1 U916 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U918 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NOR2_X1 U919 ( .A1(G237), .A2(G236), .ZN(n830) );
  NAND2_X1 U920 ( .A1(G69), .A2(n830), .ZN(n831) );
  XNOR2_X1 U921 ( .A(KEYINPUT89), .B(n831), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n832), .A2(G108), .ZN(n844) );
  NAND2_X1 U923 ( .A1(n844), .A2(G567), .ZN(n838) );
  NOR2_X1 U924 ( .A1(G220), .A2(G219), .ZN(n833) );
  XOR2_X1 U925 ( .A(KEYINPUT22), .B(n833), .Z(n834) );
  NOR2_X1 U926 ( .A1(G218), .A2(n834), .ZN(n835) );
  NAND2_X1 U927 ( .A1(G96), .A2(n835), .ZN(n845) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n845), .ZN(n836) );
  XNOR2_X1 U929 ( .A(KEYINPUT88), .B(n836), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(n847) );
  NAND2_X1 U931 ( .A1(G661), .A2(G483), .ZN(n839) );
  NOR2_X1 U932 ( .A1(n847), .A2(n839), .ZN(n843) );
  NAND2_X1 U933 ( .A1(n843), .A2(G36), .ZN(G176) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U936 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n843), .A2(n842), .ZN(G188) );
  INV_X1 U940 ( .A(G108), .ZN(G238) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  NOR2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n846), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  INV_X1 U945 ( .A(n847), .ZN(G319) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1956), .B(G1961), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1976), .B(G1971), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U958 ( .A(G1966), .B(G1981), .Z(n859) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U962 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U964 ( .A(G1986), .B(G2474), .Z(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n892), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n891), .A2(G112), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G100), .A2(n895), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G136), .A2(n896), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(G162) );
  XNOR2_X1 U974 ( .A(G162), .B(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(G160), .B(G164), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n934), .B(n876), .ZN(n886) );
  NAND2_X1 U978 ( .A1(G103), .A2(n895), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G139), .A2(n896), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G115), .A2(n891), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G127), .A2(n892), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n928) );
  XOR2_X1 U986 ( .A(n884), .B(n928), .Z(n885) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U988 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n888) );
  XNOR2_X1 U989 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U991 ( .A(n890), .B(n889), .Z(n906) );
  NAND2_X1 U992 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G130), .A2(n892), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U995 ( .A1(G106), .A2(n895), .ZN(n898) );
  NAND2_X1 U996 ( .A1(G142), .A2(n896), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(n899), .Z(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT45), .B(n900), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n908), .B(n993), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n909), .B(n994), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(G286), .B(G171), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n912), .ZN(G397) );
  XOR2_X1 U1009 ( .A(G2451), .B(G2430), .Z(n914) );
  XNOR2_X1 U1010 ( .A(G2438), .B(G2443), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n920) );
  XOR2_X1 U1012 ( .A(G2435), .B(G2454), .Z(n916) );
  XNOR2_X1 U1013 ( .A(G1341), .B(G1348), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1015 ( .A(G2446), .B(G2427), .Z(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1017 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n921), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  INV_X1 U1027 ( .A(n927), .ZN(G401) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n977) );
  XOR2_X1 U1029 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(KEYINPUT50), .B(n931), .ZN(n951) );
  XOR2_X1 U1033 ( .A(G160), .B(G2084), .Z(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT115), .B(n936), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n941), .B(KEYINPUT116), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G162), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(KEYINPUT117), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT51), .B(n947), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n952), .B(KEYINPUT52), .ZN(n953) );
  XOR2_X1 U1048 ( .A(KEYINPUT118), .B(n953), .Z(n954) );
  NAND2_X1 U1049 ( .A1(n977), .A2(n954), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(G29), .ZN(n1037) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n956), .ZN(n975) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G35), .ZN(n973) );
  XNOR2_X1 U1054 ( .A(KEYINPUT119), .B(G2067), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(n957), .B(G26), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G25), .B(n958), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n959), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n969) );
  XOR2_X1 U1061 ( .A(n964), .B(G27), .Z(n966) );
  XNOR2_X1 U1062 ( .A(G32), .B(G1996), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1064 ( .A(n967), .B(KEYINPUT120), .Z(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1066 ( .A(KEYINPUT53), .B(n970), .Z(n971) );
  XNOR2_X1 U1067 ( .A(n971), .B(KEYINPUT121), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT122), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n978), .B(n977), .ZN(n980) );
  INV_X1 U1072 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(G11), .A2(n981), .ZN(n1035) );
  INV_X1 U1075 ( .A(G16), .ZN(n1031) );
  XNOR2_X1 U1076 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(n1031), .B(n982), .ZN(n1007) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G166), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G301), .B(G1961), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(G299), .B(G1956), .ZN(n983) );
  NOR2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n992) );
  INV_X1 U1083 ( .A(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(KEYINPUT124), .B(n990), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n1005) );
  XNOR2_X1 U1087 ( .A(G1348), .B(n993), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(G1341), .B(n994), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1093 ( .A(KEYINPUT57), .B(n1001), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1033) );
  XOR2_X1 U1097 ( .A(G1348), .B(KEYINPUT59), .Z(n1008) );
  XNOR2_X1 U1098 ( .A(G4), .B(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G6), .B(G1981), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G19), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G1956), .B(G20), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(KEYINPUT125), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(KEYINPUT60), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G1966), .B(G21), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(G5), .B(G1961), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(G1986), .B(G24), .ZN(n1022) );
  XNOR2_X1 U1112 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1113 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
  XOR2_X1 U1114 ( .A(G1971), .B(KEYINPUT126), .Z(n1023) );
  XNOR2_X1 U1115 ( .A(G22), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1117 ( .A(KEYINPUT58), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1118 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1119 ( .A(KEYINPUT61), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1038), .Z(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

