//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928;
  XNOR2_X1  g000(.A(G176gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT108), .B(G120gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G230gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT10), .ZN(new_n210));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT98), .ZN(new_n212));
  NAND2_X1  g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  OR2_X1    g012(.A1(G71gat), .A2(G78gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n214), .C1(new_n211), .C2(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT102), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT7), .ZN(new_n221));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222));
  XOR2_X1   g021(.A(new_n221), .B(new_n222), .Z(new_n223));
  INV_X1    g022(.A(G99gat), .ZN(new_n224));
  INV_X1    g023(.A(G106gat), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT103), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT103), .B1(new_n224), .B2(new_n225), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(KEYINPUT8), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT104), .B(G85gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n223), .B(new_n228), .C1(G92gat), .C2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G99gat), .B(G106gat), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT106), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n219), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n231), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n230), .B(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(KEYINPUT106), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n219), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n210), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n232), .A2(new_n210), .A3(new_n219), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n209), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n238), .A2(new_n208), .A3(new_n241), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n207), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT109), .ZN(new_n248));
  INV_X1    g047(.A(new_n246), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT107), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(new_n244), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n246), .B1(new_n252), .B2(new_n208), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n206), .C1(new_n253), .C2(new_n250), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G22gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G197gat), .B(G204gat), .Z(new_n261));
  INV_X1    g060(.A(KEYINPUT22), .ZN(new_n262));
  NAND2_X1  g061(.A1(G211gat), .A2(G218gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT73), .ZN(new_n265));
  INV_X1    g064(.A(new_n263), .ZN(new_n266));
  NOR2_X1   g065(.A1(G211gat), .A2(G218gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n265), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(new_n274), .B2(KEYINPUT2), .ZN(new_n275));
  INV_X1    g074(.A(G141gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT79), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G141gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n203), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n276), .A2(G148gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G141gat), .B(G148gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n271), .B(new_n274), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G228gat), .A2(G233gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT87), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n282), .A2(new_n285), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT81), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n285), .A3(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n264), .A2(new_n268), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n264), .A2(new_n268), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n289), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT86), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n287), .B1(new_n303), .B2(new_n304), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n298), .B(new_n300), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n294), .A2(new_n296), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n265), .B(new_n268), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n289), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n286), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n293), .B1(new_n312), .B2(new_n292), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT31), .B(G50gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n308), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n308), .B2(new_n313), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n260), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n308), .A2(new_n313), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n314), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(new_n259), .A3(new_n316), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n300), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n299), .B1(new_n282), .B2(new_n285), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  INV_X1    g126(.A(G134gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT67), .ZN(new_n329));
  XNOR2_X1  g128(.A(G113gat), .B(G120gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(KEYINPUT1), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G120gat), .ZN(new_n334));
  INV_X1    g133(.A(G120gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(G113gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n332), .B(new_n328), .C1(new_n334), .C2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n327), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n331), .A2(new_n327), .A3(new_n337), .ZN(new_n339));
  OAI22_X1  g138(.A1(new_n325), .A2(new_n326), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n339), .A2(new_n338), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n288), .B(new_n343), .C1(new_n311), .C2(new_n286), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n331), .A2(new_n337), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G127gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n327), .A3(new_n337), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n297), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n342), .B(new_n344), .C1(new_n341), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n350), .A2(KEYINPUT5), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n298), .A2(new_n300), .B1(new_n346), .B2(new_n347), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n341), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n340), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n348), .A2(new_n341), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n344), .A2(new_n351), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n286), .A2(new_n339), .A3(new_n338), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n352), .B1(new_n363), .B2(new_n348), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT83), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n352), .C1(new_n363), .C2(new_n348), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n362), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n361), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n353), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G57gat), .B(G85gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n377), .B(new_n353), .C1(new_n370), .C2(new_n371), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(KEYINPUT6), .A3(new_n378), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n385));
  NOR2_X1   g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(KEYINPUT23), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  AOI22_X1  g190(.A1(KEYINPUT66), .A2(new_n391), .B1(new_n386), .B2(KEYINPUT23), .ZN(new_n392));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT24), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n391), .A2(KEYINPUT66), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n390), .A2(new_n392), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT25), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT26), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT27), .B(G183gat), .ZN(new_n407));
  INV_X1    g206(.A(G190gat), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT28), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT28), .B(new_n408), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n393), .B(new_n406), .C1(new_n409), .C2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n395), .A2(new_n396), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT64), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT25), .B1(new_n386), .B2(KEYINPUT23), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n404), .A3(new_n390), .A4(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n401), .A2(new_n414), .A3(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n424), .B(KEYINPUT74), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n423), .A2(new_n289), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n309), .B(new_n427), .C1(new_n428), .C2(new_n424), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n429), .A2(KEYINPUT76), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n423), .A2(new_n424), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n428), .A2(new_n426), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n309), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G8gat), .B(G36gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n438), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT77), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n435), .A2(new_n436), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n270), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(new_n431), .A3(new_n430), .A4(new_n442), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n441), .B1(new_n432), .B2(new_n437), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n443), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n324), .B1(new_n384), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n423), .A2(new_n343), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n423), .A2(new_n343), .ZN(new_n458));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n423), .A2(KEYINPUT68), .A3(new_n343), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT34), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n461), .A2(KEYINPUT34), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n469));
  INV_X1    g268(.A(new_n459), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT33), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT69), .B(G71gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G43gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n471), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  AOI221_X4 g277(.A(new_n468), .B1(KEYINPUT33), .B2(new_n476), .C1(new_n469), .C2(new_n470), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n467), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n461), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT70), .B1(new_n461), .B2(KEYINPUT34), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n423), .A2(KEYINPUT68), .A3(new_n343), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT68), .B1(new_n423), .B2(new_n343), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n423), .A2(new_n343), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT32), .B1(new_n487), .B2(new_n459), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n487), .B2(new_n459), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(new_n476), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n471), .B1(new_n472), .B2(new_n477), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n483), .A2(new_n491), .A3(new_n492), .A4(new_n465), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n480), .A2(new_n493), .A3(KEYINPUT72), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n467), .C1(new_n478), .C2(new_n479), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n493), .A3(KEYINPUT71), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT71), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n467), .C1(new_n478), .C2(new_n479), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(KEYINPUT36), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT88), .B1(new_n454), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n500), .A2(KEYINPUT36), .A3(new_n502), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT36), .B1(new_n494), .B2(new_n496), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n452), .B1(new_n383), .B2(new_n382), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n324), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT37), .B1(new_n432), .B2(new_n437), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n446), .A2(new_n513), .A3(new_n431), .A4(new_n430), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n441), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n515), .A2(new_n516), .B1(new_n438), .B2(new_n442), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n445), .A2(new_n309), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n270), .B(new_n427), .C1(new_n428), .C2(new_n424), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(KEYINPUT37), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n516), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n514), .A2(new_n520), .A3(new_n441), .A4(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n517), .A2(new_n382), .A3(new_n383), .A4(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT39), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n350), .A2(new_n524), .A3(new_n352), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n525), .A2(new_n377), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n350), .A2(new_n352), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n363), .A2(new_n348), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(KEYINPUT39), .C1(new_n352), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT40), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n526), .A2(new_n529), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT40), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n452), .A2(new_n532), .A3(new_n379), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n523), .A2(new_n535), .A3(new_n324), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n505), .A2(new_n511), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n323), .B1(new_n502), .B2(new_n500), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n324), .B(new_n497), .C1(new_n510), .C2(KEYINPUT91), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n384), .A2(new_n453), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n540), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n257), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(KEYINPUT93), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT15), .ZN(new_n553));
  INV_X1    g352(.A(G29gat), .ZN(new_n554));
  INV_X1    g353(.A(G36gat), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR3_X1   g356(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT94), .ZN(new_n559));
  OAI221_X1 g358(.A(new_n553), .B1(new_n554), .B2(new_n555), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  OAI22_X1  g359(.A1(new_n557), .A2(new_n558), .B1(new_n554), .B2(new_n555), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT15), .A3(new_n551), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n549), .B(new_n550), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n549), .A2(new_n550), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n550), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(new_n562), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n232), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n560), .A2(new_n562), .ZN(new_n570));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT100), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n570), .A2(new_n236), .B1(KEYINPUT41), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G190gat), .B(G218gat), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT105), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n578), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n569), .A2(new_n581), .A3(new_n574), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(KEYINPUT101), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n548), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n548), .A3(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n239), .A2(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G211gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G15gat), .B(G22gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT16), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(G1gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(G1gat), .B2(new_n597), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G8gat), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n239), .B2(KEYINPUT21), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n596), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT99), .B(G183gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n605), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n570), .A2(KEYINPUT95), .A3(KEYINPUT17), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n601), .B1(new_n611), .B2(new_n567), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n570), .A2(new_n601), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n570), .B(new_n601), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n613), .B(KEYINPUT13), .Z(new_n619));
  AOI22_X1  g418(.A1(new_n617), .A2(KEYINPUT18), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n617), .B2(KEYINPUT18), .ZN(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G197gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT11), .B(G169gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT92), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  INV_X1    g427(.A(new_n601), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n563), .B2(new_n568), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(new_n613), .A3(new_n615), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT18), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(KEYINPUT97), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n620), .A2(new_n622), .A3(new_n628), .A4(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n631), .A2(KEYINPUT96), .A3(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n619), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n631), .B2(new_n632), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT96), .B1(new_n631), .B2(new_n632), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n634), .B1(new_n639), .B2(new_n628), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n610), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n547), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n384), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g445(.A1(new_n643), .A2(new_n452), .ZN(new_n647));
  NAND2_X1  g446(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n648));
  INV_X1    g447(.A(G8gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n598), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n653), .B(new_n654), .C1(new_n649), .C2(new_n647), .ZN(G1325gat));
  AOI21_X1  g454(.A(G15gat), .B1(new_n643), .B2(new_n497), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n504), .A2(G15gat), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n643), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n323), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  AOI21_X1  g460(.A(new_n591), .B1(new_n537), .B2(new_n546), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n257), .A2(new_n641), .A3(new_n609), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n554), .A3(new_n644), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT45), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n508), .B1(new_n510), .B2(new_n324), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n523), .A2(new_n535), .A3(new_n324), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT110), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n454), .A2(new_n504), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n536), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n324), .A2(new_n497), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n543), .B2(new_n544), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT35), .B1(new_n510), .B2(KEYINPUT91), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n670), .A2(new_n673), .B1(new_n540), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n667), .B1(new_n678), .B2(new_n591), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n663), .ZN(new_n681));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681), .B2(new_n384), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n682), .ZN(G1328gat));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n555), .A3(new_n452), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT46), .Z(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n681), .B2(new_n453), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1329gat));
  XOR2_X1   g486(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n537), .A2(new_n546), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n586), .A2(new_n548), .A3(new_n587), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n588), .ZN(new_n692));
  INV_X1    g491(.A(new_n497), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n690), .A2(new_n692), .A3(new_n663), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT112), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT112), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n662), .A2(new_n697), .A3(new_n663), .A4(new_n694), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n696), .A2(KEYINPUT113), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT113), .B1(new_n696), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G43gat), .B1(new_n681), .B2(new_n508), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n689), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n696), .A2(new_n698), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT114), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT113), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n696), .A2(KEYINPUT113), .A3(new_n698), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n702), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n688), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT114), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n704), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n706), .A2(new_n714), .ZN(G1330gat));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716));
  OAI21_X1  g515(.A(G50gat), .B1(new_n681), .B2(new_n324), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT115), .ZN(new_n718));
  INV_X1    g517(.A(G50gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n664), .A2(new_n719), .A3(new_n323), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n723), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(KEYINPUT48), .A3(new_n721), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1331gat));
  NOR3_X1   g526(.A1(new_n678), .A2(new_n640), .A3(new_n610), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n257), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n644), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g531(.A(new_n453), .B(new_n729), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n729), .B2(new_n508), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n693), .A2(G71gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g538(.A1(new_n730), .A2(new_n323), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n609), .A2(new_n640), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n679), .A2(new_n257), .A3(new_n680), .A4(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n229), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n743), .A2(new_n384), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n670), .A2(new_n673), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n546), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n692), .A3(new_n742), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT51), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n747), .A2(new_n750), .A3(new_n692), .A4(new_n742), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n644), .A3(new_n257), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n745), .B1(new_n753), .B2(new_n744), .ZN(G1336gat));
  OAI21_X1  g553(.A(G92gat), .B1(new_n743), .B2(new_n453), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n453), .A2(G92gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n749), .A2(new_n751), .A3(new_n257), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760));
  OR3_X1    g559(.A1(new_n743), .A2(new_n760), .A3(new_n508), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n743), .B2(new_n508), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(G99gat), .A3(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n752), .A2(new_n224), .A3(new_n497), .A4(new_n257), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1338gat));
  NOR2_X1   g564(.A1(new_n324), .A2(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n257), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT117), .Z(new_n768));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G106gat), .B1(new_n743), .B2(new_n324), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n749), .A2(new_n751), .A3(new_n257), .A4(new_n766), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n772), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n771), .A2(new_n772), .B1(new_n775), .B2(new_n776), .ZN(G1339gat));
  INV_X1    g576(.A(new_n609), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n206), .B1(new_n245), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n242), .A2(new_n209), .A3(new_n244), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n232), .A2(new_n233), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n236), .A2(KEYINPUT106), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n783), .A3(new_n219), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT10), .B1(new_n784), .B2(new_n240), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n208), .B1(new_n785), .B2(new_n243), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n781), .A2(new_n786), .A3(KEYINPUT54), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n254), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n780), .A2(new_n787), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n788), .A2(new_n254), .A3(KEYINPUT119), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n791), .A2(new_n640), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n626), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n613), .B1(new_n630), .B2(new_n615), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n618), .A2(new_n619), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n634), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n248), .B2(new_n255), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n692), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n791), .A2(new_n801), .A3(new_n794), .A4(new_n795), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n591), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n778), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n591), .A2(new_n641), .A3(new_n609), .A4(new_n256), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n674), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n384), .A2(new_n452), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT120), .Z(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n641), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n807), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n538), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n809), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n333), .A3(new_n640), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(G1340gat));
  OAI21_X1  g616(.A(G120gat), .B1(new_n811), .B2(new_n256), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n335), .A3(new_n257), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1341gat));
  XOR2_X1   g619(.A(KEYINPUT67), .B(G127gat), .Z(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n815), .B2(new_n609), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n811), .A2(new_n778), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n821), .ZN(G1342gat));
  OAI21_X1  g623(.A(G134gat), .B1(new_n811), .B2(new_n591), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n815), .A2(new_n328), .A3(new_n692), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(G1343gat));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n323), .ZN(new_n830));
  XOR2_X1   g629(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n788), .A2(new_n254), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT122), .B1(new_n792), .B2(new_n793), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n836), .B(KEYINPUT55), .C1(new_n780), .C2(new_n787), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n834), .B(new_n640), .C1(new_n835), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n802), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n591), .ZN(new_n840));
  INV_X1    g639(.A(new_n795), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT119), .B1(new_n788), .B2(new_n254), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n692), .A3(new_n801), .A4(new_n794), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n609), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n807), .ZN(new_n846));
  OAI211_X1 g645(.A(KEYINPUT57), .B(new_n323), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT123), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n692), .B1(new_n838), .B2(new_n802), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n778), .B1(new_n849), .B2(new_n805), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n324), .B1(new_n850), .B2(new_n807), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT57), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n508), .A2(new_n809), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n640), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n277), .A2(new_n279), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n830), .A2(new_n855), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n276), .A3(new_n640), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT58), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1344gat));
  OR2_X1    g665(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n324), .B1(new_n806), .B2(new_n807), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n831), .ZN(new_n869));
  AOI211_X1 g668(.A(new_n256), .B(new_n855), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT59), .B1(new_n870), .B2(new_n203), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n257), .A3(new_n856), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(G148gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n203), .A3(new_n257), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1345gat));
  AOI21_X1  g676(.A(G155gat), .B1(new_n860), .B2(new_n609), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n854), .A2(new_n856), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n778), .A2(new_n272), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(G1346gat));
  AOI21_X1  g680(.A(G162gat), .B1(new_n860), .B2(new_n692), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n591), .A2(new_n273), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n879), .B2(new_n883), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n644), .A2(new_n453), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n808), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G169gat), .B1(new_n886), .B2(new_n641), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n814), .A2(new_n885), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n641), .A2(G169gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1348gat));
  NOR2_X1   g689(.A1(new_n888), .A2(new_n256), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n257), .A2(G176gat), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n891), .A2(G176gat), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT124), .Z(G1349gat));
  OAI21_X1  g693(.A(G183gat), .B1(new_n886), .B2(new_n778), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n609), .A2(new_n407), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n897), .B(new_n898), .Z(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n886), .B2(new_n591), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(KEYINPUT61), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(KEYINPUT61), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n692), .A2(new_n408), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n901), .A2(new_n902), .B1(new_n888), .B2(new_n903), .ZN(G1351gat));
  NOR3_X1   g703(.A1(new_n504), .A2(new_n644), .A3(new_n453), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n868), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G197gat), .B1(new_n906), .B2(new_n640), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n905), .B(KEYINPUT126), .Z(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n867), .B2(new_n869), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n640), .A2(G197gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(G1352gat));
  NAND2_X1  g710(.A1(new_n867), .A2(new_n869), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n257), .ZN(new_n913));
  OAI21_X1  g712(.A(G204gat), .B1(new_n913), .B2(new_n908), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n868), .A2(new_n905), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(G204gat), .A3(new_n256), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n915), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(KEYINPUT127), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(KEYINPUT127), .ZN(new_n920));
  OAI221_X1 g719(.A(new_n914), .B1(new_n915), .B2(new_n917), .C1(new_n919), .C2(new_n920), .ZN(G1353gat));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n595), .A3(new_n609), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n912), .A2(new_n609), .A3(new_n905), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n923), .B2(G211gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n906), .B2(new_n692), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n692), .A2(G218gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n909), .B2(new_n928), .ZN(G1355gat));
endmodule


