

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789;

  NAND2_X1 U367 ( .A1(n414), .A2(n353), .ZN(n385) );
  INV_X1 U368 ( .A(n651), .ZN(n652) );
  XNOR2_X1 U369 ( .A(n646), .B(n415), .ZN(n414) );
  NOR2_X2 U370 ( .A1(n593), .A2(n600), .ZN(n571) );
  NAND2_X2 U371 ( .A1(n345), .A2(n406), .ZN(n619) );
  XNOR2_X2 U372 ( .A(n637), .B(n428), .ZN(n732) );
  XNOR2_X2 U373 ( .A(n367), .B(n397), .ZN(n362) );
  NOR2_X1 U374 ( .A1(n623), .A2(n557), .ZN(n558) );
  XNOR2_X1 U375 ( .A(n558), .B(KEYINPUT0), .ZN(n572) );
  AND2_X1 U376 ( .A1(n391), .A2(n698), .ZN(n390) );
  XNOR2_X1 U377 ( .A(n477), .B(n476), .ZN(n595) );
  XNOR2_X1 U378 ( .A(n539), .B(n538), .ZN(n770) );
  XNOR2_X1 U379 ( .A(G146), .B(G125), .ZN(n541) );
  NAND2_X1 U380 ( .A1(n399), .A2(n398), .ZN(n789) );
  NAND2_X1 U381 ( .A1(n421), .A2(n347), .ZN(n578) );
  AND2_X1 U382 ( .A1(n401), .A2(n400), .ZN(n399) );
  XNOR2_X1 U383 ( .A(n574), .B(n357), .ZN(n421) );
  BUF_X1 U384 ( .A(n572), .Z(n573) );
  NAND2_X1 U385 ( .A1(n572), .A2(n561), .ZN(n563) );
  AND2_X1 U386 ( .A1(n461), .A2(n457), .ZN(n456) );
  NAND2_X1 U387 ( .A1(n434), .A2(n437), .ZN(n433) );
  XNOR2_X1 U388 ( .A(n548), .B(n547), .ZN(n663) );
  XNOR2_X1 U389 ( .A(n498), .B(KEYINPUT25), .ZN(n499) );
  XNOR2_X1 U390 ( .A(n777), .B(G146), .ZN(n397) );
  XNOR2_X1 U391 ( .A(n471), .B(G134), .ZN(n777) );
  NOR2_X1 U392 ( .A1(n460), .A2(n459), .ZN(n458) );
  AND2_X1 U393 ( .A1(n372), .A2(KEYINPUT91), .ZN(n459) );
  OR2_X1 U394 ( .A1(n663), .A2(n462), .ZN(n461) );
  XNOR2_X1 U395 ( .A(n367), .B(n770), .ZN(n548) );
  INV_X1 U396 ( .A(G237), .ZN(n531) );
  NAND2_X1 U397 ( .A1(n392), .A2(KEYINPUT30), .ZN(n391) );
  OR2_X1 U398 ( .A1(n688), .A2(G902), .ZN(n477) );
  NAND2_X1 U399 ( .A1(G472), .A2(G902), .ZN(n437) );
  NAND2_X1 U400 ( .A1(n480), .A2(n436), .ZN(n435) );
  AND2_X1 U401 ( .A1(n626), .A2(n447), .ZN(n444) );
  OR2_X1 U402 ( .A1(n626), .A2(n447), .ZN(n441) );
  NOR2_X1 U403 ( .A1(n789), .A2(n788), .ZN(n402) );
  NAND2_X1 U404 ( .A1(n651), .A2(n463), .ZN(n462) );
  INV_X1 U405 ( .A(n550), .ZN(n463) );
  NAND2_X1 U406 ( .A1(n450), .A2(n464), .ZN(n372) );
  NAND2_X1 U407 ( .A1(n652), .A2(n550), .ZN(n464) );
  INV_X1 U408 ( .A(KEYINPUT103), .ZN(n409) );
  XNOR2_X1 U409 ( .A(n621), .B(KEYINPUT28), .ZN(n371) );
  AND2_X1 U410 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U411 ( .A1(n432), .A2(n409), .ZN(n407) );
  XNOR2_X1 U412 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X1 U413 ( .A(n479), .B(G137), .ZN(n395) );
  XNOR2_X1 U414 ( .A(n539), .B(n348), .ZN(n396) );
  XNOR2_X1 U415 ( .A(G110), .B(G107), .ZN(n768) );
  XNOR2_X1 U416 ( .A(n381), .B(n380), .ZN(n491) );
  XNOR2_X1 U417 ( .A(KEYINPUT78), .B(KEYINPUT85), .ZN(n381) );
  XNOR2_X1 U418 ( .A(G119), .B(KEYINPUT98), .ZN(n380) );
  XNOR2_X1 U419 ( .A(G128), .B(G110), .ZN(n487) );
  XNOR2_X1 U420 ( .A(n425), .B(KEYINPUT23), .ZN(n424) );
  INV_X1 U421 ( .A(KEYINPUT24), .ZN(n425) );
  INV_X1 U422 ( .A(KEYINPUT97), .ZN(n418) );
  XNOR2_X1 U423 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n489) );
  XOR2_X1 U424 ( .A(G131), .B(KEYINPUT70), .Z(n514) );
  XNOR2_X1 U425 ( .A(G104), .B(KEYINPUT79), .ZN(n474) );
  XNOR2_X1 U426 ( .A(n473), .B(KEYINPUT71), .ZN(n494) );
  INV_X1 U427 ( .A(KEYINPUT41), .ZN(n428) );
  NOR2_X1 U428 ( .A1(n718), .A2(n721), .ZN(n637) );
  NAND2_X1 U429 ( .A1(n461), .A2(n413), .ZN(n553) );
  NAND2_X1 U430 ( .A1(n390), .A2(n386), .ZN(n641) );
  AND2_X1 U431 ( .A1(n388), .A2(n366), .ZN(n386) );
  NAND2_X1 U432 ( .A1(n371), .A2(n622), .ZN(n636) );
  INV_X1 U433 ( .A(n595), .ZN(n622) );
  INV_X1 U434 ( .A(n624), .ZN(n370) );
  AND2_X1 U435 ( .A1(n371), .A2(n369), .ZN(n368) );
  NAND2_X1 U436 ( .A1(KEYINPUT47), .A2(n627), .ZN(n626) );
  NOR2_X1 U437 ( .A1(G953), .A2(G237), .ZN(n505) );
  AND2_X1 U438 ( .A1(n445), .A2(n443), .ZN(n442) );
  INV_X1 U439 ( .A(n761), .ZN(n439) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n481) );
  XNOR2_X1 U441 ( .A(G902), .B(KEYINPUT94), .ZN(n496) );
  INV_X1 U442 ( .A(KEYINPUT4), .ZN(n361) );
  XNOR2_X1 U443 ( .A(KEYINPUT70), .B(G131), .ZN(n471) );
  INV_X1 U444 ( .A(KEYINPUT48), .ZN(n415) );
  NOR2_X1 U445 ( .A1(n709), .A2(n412), .ZN(n710) );
  NAND2_X1 U446 ( .A1(n452), .A2(n451), .ZN(n460) );
  NAND2_X1 U447 ( .A1(n552), .A2(KEYINPUT91), .ZN(n451) );
  OR2_X1 U448 ( .A1(n663), .A2(n453), .ZN(n452) );
  NOR2_X1 U449 ( .A1(n615), .A2(n568), .ZN(n503) );
  NOR2_X1 U450 ( .A1(n715), .A2(n422), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n595), .B(n478), .ZN(n699) );
  XOR2_X1 U452 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n520) );
  XNOR2_X1 U453 ( .A(G134), .B(G122), .ZN(n519) );
  XOR2_X1 U454 ( .A(G107), .B(G116), .Z(n522) );
  INV_X1 U455 ( .A(KEYINPUT40), .ZN(n404) );
  NAND2_X1 U456 ( .A1(n643), .A2(n404), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n517), .B(n423), .ZN(n592) );
  XNOR2_X1 U458 ( .A(n518), .B(G475), .ZN(n423) );
  INV_X1 U459 ( .A(KEYINPUT6), .ZN(n411) );
  BUF_X1 U460 ( .A(n699), .Z(n393) );
  XNOR2_X1 U461 ( .A(n488), .B(n418), .ZN(n417) );
  XNOR2_X1 U462 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U463 ( .A(n475), .B(n365), .ZN(n364) );
  XNOR2_X1 U464 ( .A(n494), .B(n346), .ZN(n365) );
  NAND2_X1 U465 ( .A1(n384), .A2(KEYINPUT2), .ZN(n655) );
  XNOR2_X1 U466 ( .A(n403), .B(n639), .ZN(n788) );
  NOR2_X1 U467 ( .A1(n641), .A2(n553), .ZN(n431) );
  XOR2_X1 U468 ( .A(n643), .B(KEYINPUT106), .Z(n755) );
  AND2_X1 U469 ( .A1(n407), .A2(n405), .ZN(n345) );
  XOR2_X1 U470 ( .A(n474), .B(KEYINPUT80), .Z(n346) );
  XOR2_X1 U471 ( .A(n576), .B(KEYINPUT105), .Z(n347) );
  XNOR2_X1 U472 ( .A(KEYINPUT77), .B(KEYINPUT5), .ZN(n348) );
  AND2_X1 U473 ( .A1(n567), .A2(n632), .ZN(n349) );
  AND2_X1 U474 ( .A1(n565), .A2(n564), .ZN(n350) );
  OR2_X1 U475 ( .A1(n627), .A2(KEYINPUT47), .ZN(n351) );
  AND2_X1 U476 ( .A1(n698), .A2(n622), .ZN(n352) );
  AND2_X1 U477 ( .A1(n650), .A2(n649), .ZN(n353) );
  OR2_X1 U478 ( .A1(n643), .A2(n404), .ZN(n354) );
  INV_X1 U479 ( .A(G902), .ZN(n436) );
  OR2_X1 U480 ( .A1(n615), .A2(n387), .ZN(n355) );
  XOR2_X1 U481 ( .A(KEYINPUT81), .B(KEYINPUT32), .Z(n356) );
  XOR2_X1 U482 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n357) );
  NOR2_X1 U483 ( .A1(n636), .A2(n624), .ZN(n748) );
  INV_X1 U484 ( .A(KEYINPUT30), .ZN(n422) );
  OR2_X1 U485 ( .A1(n651), .A2(KEYINPUT87), .ZN(n358) );
  INV_X1 U486 ( .A(KEYINPUT84), .ZN(n447) );
  NAND2_X1 U487 ( .A1(n652), .A2(KEYINPUT2), .ZN(n359) );
  BUF_X1 U488 ( .A(n780), .Z(n427) );
  NOR2_X1 U489 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U490 ( .A1(n429), .A2(n375), .ZN(n374) );
  NOR2_X1 U491 ( .A1(n653), .A2(n358), .ZN(n375) );
  BUF_X1 U492 ( .A(n677), .Z(n685) );
  XNOR2_X2 U493 ( .A(n360), .B(G101), .ZN(n367) );
  XNOR2_X1 U494 ( .A(n360), .B(KEYINPUT125), .ZN(n776) );
  XNOR2_X2 U495 ( .A(n521), .B(n361), .ZN(n360) );
  XNOR2_X1 U496 ( .A(n364), .B(n362), .ZN(n688) );
  XNOR2_X1 U497 ( .A(n394), .B(n362), .ZN(n670) );
  NAND2_X1 U498 ( .A1(n363), .A2(n373), .ZN(n426) );
  XNOR2_X1 U499 ( .A(n363), .B(G119), .ZN(G21) );
  XNOR2_X2 U500 ( .A(n468), .B(n356), .ZN(n363) );
  NAND2_X1 U501 ( .A1(n413), .A2(n456), .ZN(n455) );
  NOR2_X1 U502 ( .A1(n595), .A2(n355), .ZN(n366) );
  NAND2_X1 U503 ( .A1(n370), .A2(n368), .ZN(n627) );
  AND2_X1 U504 ( .A1(n625), .A2(n622), .ZN(n369) );
  INV_X1 U505 ( .A(n372), .ZN(n413) );
  XNOR2_X1 U506 ( .A(n373), .B(G110), .ZN(G12) );
  XNOR2_X2 U507 ( .A(n469), .B(KEYINPUT104), .ZN(n373) );
  NAND2_X1 U508 ( .A1(n376), .A2(n374), .ZN(n383) );
  NAND2_X1 U509 ( .A1(n378), .A2(n377), .ZN(n376) );
  NOR2_X2 U510 ( .A1(n780), .A2(n430), .ZN(n377) );
  NAND2_X1 U511 ( .A1(n379), .A2(n652), .ZN(n378) );
  INV_X1 U512 ( .A(n653), .ZN(n379) );
  XNOR2_X2 U513 ( .A(n614), .B(n613), .ZN(n653) );
  XNOR2_X2 U514 ( .A(n385), .B(KEYINPUT88), .ZN(n780) );
  NAND2_X1 U515 ( .A1(n382), .A2(n359), .ZN(n466) );
  XNOR2_X1 U516 ( .A(n383), .B(n467), .ZN(n382) );
  INV_X1 U517 ( .A(n385), .ZN(n384) );
  NAND2_X1 U518 ( .A1(n619), .A2(n389), .ZN(n388) );
  AND2_X1 U519 ( .A1(n715), .A2(n422), .ZN(n389) );
  INV_X1 U520 ( .A(n619), .ZN(n392) );
  XNOR2_X2 U521 ( .A(n416), .B(n569), .ZN(n698) );
  OR2_X1 U522 ( .A1(n648), .A2(n354), .ZN(n398) );
  NAND2_X1 U523 ( .A1(n648), .A2(n404), .ZN(n401) );
  XNOR2_X1 U524 ( .A(n402), .B(n470), .ZN(n644) );
  NAND2_X1 U525 ( .A1(n732), .A2(n638), .ZN(n403) );
  NAND2_X1 U526 ( .A1(n433), .A2(n409), .ZN(n405) );
  NAND2_X1 U527 ( .A1(n408), .A2(n410), .ZN(n406) );
  NOR2_X1 U528 ( .A1(n432), .A2(n433), .ZN(n596) );
  NOR2_X1 U529 ( .A1(n433), .A2(n409), .ZN(n408) );
  INV_X1 U530 ( .A(n432), .ZN(n410) );
  XNOR2_X1 U531 ( .A(n596), .B(n411), .ZN(n600) );
  INV_X1 U532 ( .A(n596), .ZN(n412) );
  NAND2_X1 U533 ( .A1(n568), .A2(n702), .ZN(n416) );
  XNOR2_X1 U534 ( .A(n493), .B(n417), .ZN(n495) );
  XNOR2_X1 U535 ( .A(n628), .B(KEYINPUT19), .ZN(n623) );
  NAND2_X1 U536 ( .A1(n419), .A2(n585), .ZN(n420) );
  NAND2_X1 U537 ( .A1(n581), .A2(KEYINPUT66), .ZN(n419) );
  NOR2_X2 U538 ( .A1(n678), .A2(G902), .ZN(n500) );
  NAND2_X1 U539 ( .A1(n420), .A2(n589), .ZN(n612) );
  NOR2_X1 U540 ( .A1(n440), .A2(n439), .ZN(n438) );
  XNOR2_X1 U541 ( .A(n424), .B(n487), .ZN(n488) );
  NAND2_X1 U542 ( .A1(n442), .A2(n438), .ZN(n635) );
  NAND2_X1 U543 ( .A1(n351), .A2(n441), .ZN(n440) );
  XNOR2_X2 U544 ( .A(n563), .B(n562), .ZN(n603) );
  XNOR2_X2 U545 ( .A(n426), .B(n580), .ZN(n608) );
  XNOR2_X2 U546 ( .A(n578), .B(n577), .ZN(n590) );
  NOR2_X1 U547 ( .A1(n427), .A2(n654), .ZN(n694) );
  INV_X1 U548 ( .A(n780), .ZN(n429) );
  INV_X1 U549 ( .A(KEYINPUT87), .ZN(n430) );
  XNOR2_X1 U550 ( .A(n431), .B(n616), .ZN(n617) );
  NOR2_X1 U551 ( .A1(n670), .A2(n435), .ZN(n432) );
  NAND2_X1 U552 ( .A1(n670), .A2(G472), .ZN(n434) );
  NAND2_X1 U553 ( .A1(n752), .A2(n444), .ZN(n443) );
  NAND2_X1 U554 ( .A1(n446), .A2(KEYINPUT84), .ZN(n445) );
  INV_X1 U555 ( .A(n752), .ZN(n446) );
  XNOR2_X2 U556 ( .A(n449), .B(n448), .ZN(n539) );
  XNOR2_X2 U557 ( .A(KEYINPUT3), .B(G119), .ZN(n448) );
  XNOR2_X2 U558 ( .A(G116), .B(G113), .ZN(n449) );
  NAND2_X1 U559 ( .A1(n663), .A2(n550), .ZN(n450) );
  NAND2_X1 U560 ( .A1(n454), .A2(KEYINPUT91), .ZN(n453) );
  INV_X1 U561 ( .A(n462), .ZN(n454) );
  NAND2_X1 U562 ( .A1(n458), .A2(n455), .ZN(n628) );
  NOR2_X1 U563 ( .A1(n552), .A2(KEYINPUT91), .ZN(n457) );
  AND2_X2 U564 ( .A1(n466), .A2(n465), .ZN(n677) );
  INV_X1 U565 ( .A(n696), .ZN(n465) );
  INV_X1 U566 ( .A(KEYINPUT86), .ZN(n467) );
  NAND2_X1 U567 ( .A1(n603), .A2(n349), .ZN(n468) );
  NAND2_X1 U568 ( .A1(n603), .A2(n350), .ZN(n469) );
  XNOR2_X1 U569 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n470) );
  INV_X1 U570 ( .A(KEYINPUT72), .ZN(n634) );
  XNOR2_X1 U571 ( .A(n635), .B(n634), .ZN(n645) );
  INV_X1 U572 ( .A(G472), .ZN(n480) );
  BUF_X1 U573 ( .A(n521), .Z(n523) );
  BUF_X1 U574 ( .A(n623), .Z(n624) );
  INV_X1 U575 ( .A(KEYINPUT109), .ZN(n616) );
  XNOR2_X2 U576 ( .A(G143), .B(G128), .ZN(n521) );
  XNOR2_X1 U577 ( .A(n768), .B(KEYINPUT73), .ZN(n545) );
  INV_X2 U578 ( .A(G953), .ZN(n736) );
  NAND2_X1 U579 ( .A1(n736), .A2(G227), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n545), .B(n472), .ZN(n475) );
  XNOR2_X1 U581 ( .A(G137), .B(G140), .ZN(n473) );
  INV_X1 U582 ( .A(G469), .ZN(n476) );
  XNOR2_X1 U583 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n478) );
  NAND2_X1 U584 ( .A1(n505), .A2(G210), .ZN(n479) );
  XOR2_X1 U585 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n482) );
  XOR2_X1 U586 ( .A(n482), .B(n481), .Z(n485) );
  NAND2_X1 U587 ( .A1(n485), .A2(G902), .ZN(n554) );
  NOR2_X1 U588 ( .A1(n554), .A2(n736), .ZN(n483) );
  XNOR2_X1 U589 ( .A(n483), .B(KEYINPUT107), .ZN(n484) );
  NOR2_X1 U590 ( .A1(G900), .A2(n484), .ZN(n486) );
  NAND2_X1 U591 ( .A1(G952), .A2(n485), .ZN(n728) );
  NOR2_X1 U592 ( .A1(n728), .A2(G953), .ZN(n556) );
  NOR2_X1 U593 ( .A1(n486), .A2(n556), .ZN(n615) );
  NAND2_X1 U594 ( .A1(n736), .A2(G234), .ZN(n490) );
  XNOR2_X1 U595 ( .A(n490), .B(n489), .ZN(n526) );
  NAND2_X1 U596 ( .A1(n526), .A2(G221), .ZN(n492) );
  XOR2_X1 U597 ( .A(KEYINPUT10), .B(n541), .Z(n504) );
  XNOR2_X1 U598 ( .A(n494), .B(n504), .ZN(n778) );
  XNOR2_X1 U599 ( .A(n495), .B(n778), .ZN(n678) );
  XNOR2_X1 U600 ( .A(n496), .B(KEYINPUT15), .ZN(n651) );
  NAND2_X1 U601 ( .A1(G234), .A2(n651), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n497), .B(KEYINPUT20), .ZN(n501) );
  NAND2_X1 U603 ( .A1(n501), .A2(G217), .ZN(n498) );
  XNOR2_X2 U604 ( .A(n500), .B(n499), .ZN(n568) );
  AND2_X1 U605 ( .A1(n501), .A2(G221), .ZN(n502) );
  XNOR2_X1 U606 ( .A(n502), .B(KEYINPUT21), .ZN(n702) );
  NAND2_X1 U607 ( .A1(n503), .A2(n702), .ZN(n618) );
  NOR2_X1 U608 ( .A1(n600), .A2(n618), .ZN(n530) );
  XNOR2_X1 U609 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n518) );
  INV_X1 U610 ( .A(n504), .ZN(n513) );
  XOR2_X1 U611 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n507) );
  NAND2_X1 U612 ( .A1(G214), .A2(n505), .ZN(n506) );
  XNOR2_X1 U613 ( .A(n507), .B(n506), .ZN(n511) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(G140), .Z(n509) );
  XNOR2_X1 U615 ( .A(G113), .B(G143), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U618 ( .A(n513), .B(n512), .ZN(n516) );
  XNOR2_X2 U619 ( .A(G122), .B(G104), .ZN(n537) );
  XOR2_X1 U620 ( .A(n537), .B(n514), .Z(n515) );
  XNOR2_X1 U621 ( .A(n516), .B(n515), .ZN(n656) );
  NOR2_X1 U622 ( .A1(G902), .A2(n656), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n520), .B(n519), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U625 ( .A(n525), .B(n524), .ZN(n528) );
  NAND2_X1 U626 ( .A1(n526), .A2(G217), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n528), .B(n527), .ZN(n682) );
  NOR2_X1 U628 ( .A1(G902), .A2(n682), .ZN(n529) );
  XNOR2_X1 U629 ( .A(G478), .B(n529), .ZN(n591) );
  NAND2_X1 U630 ( .A1(n592), .A2(n591), .ZN(n643) );
  NAND2_X1 U631 ( .A1(n530), .A2(n755), .ZN(n630) );
  INV_X1 U632 ( .A(n630), .ZN(n532) );
  NAND2_X1 U633 ( .A1(n436), .A2(n531), .ZN(n549) );
  NAND2_X1 U634 ( .A1(n549), .A2(G214), .ZN(n715) );
  NAND2_X1 U635 ( .A1(n532), .A2(n715), .ZN(n533) );
  NOR2_X1 U636 ( .A1(n393), .A2(n533), .ZN(n534) );
  XOR2_X1 U637 ( .A(KEYINPUT43), .B(n534), .Z(n535) );
  XNOR2_X1 U638 ( .A(n535), .B(KEYINPUT108), .ZN(n551) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n536) );
  XNOR2_X1 U640 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U641 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n541), .B(n540), .ZN(n544) );
  NAND2_X1 U643 ( .A1(n736), .A2(G224), .ZN(n542) );
  XNOR2_X1 U644 ( .A(n542), .B(KEYINPUT95), .ZN(n543) );
  XNOR2_X1 U645 ( .A(n544), .B(n543), .ZN(n546) );
  XNOR2_X1 U646 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U647 ( .A1(n549), .A2(G210), .ZN(n550) );
  NAND2_X1 U648 ( .A1(n551), .A2(n553), .ZN(n649) );
  XNOR2_X1 U649 ( .A(n649), .B(G140), .ZN(G42) );
  INV_X1 U650 ( .A(n715), .ZN(n552) );
  XOR2_X1 U651 ( .A(G898), .B(KEYINPUT96), .Z(n765) );
  NAND2_X1 U652 ( .A1(G953), .A2(n765), .ZN(n771) );
  NOR2_X1 U653 ( .A1(n554), .A2(n771), .ZN(n555) );
  NOR2_X1 U654 ( .A1(n556), .A2(n555), .ZN(n557) );
  INV_X1 U655 ( .A(n591), .ZN(n575) );
  NOR2_X1 U656 ( .A1(n592), .A2(n575), .ZN(n559) );
  XNOR2_X1 U657 ( .A(n559), .B(KEYINPUT101), .ZN(n718) );
  INV_X1 U658 ( .A(n702), .ZN(n560) );
  NOR2_X1 U659 ( .A1(n718), .A2(n560), .ZN(n561) );
  INV_X1 U660 ( .A(KEYINPUT22), .ZN(n562) );
  NOR2_X1 U661 ( .A1(n619), .A2(n568), .ZN(n565) );
  INV_X1 U662 ( .A(n393), .ZN(n564) );
  XNOR2_X1 U663 ( .A(n568), .B(KEYINPUT102), .ZN(n703) );
  INV_X1 U664 ( .A(n703), .ZN(n566) );
  AND2_X1 U665 ( .A1(n600), .A2(n566), .ZN(n567) );
  XNOR2_X1 U666 ( .A(n393), .B(KEYINPUT92), .ZN(n632) );
  INV_X1 U667 ( .A(KEYINPUT68), .ZN(n569) );
  NAND2_X1 U668 ( .A1(n698), .A2(n699), .ZN(n593) );
  INV_X1 U669 ( .A(KEYINPUT33), .ZN(n570) );
  XNOR2_X1 U670 ( .A(n571), .B(n570), .ZN(n731) );
  NAND2_X1 U671 ( .A1(n731), .A2(n573), .ZN(n574) );
  AND2_X1 U672 ( .A1(n592), .A2(n575), .ZN(n576) );
  INV_X1 U673 ( .A(KEYINPUT35), .ZN(n577) );
  XOR2_X1 U674 ( .A(G122), .B(KEYINPUT127), .Z(n579) );
  XNOR2_X1 U675 ( .A(n590), .B(n579), .ZN(G24) );
  INV_X1 U676 ( .A(KEYINPUT90), .ZN(n580) );
  INV_X1 U677 ( .A(n608), .ZN(n581) );
  INV_X1 U678 ( .A(n590), .ZN(n583) );
  INV_X1 U679 ( .A(KEYINPUT89), .ZN(n582) );
  NAND2_X1 U680 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U681 ( .A1(n584), .A2(KEYINPUT44), .ZN(n585) );
  NAND2_X1 U682 ( .A1(n608), .A2(n590), .ZN(n588) );
  NOR2_X1 U683 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n586) );
  AND2_X1 U684 ( .A1(n586), .A2(KEYINPUT66), .ZN(n587) );
  NAND2_X1 U685 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X1 U686 ( .A1(n590), .A2(KEYINPUT89), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n592), .A2(n591), .ZN(n757) );
  INV_X1 U688 ( .A(n757), .ZN(n647) );
  NAND2_X1 U689 ( .A1(n643), .A2(n647), .ZN(n625) );
  INV_X1 U690 ( .A(n625), .ZN(n720) );
  NOR2_X1 U691 ( .A1(n596), .A2(n593), .ZN(n711) );
  NAND2_X1 U692 ( .A1(n573), .A2(n711), .ZN(n594) );
  XNOR2_X1 U693 ( .A(n594), .B(KEYINPUT31), .ZN(n758) );
  INV_X1 U694 ( .A(n573), .ZN(n598) );
  NAND2_X1 U695 ( .A1(n352), .A2(n596), .ZN(n597) );
  NOR2_X1 U696 ( .A1(n598), .A2(n597), .ZN(n744) );
  NOR2_X1 U697 ( .A1(n758), .A2(n744), .ZN(n599) );
  NOR2_X1 U698 ( .A1(n720), .A2(n599), .ZN(n604) );
  NAND2_X1 U699 ( .A1(n600), .A2(n703), .ZN(n601) );
  NOR2_X1 U700 ( .A1(n601), .A2(n393), .ZN(n602) );
  AND2_X1 U701 ( .A1(n603), .A2(n602), .ZN(n741) );
  OR2_X1 U702 ( .A1(n604), .A2(n741), .ZN(n605) );
  NOR2_X1 U703 ( .A1(n606), .A2(n605), .ZN(n610) );
  INV_X1 U704 ( .A(KEYINPUT66), .ZN(n607) );
  NAND2_X1 U705 ( .A1(n608), .A2(n607), .ZN(n609) );
  AND2_X1 U706 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U707 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X1 U708 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n613) );
  NAND2_X1 U709 ( .A1(n617), .A2(n347), .ZN(n752) );
  INV_X1 U710 ( .A(n618), .ZN(n620) );
  INV_X1 U711 ( .A(n628), .ZN(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U713 ( .A(n631), .B(KEYINPUT36), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n761) );
  XOR2_X1 U715 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n639) );
  INV_X1 U716 ( .A(n636), .ZN(n638) );
  XOR2_X1 U717 ( .A(KEYINPUT38), .B(n553), .Z(n640) );
  INV_X1 U718 ( .A(n640), .ZN(n716) );
  NAND2_X1 U719 ( .A1(n716), .A2(n715), .ZN(n721) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT39), .ZN(n648) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n762) );
  INV_X1 U723 ( .A(n762), .ZN(n650) );
  BUF_X1 U724 ( .A(n653), .Z(n654) );
  NOR2_X1 U725 ( .A1(n654), .A2(n655), .ZN(n696) );
  NAND2_X1 U726 ( .A1(n677), .A2(G475), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT59), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(n660) );
  INV_X1 U729 ( .A(G952), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n659), .A2(G953), .ZN(n680) );
  NAND2_X1 U731 ( .A1(n660), .A2(n680), .ZN(n662) );
  XNOR2_X1 U732 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(G60) );
  NAND2_X1 U734 ( .A1(n677), .A2(G210), .ZN(n666) );
  XNOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n663), .B(n664), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n667), .A2(n680), .ZN(n669) );
  XNOR2_X1 U739 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(G51) );
  NAND2_X1 U741 ( .A1(n677), .A2(G472), .ZN(n673) );
  XNOR2_X1 U742 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n670), .B(n671), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n674), .A2(n680), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT93), .B(KEYINPUT63), .Z(n675) );
  XNOR2_X1 U747 ( .A(n676), .B(n675), .ZN(G57) );
  NAND2_X1 U748 ( .A1(n685), .A2(G217), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n678), .B(n679), .ZN(n681) );
  INV_X1 U750 ( .A(n680), .ZN(n691) );
  NOR2_X1 U751 ( .A1(n681), .A2(n691), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n685), .A2(G478), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n684), .A2(n691), .ZN(G63) );
  NAND2_X1 U755 ( .A1(n685), .A2(G469), .ZN(n690) );
  XOR2_X1 U756 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT58), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U759 ( .A(n690), .B(n689), .ZN(n692) );
  NOR2_X1 U760 ( .A1(n692), .A2(n691), .ZN(G54) );
  XOR2_X1 U761 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n693) );
  NOR2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U763 ( .A(n695), .B(KEYINPUT82), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n739) );
  NOR2_X1 U765 ( .A1(n393), .A2(n698), .ZN(n701) );
  XNOR2_X1 U766 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n701), .B(n700), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n705) );
  XNOR2_X1 U769 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n704) );
  XNOR2_X1 U770 ( .A(n705), .B(n704), .ZN(n706) );
  XOR2_X1 U771 ( .A(KEYINPUT116), .B(n706), .Z(n707) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U774 ( .A(n712), .B(KEYINPUT118), .ZN(n713) );
  XNOR2_X1 U775 ( .A(n713), .B(KEYINPUT51), .ZN(n714) );
  NAND2_X1 U776 ( .A1(n732), .A2(n714), .ZN(n726) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U778 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U779 ( .A(n719), .B(KEYINPUT119), .ZN(n723) );
  OR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U781 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U782 ( .A1(n731), .A2(n724), .ZN(n725) );
  NAND2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U784 ( .A(KEYINPUT52), .B(n727), .ZN(n730) );
  INV_X1 U785 ( .A(n728), .ZN(n729) );
  NAND2_X1 U786 ( .A1(n730), .A2(n729), .ZN(n734) );
  NAND2_X1 U787 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U789 ( .A(KEYINPUT120), .B(n735), .Z(n737) );
  NAND2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U793 ( .A(G101), .B(n741), .Z(G3) );
  NAND2_X1 U794 ( .A1(n755), .A2(n744), .ZN(n742) );
  XNOR2_X1 U795 ( .A(n742), .B(KEYINPUT112), .ZN(n743) );
  XNOR2_X1 U796 ( .A(G104), .B(n743), .ZN(G6) );
  XOR2_X1 U797 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n746) );
  NAND2_X1 U798 ( .A1(n744), .A2(n757), .ZN(n745) );
  XNOR2_X1 U799 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U800 ( .A(G107), .B(n747), .ZN(G9) );
  XOR2_X1 U801 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n750) );
  NAND2_X1 U802 ( .A1(n748), .A2(n757), .ZN(n749) );
  XNOR2_X1 U803 ( .A(n750), .B(n749), .ZN(n751) );
  XOR2_X1 U804 ( .A(G128), .B(n751), .Z(G30) );
  XNOR2_X1 U805 ( .A(n752), .B(G143), .ZN(G45) );
  NAND2_X1 U806 ( .A1(n748), .A2(n755), .ZN(n753) );
  XNOR2_X1 U807 ( .A(n753), .B(KEYINPUT114), .ZN(n754) );
  XNOR2_X1 U808 ( .A(G146), .B(n754), .ZN(G48) );
  NAND2_X1 U809 ( .A1(n755), .A2(n758), .ZN(n756) );
  XNOR2_X1 U810 ( .A(n756), .B(G113), .ZN(G15) );
  NAND2_X1 U811 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n759), .B(G116), .ZN(G18) );
  XOR2_X1 U813 ( .A(G125), .B(KEYINPUT37), .Z(n760) );
  XNOR2_X1 U814 ( .A(n761), .B(n760), .ZN(G27) );
  XOR2_X1 U815 ( .A(G134), .B(n762), .Z(G36) );
  NOR2_X1 U816 ( .A1(n654), .A2(G953), .ZN(n767) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n763) );
  XOR2_X1 U818 ( .A(KEYINPUT61), .B(n763), .Z(n764) );
  NOR2_X1 U819 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U820 ( .A1(n767), .A2(n766), .ZN(n774) );
  XNOR2_X1 U821 ( .A(n768), .B(G101), .ZN(n769) );
  XNOR2_X1 U822 ( .A(n770), .B(n769), .ZN(n772) );
  NAND2_X1 U823 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U824 ( .A(n774), .B(n773), .ZN(n775) );
  XNOR2_X1 U825 ( .A(KEYINPUT124), .B(n775), .ZN(G69) );
  XNOR2_X1 U826 ( .A(n777), .B(n776), .ZN(n779) );
  XNOR2_X1 U827 ( .A(n779), .B(n778), .ZN(n782) );
  XOR2_X1 U828 ( .A(n427), .B(n782), .Z(n781) );
  NOR2_X1 U829 ( .A1(G953), .A2(n781), .ZN(n786) );
  XNOR2_X1 U830 ( .A(G227), .B(n782), .ZN(n784) );
  NAND2_X1 U831 ( .A1(G900), .A2(G953), .ZN(n783) );
  NOR2_X1 U832 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U833 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U834 ( .A(KEYINPUT126), .B(n787), .ZN(G72) );
  XOR2_X1 U835 ( .A(G137), .B(n788), .Z(G39) );
  XOR2_X1 U836 ( .A(n789), .B(G131), .Z(G33) );
endmodule

