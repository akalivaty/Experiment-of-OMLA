//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  XOR2_X1   g000(.A(KEYINPUT26), .B(G101), .Z(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT29), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .A3(G143), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT0), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n205), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n203), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT65), .B1(new_n198), .B2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n201), .A3(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n206), .A3(new_n200), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n201), .A2(G143), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n210), .B2(new_n212), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT66), .A3(new_n206), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n209), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  INV_X1    g035(.A(G134), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G137), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(G137), .ZN(new_n224));
  INV_X1    g038(.A(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT11), .A3(G134), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G131), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n226), .A3(new_n229), .A4(new_n224), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n220), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n223), .A2(new_n226), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n229), .A4(new_n224), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n218), .A2(new_n240), .A3(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n203), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n224), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n222), .A2(G137), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n234), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT2), .B(G113), .Z(new_n252));
  XNOR2_X1  g066(.A(G116), .B(G119), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(KEYINPUT68), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(new_n252), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n262));
  INV_X1    g076(.A(new_n249), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n203), .A2(new_n207), .A3(new_n208), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n218), .A2(KEYINPUT66), .A3(new_n206), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT66), .B1(new_n218), .B2(new_n206), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n227), .A2(G131), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n237), .B2(new_n238), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n264), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n220), .A2(KEYINPUT69), .A3(new_n233), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n257), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n268), .A2(new_n270), .A3(new_n264), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT69), .B1(new_n220), .B2(new_n233), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n257), .B(new_n249), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n273), .B2(new_n257), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n275), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(new_n280), .A3(new_n257), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT74), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n274), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n262), .B1(new_n286), .B2(new_n259), .ZN(new_n287));
  INV_X1    g101(.A(new_n274), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n283), .A2(KEYINPUT74), .A3(new_n284), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT74), .B1(new_n283), .B2(new_n284), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n196), .B(new_n261), .C1(new_n287), .C2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT30), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n234), .A2(new_n295), .A3(new_n249), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n273), .B2(new_n295), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n256), .A2(new_n297), .B1(new_n283), .B2(new_n284), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n194), .B1(new_n298), .B2(new_n192), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n283), .A2(KEYINPUT28), .A3(new_n284), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n251), .A2(new_n257), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n259), .B2(new_n258), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n192), .B(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n299), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n297), .A2(new_n256), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n283), .A2(new_n284), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n310), .B2(new_n193), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT73), .B1(new_n311), .B2(new_n304), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n294), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G472), .B1(new_n293), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n303), .B1(new_n300), .B2(new_n302), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n309), .A3(new_n192), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT31), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT31), .A4(new_n192), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(G472), .A2(G902), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT32), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n316), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT31), .B1(new_n298), .B2(new_n192), .ZN(new_n326));
  AND4_X1   g140(.A1(KEYINPUT31), .A2(new_n308), .A3(new_n309), .A4(new_n192), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT32), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n322), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n314), .A2(new_n315), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G472), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n286), .A2(new_n262), .A3(new_n259), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT75), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n195), .B(new_n260), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n306), .B1(new_n299), .B2(new_n305), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n311), .A2(KEYINPUT73), .A3(new_n304), .ZN(new_n338));
  AOI21_X1  g152(.A(G902), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n333), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n324), .A2(new_n330), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n348), .A3(G140), .ZN(new_n349));
  INV_X1    g163(.A(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n344), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n348), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n353), .A2(KEYINPUT16), .A3(G140), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n201), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT78), .B(G125), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n344), .A3(new_n350), .ZN(new_n357));
  NOR2_X1   g171(.A1(G125), .A2(G140), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n356), .B2(G140), .ZN(new_n359));
  OAI211_X1 g173(.A(G146), .B(new_n357), .C1(new_n359), .C2(new_n344), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(KEYINPUT79), .A3(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(G119), .B(G128), .Z(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT77), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT24), .B(G110), .Z(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n352), .A2(new_n354), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G146), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n369), .A2(new_n205), .A3(G119), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n369), .B1(G119), .B2(new_n205), .ZN(new_n371));
  OAI22_X1  g185(.A1(new_n370), .A2(new_n371), .B1(G119), .B2(new_n205), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G110), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n361), .A2(new_n365), .A3(new_n368), .A4(new_n373), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT80), .B(G110), .Z(new_n375));
  OAI22_X1  g189(.A1(new_n363), .A2(new_n364), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(G125), .A2(G140), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n351), .A2(KEYINPUT81), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT81), .B1(new_n351), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n201), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n360), .A3(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n374), .A2(KEYINPUT82), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT82), .B1(new_n374), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(G221), .A3(G234), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT22), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(G137), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT83), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n374), .A2(new_n381), .A3(new_n388), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n391));
  INV_X1    g205(.A(new_n388), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n391), .B(new_n392), .C1(new_n382), .C2(new_n383), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n389), .A2(new_n294), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G217), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(G234), .B2(new_n294), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n399), .A2(G902), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G214), .B1(G237), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G107), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G104), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT3), .ZN(new_n412));
  INV_X1    g226(.A(G104), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G107), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n414), .B2(new_n412), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT86), .B(KEYINPUT3), .C1(new_n413), .C2(G107), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G101), .ZN(new_n420));
  INV_X1    g234(.A(G101), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n415), .A2(new_n417), .A3(new_n421), .A4(new_n418), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(KEYINPUT4), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n424), .A3(G101), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n256), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT88), .B(KEYINPUT5), .Z(new_n427));
  INV_X1    g241(.A(G116), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(G119), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n430), .A2(G113), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT68), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n253), .B(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n431), .B1(new_n433), .B2(new_n427), .ZN(new_n434));
  OAI21_X1  g248(.A(G101), .B1(new_n414), .B2(new_n411), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n422), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n437), .A3(new_n254), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(G110), .B(G122), .Z(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n440), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n426), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n245), .A2(new_n353), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n268), .B2(new_n353), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n385), .A2(G224), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n446), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n439), .A2(new_n450), .A3(new_n440), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT89), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n444), .A2(new_n449), .A3(new_n454), .A4(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n431), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n254), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n437), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n440), .B(KEYINPUT8), .Z(new_n461));
  NAND3_X1  g275(.A1(new_n434), .A2(new_n254), .A3(new_n436), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n446), .A2(KEYINPUT7), .A3(new_n448), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n443), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n446), .B1(KEYINPUT7), .B2(new_n448), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n456), .A2(new_n294), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n453), .B2(new_n455), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n469), .A3(new_n467), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n409), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n361), .A2(new_n368), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n188), .A2(G214), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n198), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n229), .A3(new_n476), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n475), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  XOR2_X1   g300(.A(G113), .B(G122), .Z(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT92), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(new_n413), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n359), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n380), .B1(new_n491), .B2(new_n201), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(KEYINPUT90), .A3(new_n476), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT18), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n493), .A2(new_n494), .A3(new_n229), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n229), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n477), .A2(new_n478), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(KEYINPUT90), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n492), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n486), .A2(new_n490), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n490), .B1(new_n486), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n294), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G475), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT19), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n378), .B2(new_n379), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n349), .A2(KEYINPUT19), .A3(new_n351), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n201), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n479), .A2(new_n484), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n360), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT91), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n499), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n489), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(G475), .B1(new_n515), .B2(new_n500), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n516), .A2(new_n517), .A3(new_n294), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n516), .B2(new_n294), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n504), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g334(.A(KEYINPUT9), .B(G234), .Z(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n522), .A2(new_n398), .A3(G953), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n524));
  NOR2_X1   g338(.A1(new_n205), .A2(G143), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT94), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n198), .A2(G128), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n524), .B2(new_n526), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n525), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G134), .ZN(new_n534));
  XNOR2_X1  g348(.A(G116), .B(G122), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G107), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n410), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n525), .A2(new_n528), .A3(G134), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT95), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT96), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n533), .A2(G134), .B1(new_n537), .B2(new_n538), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n541), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n525), .A2(new_n528), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n222), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n428), .A2(KEYINPUT14), .A3(G122), .ZN(new_n550));
  OAI211_X1 g364(.A(G107), .B(new_n550), .C1(new_n536), .C2(KEYINPUT14), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n538), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n523), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n552), .ZN(new_n554));
  INV_X1    g368(.A(new_n523), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n554), .B(new_n555), .C1(new_n543), .C2(new_n546), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n294), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(G478), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  OAI221_X1 g374(.A(new_n294), .B1(KEYINPUT15), .B2(new_n560), .C1(new_n553), .C2(new_n556), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n385), .A2(G952), .ZN(new_n563));
  NAND2_X1  g377(.A1(G234), .A2(G237), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT21), .B(G898), .Z(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(G902), .A3(G953), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n520), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G221), .B1(new_n522), .B2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(G110), .B(G140), .Z(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT85), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n385), .A2(G227), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g390(.A(new_n241), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n218), .B1(G128), .B2(new_n242), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n437), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n245), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n436), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n270), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT12), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT87), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n437), .A2(new_n584), .A3(KEYINPUT10), .A4(new_n245), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n422), .A2(KEYINPUT10), .A3(new_n435), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT87), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n579), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n423), .A2(new_n220), .A3(new_n425), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n270), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n576), .B1(new_n583), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n576), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n233), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G469), .B1(new_n597), .B2(G902), .ZN(new_n598));
  INV_X1    g412(.A(G469), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n582), .A2(KEYINPUT12), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n582), .A2(KEYINPUT12), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n594), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n595), .A2(new_n233), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n576), .B1(new_n603), .B2(new_n592), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n599), .B(new_n294), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n572), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n474), .A2(new_n570), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n343), .A2(new_n407), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  AND3_X1   g424(.A1(new_n472), .A2(new_n469), .A3(new_n467), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n469), .B1(new_n472), .B2(new_n467), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n568), .B(new_n408), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT33), .B1(new_n553), .B2(new_n556), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n542), .A2(KEYINPUT96), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n545), .B1(new_n544), .B2(new_n541), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n552), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n555), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n547), .A2(new_n552), .A3(new_n523), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n621), .A3(G478), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n560), .B(new_n294), .C1(new_n553), .C2(new_n556), .ZN(new_n623));
  NAND2_X1  g437(.A1(G478), .A2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT97), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n622), .A2(new_n627), .A3(new_n623), .A4(new_n624), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n520), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT98), .B1(new_n613), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n519), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n516), .A2(new_n517), .A3(new_n294), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n632), .A2(new_n633), .B1(G475), .B2(new_n503), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n626), .B2(new_n628), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n474), .A2(new_n635), .A3(new_n636), .A4(new_n568), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n321), .B2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n328), .A2(new_n322), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n606), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n406), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(new_n562), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n520), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(new_n650), .A3(new_n569), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n471), .A2(new_n473), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n408), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT99), .B1(new_n648), .B2(new_n568), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n643), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT100), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(G9));
  AND3_X1   g473(.A1(new_n652), .A2(new_n570), .A3(new_n408), .ZN(new_n660));
  INV_X1    g474(.A(new_n641), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n392), .A2(KEYINPUT36), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n384), .B(new_n662), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n404), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n401), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n660), .A2(new_n606), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n606), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n567), .A2(G900), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n565), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n648), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n343), .A2(new_n474), .A3(new_n671), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n673), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n606), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT40), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n394), .B(new_n395), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n681), .A2(new_n399), .B1(new_n404), .B2(new_n663), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n634), .A2(new_n647), .A3(new_n409), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n652), .B(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(new_n303), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n291), .A2(new_n686), .B1(new_n192), .B2(new_n298), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n331), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n680), .A2(new_n684), .A3(new_n685), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NAND2_X1  g505(.A1(new_n635), .A2(new_n673), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n474), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n692), .A2(new_n653), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n670), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n343), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  NOR2_X1   g514(.A1(new_n602), .A2(new_n604), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n571), .A3(new_n605), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n343), .A2(new_n638), .A3(new_n407), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND4_X1  g520(.A1(new_n343), .A2(new_n407), .A3(new_n655), .A4(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND3_X1  g522(.A1(new_n652), .A2(new_n703), .A3(new_n408), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n682), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n343), .A2(new_n570), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND2_X1  g526(.A1(new_n683), .A2(new_n652), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n261), .B1(new_n287), .B2(new_n292), .ZN(new_n716));
  OAI22_X1  g530(.A1(new_n716), .A2(new_n303), .B1(new_n326), .B2(new_n327), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n322), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(new_n639), .ZN(new_n719));
  INV_X1    g533(.A(new_n703), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n569), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n715), .A2(new_n719), .A3(new_n407), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT104), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(G122), .Z(G24));
  AND4_X1   g538(.A1(new_n639), .A2(new_n710), .A3(new_n718), .A4(new_n693), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n345), .ZN(G27));
  NAND3_X1  g540(.A1(new_n471), .A2(new_n408), .A3(new_n473), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n692), .A2(new_n642), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n315), .B1(new_n314), .B2(new_n331), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT76), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n407), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT105), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n406), .B1(new_n332), .B2(new_n342), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n728), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n732), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n331), .B(KEYINPUT106), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(new_n340), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n407), .A4(new_n728), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NOR3_X1   g556(.A1(new_n642), .A2(new_n674), .A3(new_n727), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n734), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n734), .A2(KEYINPUT107), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  AND3_X1   g563(.A1(new_n629), .A2(KEYINPUT43), .A3(new_n634), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT43), .B1(new_n629), .B2(new_n634), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n641), .B(new_n665), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n611), .A2(new_n612), .A3(new_n409), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n752), .B2(new_n753), .ZN(new_n756));
  INV_X1    g570(.A(new_n605), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n597), .A2(KEYINPUT45), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n593), .B2(new_n596), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(G469), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n571), .A3(new_n678), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n754), .A2(new_n756), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n225), .ZN(G39));
  AOI21_X1  g584(.A(KEYINPUT47), .B1(new_n767), .B2(new_n571), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n772), .B(new_n572), .C1(new_n765), .C2(new_n766), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n693), .B(new_n755), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n332), .A2(new_n342), .A3(new_n406), .ZN(new_n775));
  OR3_X1    g589(.A1(new_n774), .A2(KEYINPUT108), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT108), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n350), .ZN(G42));
  NOR2_X1   g593(.A1(new_n750), .A2(new_n751), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n755), .A2(new_n564), .A3(new_n563), .A4(new_n703), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n739), .A2(new_n407), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(KEYINPUT48), .A3(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n781), .A2(new_n406), .A3(new_n689), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n635), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n563), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n786), .A2(KEYINPUT48), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n780), .A2(new_n565), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n407), .A3(new_n719), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n709), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n790), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT115), .Z(new_n796));
  NAND3_X1  g610(.A1(new_n719), .A2(new_n693), .A3(new_n710), .ZN(new_n797));
  INV_X1    g611(.A(new_n673), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n665), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n715), .A2(new_n606), .A3(new_n689), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n676), .A2(new_n699), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n332), .A2(new_n342), .B1(new_n694), .B2(KEYINPUT102), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n725), .B1(new_n804), .B2(new_n698), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n676), .A4(new_n800), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT110), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n803), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n520), .A2(new_n562), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n471), .A2(new_n813), .A3(new_n408), .A4(new_n473), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n814), .B2(new_n798), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n755), .A2(KEYINPUT109), .A3(new_n813), .A4(new_n673), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n815), .B(new_n816), .C1(new_n729), .C2(new_n730), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n639), .A2(new_n718), .A3(new_n693), .A4(new_n755), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n670), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n630), .A2(new_n649), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n407), .A3(new_n661), .A4(new_n606), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n666), .B1(new_n822), .B2(new_n613), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n609), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n704), .A2(new_n707), .A3(new_n711), .A4(new_n722), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n748), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n737), .A2(new_n740), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n830), .A2(new_n807), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(KEYINPUT53), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n823), .B1(new_n734), .B2(new_n608), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n816), .A2(new_n815), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n332), .B2(new_n342), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n671), .B1(new_n837), .B2(new_n818), .ZN(new_n838));
  AND4_X1   g652(.A1(KEYINPUT107), .A2(new_n343), .A3(new_n407), .A4(new_n743), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT107), .B1(new_n734), .B2(new_n743), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n835), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n704), .A2(new_n707), .A3(new_n711), .A4(new_n722), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n807), .A3(KEYINPUT53), .A4(new_n741), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT53), .B1(new_n811), .B2(new_n830), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n796), .A2(new_n834), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n685), .A2(new_n408), .A3(new_n720), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT112), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(new_n793), .ZN(new_n854));
  OR2_X1    g668(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(KEYINPUT113), .B2(KEYINPUT50), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n702), .A2(new_n605), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n773), .B(new_n771), .C1(new_n572), .C2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n727), .A3(new_n793), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n780), .A2(new_n682), .A3(new_n781), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n629), .A2(new_n520), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n861), .A2(new_n719), .B1(new_n788), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n854), .B2(new_n855), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n857), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT51), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n851), .A2(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n629), .A2(new_n634), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT49), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n858), .A2(new_n869), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n685), .A2(new_n868), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n689), .A2(new_n406), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n571), .A3(new_n408), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n867), .A2(new_n874), .ZN(G75));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n830), .A2(new_n845), .A3(KEYINPUT53), .A4(new_n807), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n844), .A2(KEYINPUT111), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(G210), .B(G902), .C1(new_n879), .C2(new_n847), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n385), .A2(G952), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n876), .A3(new_n881), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n444), .A2(new_n451), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n449), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT55), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n887), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n880), .A2(new_n876), .A3(new_n881), .A4(new_n889), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n882), .B(new_n883), .C1(new_n888), .C2(new_n890), .ZN(G51));
  XOR2_X1   g705(.A(new_n762), .B(KEYINPUT57), .Z(new_n892));
  AOI21_X1  g706(.A(new_n849), .B1(new_n846), .B2(new_n848), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n879), .A2(new_n847), .A3(KEYINPUT54), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n701), .B(KEYINPUT117), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n294), .B1(new_n846), .B2(new_n848), .ZN(new_n898));
  INV_X1    g712(.A(new_n761), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n883), .B1(new_n897), .B2(new_n900), .ZN(G54));
  NAND3_X1  g715(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n500), .A3(new_n515), .ZN(new_n903));
  INV_X1    g717(.A(new_n883), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n515), .A2(new_n500), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .A4(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(G60));
  NAND2_X1  g721(.A1(new_n614), .A2(new_n621), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n850), .A2(new_n834), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n624), .B(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n910), .ZN(new_n912));
  INV_X1    g726(.A(new_n893), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n850), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n911), .A2(new_n914), .A3(new_n883), .ZN(G63));
  NAND2_X1  g729(.A1(new_n846), .A2(new_n848), .ZN(new_n916));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  AOI21_X1  g732(.A(new_n403), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n663), .B(new_n918), .C1(new_n879), .C2(new_n847), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n904), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  OR3_X1    g736(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n919), .B2(new_n921), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G66));
  NAND2_X1  g739(.A1(new_n827), .A2(new_n835), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n385), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n566), .A2(G224), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n927), .B(KEYINPUT118), .C1(new_n385), .C2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(KEYINPUT118), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n885), .B1(G898), .B2(new_n385), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT119), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n930), .B(new_n932), .ZN(G69));
  AND3_X1   g747(.A1(new_n676), .A2(new_n699), .A3(new_n797), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n690), .ZN(new_n935));
  NOR2_X1   g749(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n778), .A2(new_n769), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n679), .A2(new_n727), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n734), .A2(new_n821), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n937), .A2(new_n938), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n385), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n297), .B(KEYINPUT120), .Z(new_n944));
  AND2_X1   g758(.A1(new_n506), .A2(new_n507), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n944), .B(new_n945), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n767), .A2(new_n571), .A3(new_n678), .ZN(new_n949));
  AND4_X1   g763(.A1(new_n407), .A2(new_n739), .A3(new_n715), .A4(new_n949), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n950), .B(new_n769), .C1(new_n776), .C2(new_n777), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n741), .A2(new_n748), .A3(new_n934), .ZN(new_n952));
  AOI21_X1  g766(.A(G953), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n385), .A2(G900), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT122), .Z(new_n955));
  OAI21_X1  g769(.A(new_n946), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n958), .B(new_n946), .C1(new_n953), .C2(new_n955), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n948), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n385), .B1(G227), .B2(G900), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  INV_X1    g777(.A(new_n961), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n948), .A2(new_n964), .A3(new_n956), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n948), .A2(KEYINPUT123), .A3(new_n964), .A4(new_n956), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n960), .A2(new_n970), .A3(new_n961), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n963), .A2(new_n969), .A3(new_n971), .ZN(G72));
  XNOR2_X1  g786(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n333), .A2(new_n294), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n942), .B2(new_n926), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n298), .A2(new_n193), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n951), .A2(new_n952), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n975), .B1(new_n979), .B2(new_n926), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n310), .A2(new_n192), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n883), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n981), .ZN(new_n984));
  INV_X1    g798(.A(new_n977), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(new_n985), .A3(new_n975), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n983), .B1(new_n833), .B2(new_n987), .ZN(G57));
endmodule


