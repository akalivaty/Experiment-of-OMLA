//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n203), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n213), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n204), .A2(new_n205), .ZN(new_n230));
  INV_X1    g0030(.A(G50), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n211), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n216), .A2(new_n229), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT76), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n211), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n211), .A2(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n223), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n212), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n233), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n262), .A2(KEYINPUT11), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n212), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n211), .A3(G1), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n210), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G68), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(KEYINPUT11), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n203), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT12), .ZN(new_n274));
  AND4_X1   g0074(.A1(new_n263), .A2(new_n271), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT65), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT65), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G226), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G232), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n280), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G97), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  OAI211_X1 g0095(.A(G1), .B(G13), .C1(new_n254), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n296), .A3(G274), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n293), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n218), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n276), .B1(new_n292), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n296), .B1(new_n288), .B2(new_n289), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n302), .A2(KEYINPUT13), .A3(new_n299), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G179), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n301), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(KEYINPUT14), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT71), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT14), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n306), .B2(KEYINPUT70), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT70), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(G169), .C1(new_n301), .C2(new_n303), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  INV_X1    g0115(.A(new_n289), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n283), .B1(new_n281), .B2(new_n282), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(new_n287), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n276), .B(new_n300), .C1(new_n320), .C2(new_n296), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT13), .B1(new_n302), .B2(new_n299), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT14), .B1(new_n323), .B2(new_n312), .ZN(new_n324));
  AOI211_X1 g0124(.A(KEYINPUT70), .B(new_n315), .C1(new_n321), .C2(new_n322), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n324), .A2(KEYINPUT71), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n308), .B1(new_n314), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT71), .B1(new_n324), .B2(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n306), .A2(KEYINPUT70), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n330), .A2(new_n309), .A3(KEYINPUT14), .A4(new_n313), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(new_n308), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n275), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G226), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n297), .B1(new_n298), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G1698), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n280), .A2(G222), .A3(new_n338), .A4(new_n284), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n280), .A2(G223), .A3(G1698), .A4(new_n284), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n319), .C2(new_n223), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n341), .B2(new_n291), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT69), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  OR3_X1    g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT68), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n342), .A2(G190), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n270), .A2(G50), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT66), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n269), .A2(new_n351), .B1(new_n231), .B2(new_n266), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n211), .B1(new_n230), .B2(new_n231), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT8), .B(G58), .ZN(new_n354));
  INV_X1    g0154(.A(G150), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n354), .A2(new_n258), .B1(new_n355), .B2(new_n255), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n261), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n352), .A2(KEYINPUT9), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT9), .B1(new_n352), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n345), .A2(new_n347), .A3(new_n360), .A4(new_n348), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT10), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n349), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n349), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366));
  INV_X1    g0166(.A(new_n270), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n354), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n268), .B1(KEYINPUT75), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(KEYINPUT75), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n369), .A2(new_n370), .B1(new_n266), .B2(new_n354), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n282), .B1(new_n278), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n281), .A2(KEYINPUT74), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT7), .B(new_n211), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(G20), .B1(new_n280), .B2(new_n284), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G68), .ZN(new_n378));
  INV_X1    g0178(.A(G159), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n255), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G58), .A2(G68), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n204), .A2(new_n205), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n382), .B2(G20), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT16), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n278), .A2(new_n279), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT7), .B1(new_n385), .B2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n281), .A2(new_n282), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(new_n211), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(G68), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  AOI211_X1 g0192(.A(KEYINPUT73), .B(new_n380), .C1(new_n382), .C2(G20), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT16), .B(new_n390), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n261), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n371), .B1(new_n384), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(G223), .A2(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n336), .A2(G1698), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n385), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n296), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n297), .B1(new_n298), .B2(new_n286), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G169), .ZN(new_n404));
  INV_X1    g0204(.A(G179), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n366), .B1(new_n396), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n396), .A2(new_n366), .A3(new_n406), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n384), .A2(new_n395), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n401), .A2(new_n411), .A3(new_n402), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(G200), .B2(new_n403), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n371), .A4(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n371), .C1(new_n384), .C2(new_n395), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND4_X1   g0217(.A1(new_n408), .A2(new_n409), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n352), .A2(new_n357), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n342), .B2(G169), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n405), .B2(new_n342), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n304), .A2(G190), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n275), .B(new_n423), .C1(new_n344), .C2(new_n304), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n268), .A2(new_n223), .A3(new_n367), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n223), .B2(new_n266), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n258), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n354), .A2(new_n255), .B1(new_n211), .B2(new_n223), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(KEYINPUT67), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(KEYINPUT67), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n261), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n297), .B1(new_n298), .B2(new_n224), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n319), .A2(G232), .A3(new_n338), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n319), .A2(G238), .A3(G1698), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(new_n436), .C1(new_n225), .C2(new_n319), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n434), .B1(new_n437), .B2(new_n291), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n433), .B1(new_n438), .B2(G190), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n344), .B2(new_n438), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n405), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n433), .C1(G169), .C2(new_n438), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n424), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n365), .A2(new_n418), .A3(new_n422), .A4(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n253), .B1(new_n335), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n409), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n407), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n415), .B(KEYINPUT17), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n349), .A2(new_n362), .ZN(new_n450));
  INV_X1    g0250(.A(new_n361), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n349), .A2(new_n361), .A3(new_n362), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n422), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n275), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n333), .B1(new_n332), .B2(new_n308), .ZN(new_n457));
  AOI211_X1 g0257(.A(KEYINPUT72), .B(new_n307), .C1(new_n329), .C2(new_n331), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(new_n459), .A3(KEYINPUT76), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n445), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G257), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n338), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n385), .A2(new_n463), .B1(G33), .B2(G294), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n220), .A2(G1698), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT84), .B1(new_n385), .B2(new_n465), .ZN(new_n466));
  AND4_X1   g0266(.A1(KEYINPUT84), .A2(new_n465), .A3(new_n281), .A4(new_n282), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT5), .B(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n291), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n468), .A2(new_n291), .B1(G264), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n471), .A2(new_n296), .A3(G274), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G169), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(G179), .A3(new_n474), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT85), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n476), .B2(new_n477), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n219), .A2(KEYINPUT22), .A3(G20), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n280), .A2(new_n284), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n281), .A2(new_n282), .A3(new_n211), .A4(G87), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT22), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n486), .B2(KEYINPUT22), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT82), .B(new_n485), .C1(new_n488), .C2(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR3_X1    g0294(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(KEYINPUT83), .B1(KEYINPUT23), .B2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n495), .A2(KEYINPUT83), .B1(new_n498), .B2(G20), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n483), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  AOI211_X1 g0302(.A(KEYINPUT24), .B(new_n500), .C1(new_n492), .C2(new_n493), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n261), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n264), .B(new_n267), .C1(G1), .C2(new_n254), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT25), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n267), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n225), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n506), .A2(G107), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n482), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n475), .A2(new_n344), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(G190), .B2(new_n475), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n504), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G116), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n260), .A2(new_n233), .B1(G20), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT77), .B(G97), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G33), .ZN(new_n520));
  INV_X1    g0320(.A(G283), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n211), .B1(new_n254), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n518), .B(KEYINPUT20), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n267), .A2(G116), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n506), .B2(G116), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n471), .A2(new_n470), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n296), .ZN(new_n533));
  INV_X1    g0333(.A(G270), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n474), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n474), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G303), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n280), .B2(new_n284), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G257), .A2(G1698), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n338), .A2(G264), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n387), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n291), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT80), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(KEYINPUT80), .B(new_n291), .C1(new_n541), .C2(new_n544), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n539), .A2(G190), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n539), .A2(new_n548), .A3(new_n547), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n531), .B(new_n549), .C1(new_n550), .C2(new_n344), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(G179), .A3(new_n530), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n315), .B1(new_n527), .B2(new_n529), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n539), .A2(new_n548), .A3(new_n547), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n554), .A2(new_n555), .A3(new_n553), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n551), .B(new_n552), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n385), .A2(new_n211), .A3(G68), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n519), .B2(new_n258), .ZN(new_n561));
  XOR2_X1   g0361(.A(KEYINPUT77), .B(G97), .Z(new_n562));
  NOR3_X1   g0362(.A1(new_n562), .A2(G87), .A3(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(G20), .B1(new_n316), .B2(KEYINPUT19), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n559), .B(new_n561), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(new_n261), .B1(new_n266), .B2(new_n427), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G238), .A2(G1698), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n224), .B2(G1698), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n385), .A2(new_n568), .B1(G33), .B2(G116), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(new_n296), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n296), .B(G250), .C1(G1), .C2(new_n469), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n296), .A2(G274), .A3(new_n470), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(G190), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n506), .A2(G87), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n566), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n575), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n570), .A2(G179), .A3(new_n574), .ZN(new_n581));
  INV_X1    g0381(.A(new_n427), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n506), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n566), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n315), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n578), .A2(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n267), .A2(G97), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n506), .B2(G97), .ZN(new_n588));
  INV_X1    g0388(.A(G97), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n225), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n207), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n225), .A2(KEYINPUT6), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n591), .A2(KEYINPUT6), .B1(new_n519), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n256), .A2(G77), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(G107), .B2(new_n377), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n588), .B1(new_n597), .B2(new_n264), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n280), .A2(G250), .A3(G1698), .A4(new_n284), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n281), .A2(new_n282), .A3(G244), .A4(new_n338), .ZN(new_n600));
  XOR2_X1   g0400(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n601));
  AOI22_X1  g0401(.A1(new_n600), .A2(new_n601), .B1(G33), .B2(G283), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n280), .A2(new_n284), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n338), .A2(KEYINPUT4), .A3(G244), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n291), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n472), .A2(G257), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(new_n474), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n315), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(new_n405), .A3(new_n608), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n598), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(G200), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n377), .A2(G107), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n261), .B1(new_n614), .B2(new_n596), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n606), .A2(G190), .A3(new_n608), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n613), .A2(new_n615), .A3(new_n588), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n586), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n558), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n461), .A2(new_n516), .A3(new_n619), .ZN(G372));
  INV_X1    g0420(.A(new_n448), .ZN(new_n621));
  INV_X1    g0421(.A(new_n424), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(new_n442), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n459), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n447), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n365), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(new_n422), .ZN(new_n628));
  INV_X1    g0428(.A(new_n461), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n598), .A2(new_n610), .A3(new_n611), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n574), .A2(KEYINPUT86), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT86), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n572), .B2(new_n573), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n571), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n315), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n578), .A2(new_n635), .B1(new_n584), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n630), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n584), .A2(new_n636), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(KEYINPUT87), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT87), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n584), .B2(new_n636), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n566), .A2(new_n583), .ZN(new_n645));
  INV_X1    g0445(.A(new_n581), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n585), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n580), .A2(new_n566), .A3(new_n577), .A4(new_n576), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n649), .B2(new_n612), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n639), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n612), .A2(new_n617), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n652), .A2(new_n515), .A3(new_n637), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n511), .A2(new_n478), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n552), .B1(new_n557), .B2(new_n556), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n628), .B1(new_n629), .B2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n511), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n516), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT88), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n516), .A2(KEYINPUT88), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n512), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n665), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n665), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n656), .B(new_n551), .C1(new_n531), .C2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n655), .A2(new_n530), .A3(new_n665), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n511), .A2(new_n478), .A3(new_n675), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n656), .A2(new_n665), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n669), .A2(new_n670), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(G399));
  NAND2_X1  g0485(.A1(new_n563), .A2(new_n517), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT89), .ZN(new_n687));
  INV_X1    g0487(.A(new_n214), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(G1), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n232), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT90), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n658), .B2(new_n665), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n655), .B1(new_n511), .B2(new_n478), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n652), .A2(new_n515), .A3(new_n637), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT90), .B(new_n675), .C1(new_n699), .C2(new_n651), .ZN(new_n700));
  XOR2_X1   g0500(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n652), .B(KEYINPUT93), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n515), .A2(new_n637), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n512), .A2(new_n656), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n578), .A2(new_n635), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n640), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT26), .B1(new_n708), .B2(new_n612), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n630), .A2(new_n586), .A3(new_n638), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n644), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT92), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n709), .A2(new_n713), .A3(new_n710), .A4(new_n644), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT29), .B(new_n675), .C1(new_n706), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n702), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n619), .A2(new_n512), .A3(new_n515), .A4(new_n675), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n570), .A2(new_n405), .A3(new_n574), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n473), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n609), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n550), .A2(new_n720), .A3(KEYINPUT30), .A4(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n634), .A2(new_n405), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n555), .A3(new_n475), .A4(new_n609), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n473), .A2(new_n719), .A3(new_n606), .A4(new_n608), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n555), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n728), .B2(new_n665), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n718), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n717), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n694), .B1(new_n735), .B2(G1), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT94), .Z(G364));
  XNOR2_X1  g0537(.A(new_n679), .B(KEYINPUT95), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n265), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G1), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n689), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n738), .B(new_n744), .C1(G330), .C2(new_n678), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n233), .B1(G20), .B2(new_n315), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n211), .A2(new_n405), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G200), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT97), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n411), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(G190), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT33), .B(G317), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G326), .A2(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n748), .A2(G190), .A3(new_n344), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n748), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n756), .A2(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n211), .A2(G179), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n758), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(G329), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n411), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n211), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n319), .B1(G294), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n762), .A2(new_n411), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n771), .A2(G303), .B1(new_n773), .B2(G283), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n755), .A2(new_n765), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G50), .A2(new_n752), .B1(new_n753), .B2(G68), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n763), .A2(new_n379), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n778), .A2(KEYINPUT32), .B1(new_n219), .B2(new_n770), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n767), .A2(new_n589), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n756), .A2(new_n202), .B1(new_n759), .B2(new_n223), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n603), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n772), .A2(new_n225), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n778), .B2(KEYINPUT32), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n776), .A2(new_n781), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n747), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n746), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n319), .A2(G355), .A3(new_n214), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n688), .A2(new_n385), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n692), .B2(G45), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n251), .A2(G45), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n792), .B1(G116), .B2(new_n214), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n744), .B(new_n787), .C1(new_n791), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n790), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n678), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n745), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n433), .A2(new_n665), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n440), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n442), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n442), .A2(new_n665), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n696), .A2(new_n700), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n806), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n808), .B(new_n675), .C1(new_n699), .C2(new_n651), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n743), .B1(new_n810), .B2(new_n733), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n733), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n746), .A2(new_n788), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n744), .B1(new_n223), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n385), .B1(new_n763), .B2(new_n815), .C1(new_n772), .C2(new_n203), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n767), .A2(new_n202), .B1(new_n770), .B2(new_n231), .ZN(new_n817));
  INV_X1    g0617(.A(new_n756), .ZN(new_n818));
  INV_X1    g0618(.A(new_n759), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(G143), .B1(new_n819), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(new_n753), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  INV_X1    g0622(.A(new_n752), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n820), .B1(new_n821), .B2(new_n355), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT34), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n816), .B(new_n817), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G116), .A2(new_n819), .B1(new_n764), .B2(G311), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n756), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n219), .A2(new_n772), .B1(new_n770), .B2(new_n225), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n830), .A2(new_n319), .A3(new_n831), .A4(new_n780), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G283), .A2(new_n753), .B1(new_n752), .B2(G303), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n826), .A2(new_n827), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n814), .B1(new_n747), .B2(new_n834), .C1(new_n808), .C2(new_n789), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n812), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  INV_X1    g0637(.A(KEYINPUT98), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n459), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(KEYINPUT98), .B(new_n456), .C1(new_n457), .C2(new_n458), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n275), .A2(new_n675), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n622), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n328), .A2(new_n334), .A3(new_n424), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n841), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n846), .A2(new_n732), .A3(new_n808), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n383), .B(new_n391), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n848), .B2(new_n390), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n371), .B1(new_n395), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT99), .ZN(new_n851));
  INV_X1    g0651(.A(new_n663), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT99), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n853), .B(new_n371), .C1(new_n395), .C2(new_n849), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n406), .A3(new_n854), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n415), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n396), .A2(new_n406), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n396), .A2(new_n852), .ZN(new_n861));
  AND4_X1   g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n415), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n855), .B1(new_n447), .B2(new_n448), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n862), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n847), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n396), .B(new_n852), .C1(new_n626), .C2(new_n621), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n860), .A2(new_n861), .A3(new_n415), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT37), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(new_n870), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(KEYINPUT40), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n872), .A2(new_n873), .B1(new_n847), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n461), .A2(new_n732), .ZN(new_n882));
  OAI21_X1  g0682(.A(G330), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n882), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT39), .B1(new_n867), .B2(new_n870), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT100), .ZN(new_n886));
  OR3_X1    g0686(.A1(new_n877), .A2(new_n870), .A3(KEYINPUT39), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT100), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n888), .B(KEYINPUT39), .C1(new_n867), .C2(new_n870), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n665), .B1(new_n839), .B2(new_n840), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n809), .A2(new_n805), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n846), .A2(new_n871), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n626), .A2(new_n663), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n461), .A2(new_n716), .A3(new_n702), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n628), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n896), .B(new_n898), .Z(new_n899));
  OAI22_X1  g0699(.A1(new_n884), .A2(new_n899), .B1(new_n210), .B2(new_n740), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n884), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n593), .A2(KEYINPUT35), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n593), .A2(KEYINPUT35), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(G116), .A3(new_n234), .A4(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT36), .Z(new_n905));
  NAND3_X1  g0705(.A1(new_n232), .A2(G77), .A3(new_n381), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n231), .A2(G68), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n210), .B(G13), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n901), .A2(new_n905), .A3(new_n908), .ZN(G367));
  NAND2_X1  g0709(.A1(new_n771), .A2(G116), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT46), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n385), .B1(new_n819), .B2(G283), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n818), .A2(G303), .B1(new_n764), .B2(G317), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n768), .A2(G107), .B1(new_n773), .B2(new_n562), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n829), .A2(new_n821), .B1(new_n823), .B2(new_n760), .ZN(new_n916));
  INV_X1    g0716(.A(G143), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n917), .A2(new_n823), .B1(new_n821), .B2(new_n379), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n756), .A2(new_n355), .B1(new_n759), .B2(new_n231), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G137), .B2(new_n764), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n603), .B1(G77), .B2(new_n773), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n768), .A2(G68), .B1(new_n771), .B2(G58), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n915), .A2(new_n916), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT47), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n747), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  INV_X1    g0727(.A(new_n793), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n791), .B1(new_n214), .B2(new_n427), .C1(new_n928), .C2(new_n244), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n743), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT104), .Z(new_n931));
  AND2_X1   g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n675), .B1(new_n566), .B2(new_n577), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n708), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n933), .B1(new_n641), .B2(new_n643), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n790), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n935), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n598), .A2(new_n665), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n703), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n630), .A2(new_n665), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n684), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT42), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT101), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n943), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n672), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(KEYINPUT102), .A3(new_n612), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n675), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT102), .B1(new_n949), .B2(new_n612), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n939), .B(new_n946), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT103), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n946), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n938), .B(KEYINPUT43), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n948), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n681), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n961), .A3(new_n958), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n684), .A2(new_n682), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n944), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n684), .A2(new_n682), .A3(new_n943), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n681), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n684), .B1(new_n674), .B2(new_n683), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n738), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n679), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n734), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n969), .A2(new_n681), .A3(new_n972), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n735), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n689), .B(KEYINPUT41), .Z(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n742), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n937), .B1(new_n965), .B2(new_n984), .ZN(G387));
  INV_X1    g0785(.A(new_n978), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n977), .A2(new_n734), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n689), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n977), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n671), .A2(new_n673), .A3(new_n790), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n793), .B1(new_n241), .B2(new_n469), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n319), .A2(new_n214), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n687), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n469), .B1(new_n203), .B2(new_n223), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n354), .A2(G50), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n687), .B(new_n996), .C1(KEYINPUT50), .C2(new_n995), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n993), .A2(new_n997), .B1(new_n225), .B2(new_n688), .ZN(new_n998));
  INV_X1    g0798(.A(new_n791), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n743), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n767), .A2(new_n427), .B1(new_n772), .B2(new_n589), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n756), .A2(new_n231), .B1(new_n763), .B2(new_n355), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n385), .B1(new_n759), .B2(new_n203), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n770), .A2(new_n223), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n821), .B2(new_n354), .C1(new_n379), .C2(new_n823), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G311), .A2(new_n753), .B1(new_n752), .B2(G322), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT105), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(KEYINPUT105), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n818), .A2(G317), .B1(new_n819), .B2(G303), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n767), .A2(new_n521), .B1(new_n770), .B2(new_n829), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n385), .B1(new_n764), .B2(G326), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n517), .C2(new_n772), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT49), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1006), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1000), .B1(new_n1020), .B2(new_n746), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n989), .A2(new_n742), .B1(new_n990), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n988), .A2(new_n1022), .ZN(G393));
  NAND3_X1  g0823(.A1(new_n974), .A2(new_n742), .A3(new_n979), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n791), .B1(new_n214), .B2(new_n519), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n793), .B2(new_n248), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n752), .A2(G150), .B1(G159), .B2(new_n818), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT51), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n385), .B1(new_n763), .B2(new_n917), .C1(new_n759), .C2(new_n354), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n203), .A2(new_n770), .B1(new_n772), .B2(new_n219), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G77), .B2(new_n768), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(new_n821), .C2(new_n231), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n752), .A2(G317), .B1(G311), .B2(new_n818), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n753), .A2(G303), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n770), .A2(new_n521), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n784), .B(new_n1037), .C1(G116), .C2(new_n768), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G294), .A2(new_n819), .B1(new_n764), .B2(G322), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1038), .A3(new_n603), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1028), .A2(new_n1033), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n744), .B(new_n1026), .C1(new_n1041), .C2(new_n746), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n948), .B2(new_n798), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1024), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n979), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n986), .B1(new_n1045), .B2(new_n973), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n980), .A3(new_n689), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT106), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1046), .A2(new_n980), .A3(KEYINPUT106), .A4(new_n689), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1044), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(G390));
  AOI21_X1  g0852(.A(new_n891), .B1(new_n846), .B2(new_n893), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n675), .B(new_n804), .C1(new_n706), .C2(new_n715), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(new_n805), .B1(new_n843), .B2(new_n845), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n891), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n878), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n890), .A2(new_n1053), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n733), .B(new_n806), .C1(new_n843), .C2(new_n845), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(G330), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n718), .B2(new_n731), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n846), .A2(new_n1062), .A3(new_n808), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n1055), .B2(new_n1057), .C1(new_n890), .C2(new_n1053), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n742), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n890), .A2(new_n789), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n772), .A2(new_n203), .B1(new_n763), .B2(new_n829), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT113), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n753), .A2(G107), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n818), .A2(G116), .B1(new_n819), .B2(new_n562), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n768), .A2(G77), .B1(new_n771), .B2(G87), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1070), .A2(new_n603), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1069), .B(new_n1073), .C1(G283), .C2(new_n752), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n770), .A2(new_n355), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT54), .B(G143), .Z(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT111), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1077), .B1(new_n759), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n753), .A2(G137), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n818), .A2(G132), .B1(new_n764), .B2(G125), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n768), .A2(G159), .B1(new_n773), .B2(G50), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1081), .A2(new_n319), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1080), .B(new_n1084), .C1(G128), .C2(new_n752), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n746), .B1(new_n1074), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n813), .A2(new_n354), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n743), .A3(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1065), .A2(new_n1066), .B1(new_n1067), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT109), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n335), .A2(new_n444), .A3(new_n253), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT76), .B1(new_n455), .B2(new_n459), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1062), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n897), .A2(new_n422), .A3(new_n627), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT107), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT107), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n628), .A2(new_n897), .A3(new_n1097), .A4(new_n1094), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1062), .A2(new_n808), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n843), .A2(new_n845), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1054), .A2(new_n805), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1059), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1063), .A2(new_n1100), .B1(new_n805), .B2(new_n809), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1096), .B(new_n1098), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT108), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n893), .B1(new_n1059), .B2(new_n1101), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1063), .A2(new_n805), .A3(new_n1054), .A4(new_n1100), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1110), .A2(KEYINPUT108), .A3(new_n1098), .A4(new_n1096), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1065), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1091), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(KEYINPUT109), .B(new_n1065), .C1(new_n1107), .C2(new_n1111), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT110), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1107), .A2(new_n1118), .A3(new_n1065), .A4(new_n1111), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n689), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1090), .B1(new_n1116), .B2(new_n1120), .ZN(G378));
  INV_X1    g0921(.A(new_n454), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n419), .A2(new_n852), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT55), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n1126));
  NAND2_X1  g0926(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1126), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT117), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1132), .A2(new_n788), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT118), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n813), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n743), .B1(G50), .B2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n753), .A2(G97), .B1(new_n582), .B2(new_n819), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT114), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n752), .A2(G116), .B1(G68), .B2(new_n768), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT115), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n385), .A2(G41), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n225), .B2(new_n756), .C1(new_n521), .C2(new_n763), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1004), .B(new_n1142), .C1(G58), .C2(new_n773), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT58), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n379), .B2(new_n772), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n756), .A2(new_n1149), .B1(new_n759), .B2(new_n822), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1079), .A2(new_n770), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G150), .C2(new_n768), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n752), .A2(G125), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n815), .C2(new_n821), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1148), .B1(new_n1154), .B2(KEYINPUT59), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(KEYINPUT59), .B2(new_n1154), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1145), .A2(KEYINPUT58), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1141), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1158), .B(new_n231), .C1(G33), .C2(G41), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1146), .A2(new_n1156), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1136), .B1(new_n1160), .B2(new_n746), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OR3_X1    g0962(.A1(new_n1133), .A2(new_n1134), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1134), .B1(new_n1133), .B2(new_n1162), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1131), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n881), .B2(new_n1061), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n880), .A2(G330), .A3(new_n1132), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1166), .A2(new_n896), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n896), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1163), .B(new_n1164), .C1(new_n1170), .C2(new_n1066), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT108), .B1(new_n1173), .B2(new_n1110), .ZN(new_n1175));
  AND4_X1   g0975(.A1(KEYINPUT108), .A2(new_n1110), .A3(new_n1098), .A4(new_n1096), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1113), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT109), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1112), .A2(new_n1091), .A3(new_n1113), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1172), .B1(new_n1180), .B2(new_n1170), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n896), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1166), .A2(new_n896), .A3(new_n1167), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1172), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1173), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n690), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1171), .B1(new_n1181), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n1110), .A2(new_n742), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n743), .B1(G68), .B2(new_n1135), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G116), .A2(new_n753), .B1(new_n752), .B2(G294), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n756), .A2(new_n521), .B1(new_n759), .B2(new_n225), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G303), .B2(new_n764), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n319), .B1(G77), .B2(new_n773), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n768), .A2(new_n582), .B1(new_n771), .B2(G97), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n385), .B1(new_n772), .B2(new_n202), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT120), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n759), .A2(new_n355), .B1(new_n763), .B2(new_n1149), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G50), .B2(new_n768), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(new_n379), .C2(new_n770), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT121), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n752), .A2(G132), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n822), .B2(new_n756), .C1(new_n821), .C2(new_n1079), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1198), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1192), .B1(new_n1207), .B2(new_n746), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n846), .B2(new_n789), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1191), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1173), .A2(new_n1110), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT119), .Z(new_n1212));
  NOR2_X1   g1012(.A1(new_n1112), .A2(new_n982), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1210), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(G381));
  AND3_X1   g1015(.A1(new_n954), .A2(new_n961), .A3(new_n958), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n961), .B1(new_n954), .B2(new_n958), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n984), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1218), .A2(new_n1219), .B1(new_n936), .B2(new_n932), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G393), .A2(G396), .ZN(new_n1221));
  AND4_X1   g1021(.A1(new_n836), .A2(new_n1220), .A3(new_n1051), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(G378), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1189), .A4(new_n1214), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n664), .A2(G213), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT122), .Z(new_n1226));
  NAND3_X1  g1026(.A1(new_n1189), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(G407), .A2(G213), .A3(new_n1227), .ZN(G409));
  AOI21_X1  g1028(.A(new_n800), .B1(new_n988), .B2(new_n1022), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1221), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1220), .A2(G390), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G387), .A2(new_n1051), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT126), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1231), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(KEYINPUT126), .B(new_n1230), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1187), .A2(new_n983), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1239), .B2(new_n742), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G378), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT123), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1189), .B2(G378), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n689), .B1(new_n1180), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1239), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1242), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(KEYINPUT123), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1244), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1226), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(KEYINPUT127), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT127), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1250), .A2(KEYINPUT123), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1181), .A2(new_n1188), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1257), .A2(new_n1245), .A3(G378), .A4(new_n1242), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1243), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1255), .B1(new_n1259), .B2(new_n1226), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n690), .B1(new_n1211), .B2(KEYINPUT60), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1111), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1212), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT124), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1212), .A2(new_n1266), .A3(new_n1263), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1262), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  OR3_X1    g1068(.A1(new_n1268), .A2(new_n836), .A3(new_n1210), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n836), .B1(new_n1268), .B2(new_n1210), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1254), .A2(new_n1260), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1272), .B1(new_n1275), .B2(new_n1271), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1226), .A2(G2897), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1278), .B(KEYINPUT125), .Z(new_n1279));
  AND3_X1   g1079(.A1(new_n1269), .A2(new_n1270), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT127), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1259), .A2(new_n1255), .A3(new_n1226), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1238), .B1(new_n1277), .B2(new_n1287), .ZN(new_n1288));
  OR3_X1    g1088(.A1(new_n1236), .A2(new_n1237), .A3(KEYINPUT61), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1275), .B2(new_n1282), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1271), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1254), .A2(new_n1260), .A3(KEYINPUT63), .A4(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1275), .A2(new_n1271), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1290), .B(new_n1292), .C1(KEYINPUT63), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1288), .A2(new_n1294), .ZN(G405));
  AOI22_X1  g1095(.A1(new_n1256), .A2(new_n1258), .B1(new_n1223), .B2(G375), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1238), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1238), .A2(new_n1296), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1291), .ZN(G402));
endmodule


