//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(G8gat), .B1(new_n204), .B2(KEYINPUT88), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G1gat), .B2(new_n203), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n205), .B(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT86), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n216), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n218), .B2(new_n219), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n212), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  INV_X1    g023(.A(new_n212), .ZN(new_n225));
  INV_X1    g024(.A(new_n214), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(new_n213), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n211), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n225), .A2(new_n221), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n223), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n224), .B1(new_n223), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n209), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT89), .B(new_n209), .C1(new_n230), .C2(new_n231), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n223), .A2(new_n229), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT90), .B1(new_n239), .B2(new_n209), .ZN(new_n240));
  INV_X1    g039(.A(new_n209), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n229), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n238), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI211_X1 g047(.A(new_n247), .B(new_n238), .C1(new_n240), .C2(new_n244), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n240), .A2(new_n244), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n239), .A2(new_n209), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n237), .B(KEYINPUT13), .Z(new_n253));
  AOI22_X1  g052(.A1(new_n249), .A2(new_n236), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT12), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n248), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n248), .B2(new_n254), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n202), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n254), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n259), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n254), .A3(new_n260), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT91), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(G99gat), .A2(G106gat), .ZN(new_n271));
  INV_X1    g070(.A(G85gat), .ZN(new_n272));
  INV_X1    g071(.A(G92gat), .ZN(new_n273));
  AOI22_X1  g072(.A1(KEYINPUT8), .A2(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n272), .B2(new_n273), .ZN(new_n276));
  NAND4_X1  g075(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G99gat), .B(G106gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n274), .A2(new_n279), .A3(new_n276), .A4(new_n277), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n281), .A2(KEYINPUT98), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT98), .B1(new_n281), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n270), .B1(new_n239), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n230), .A2(new_n231), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n286), .ZN(new_n289));
  XOR2_X1   g088(.A(G190gat), .B(G218gat), .Z(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G134gat), .B(G162gat), .Z(new_n294));
  AOI21_X1  g093(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n296), .A2(KEYINPUT101), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n292), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(KEYINPUT101), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n300), .B(KEYINPUT102), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n302), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G57gat), .B(G64gat), .Z(new_n307));
  NAND2_X1  g106(.A1(G71gat), .A2(G78gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT92), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT93), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  OR2_X1    g113(.A1(G71gat), .A2(G78gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n316));
  AND4_X1   g115(.A1(new_n312), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n314), .A2(new_n316), .B1(new_n315), .B2(new_n312), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n308), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n315), .A2(KEYINPUT94), .A3(new_n308), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(new_n310), .A3(new_n307), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G231gat), .A2(G233gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G127gat), .B(G155gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT20), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n329), .B(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n209), .B1(new_n326), .B2(new_n325), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT96), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n332), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G183gat), .B(G211gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n335), .B(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n306), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G120gat), .B(G148gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G176gat), .B(G204gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G230gat), .A2(G233gat), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n281), .A2(new_n282), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n279), .A2(KEYINPUT103), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(new_n319), .A3(new_n324), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n319), .A2(new_n324), .A3(new_n348), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n281), .A2(new_n282), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n346), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n353), .A2(KEYINPUT104), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n352), .ZN(new_n355));
  INV_X1    g154(.A(new_n346), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT104), .A3(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n352), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n325), .A2(new_n360), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n285), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n356), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n345), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n346), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n354), .A2(KEYINPUT105), .A3(new_n357), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT105), .B1(new_n354), .B2(new_n357), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n344), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n341), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT77), .ZN(new_n378));
  XNOR2_X1  g177(.A(G197gat), .B(G204gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380));
  INV_X1    g179(.A(G211gat), .ZN(new_n381));
  INV_X1    g180(.A(G218gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n377), .A2(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n377), .A2(KEYINPUT77), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n386), .A2(new_n383), .A3(new_n379), .A4(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT26), .ZN(new_n392));
  NAND2_X1  g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT71), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT70), .ZN(new_n400));
  INV_X1    g199(.A(G183gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT27), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G183gat), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n400), .B1(new_n403), .B2(G183gat), .ZN(new_n406));
  INV_X1    g205(.A(G190gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n399), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(G190gat), .B1(new_n402), .B2(new_n400), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT27), .B(G183gat), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n410), .B(KEYINPUT71), .C1(new_n400), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT28), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(KEYINPUT28), .A3(new_n407), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n398), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n414), .A2(KEYINPUT72), .A3(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n391), .A2(KEYINPUT23), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n391), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT67), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n391), .A2(KEYINPUT23), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n424), .A3(new_n395), .A4(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n395), .A2(new_n427), .A3(new_n421), .A4(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT67), .ZN(new_n430));
  INV_X1    g229(.A(new_n397), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n432));
  OAI211_X1 g231(.A(KEYINPUT64), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n433));
  MUX2_X1   g232(.A(new_n431), .B(new_n432), .S(new_n433), .Z(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT25), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n395), .B(KEYINPUT68), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n397), .A2(KEYINPUT69), .A3(KEYINPUT24), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(KEYINPUT23), .B2(new_n391), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n401), .A2(new_n407), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n441), .B(new_n397), .C1(KEYINPUT69), .C2(KEYINPUT24), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT25), .A4(new_n421), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n437), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G226gat), .ZN(new_n447));
  INV_X1    g246(.A(G233gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n420), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n420), .A2(new_n446), .B1(new_n453), .B2(new_n450), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n390), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n414), .A2(KEYINPUT72), .A3(new_n415), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT72), .B1(new_n414), .B2(new_n415), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(new_n398), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n444), .B1(new_n435), .B2(new_n436), .ZN(new_n459));
  OAI22_X1  g258(.A1(new_n458), .A2(new_n459), .B1(KEYINPUT29), .B2(new_n449), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n389), .A3(new_n451), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n455), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n460), .A2(KEYINPUT78), .A3(new_n389), .A4(new_n451), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n376), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n375), .B(KEYINPUT79), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  OAI22_X1  g267(.A1(new_n465), .A2(KEYINPUT30), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G127gat), .B(G134gat), .Z(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G120gat), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n472), .A2(KEYINPUT1), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n472), .A2(KEYINPUT1), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT73), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(KEYINPUT73), .A3(new_n471), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(G141gat), .B(G148gat), .Z(new_n481));
  XNOR2_X1  g280(.A(G155gat), .B(G162gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT2), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT80), .B(G155gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n485), .B2(G162gat), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n482), .ZN(new_n488));
  INV_X1    g287(.A(new_n481), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(KEYINPUT2), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n480), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G225gat), .A2(G233gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT5), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n480), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n487), .A2(new_n496), .A3(new_n490), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n487), .A2(new_n490), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n493), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G1gat), .B(G29gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT0), .ZN(new_n508));
  XNOR2_X1  g307(.A(G57gat), .B(G85gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n501), .B(KEYINPUT4), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(KEYINPUT5), .A3(new_n493), .A4(new_n499), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n511), .B1(new_n506), .B2(new_n513), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n465), .A2(KEYINPUT30), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n470), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT34), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n480), .B1(new_n458), .B2(new_n459), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n420), .A2(new_n446), .A3(new_n495), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G227gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(new_n448), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n523), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  AOI211_X1 g329(.A(KEYINPUT34), .B(new_n528), .C1(new_n524), .C2(new_n525), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(new_n528), .A3(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT33), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G15gat), .B(G43gat), .Z(new_n537));
  XNOR2_X1  g336(.A(G71gat), .B(G99gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n533), .B(KEYINPUT32), .C1(new_n535), .C2(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n532), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n532), .B1(new_n542), .B2(new_n540), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n389), .B1(new_n453), .B2(new_n497), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n385), .A2(new_n453), .A3(new_n388), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n500), .B1(new_n496), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(G228gat), .B(G233gat), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n497), .A2(new_n453), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT83), .B1(new_n552), .B2(new_n389), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT82), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G228gat), .A2(G233gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n548), .B2(new_n554), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n549), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G50gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G78gat), .B(G106gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n560), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n549), .B(new_n564), .C1(new_n556), .C2(new_n558), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n561), .B2(new_n565), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR4_X1   g367(.A1(new_n522), .A2(new_n545), .A3(KEYINPUT35), .A4(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n543), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT75), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n540), .A2(new_n542), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT74), .ZN(new_n573));
  INV_X1    g372(.A(new_n532), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n540), .A2(new_n575), .A3(new_n542), .ZN(new_n576));
  AND4_X1   g375(.A1(new_n571), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n532), .B1(new_n572), .B2(KEYINPUT74), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n571), .B1(new_n578), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n570), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT85), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n522), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n570), .B(KEYINPUT85), .C1(new_n577), .C2(new_n579), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n569), .B1(new_n585), .B2(KEYINPUT35), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n522), .A2(new_n568), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n514), .A2(new_n515), .ZN(new_n588));
  INV_X1    g387(.A(new_n518), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n516), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n465), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n466), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n461), .A2(KEYINPUT84), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n455), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n461), .A2(KEYINPUT84), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT37), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n594), .A2(new_n598), .A3(new_n467), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n463), .A2(KEYINPUT37), .A3(new_n464), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n594), .A2(KEYINPUT38), .A3(new_n376), .A4(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n592), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n504), .A2(new_n605), .A3(new_n505), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n493), .B1(new_n512), .B2(new_n499), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n492), .A2(new_n493), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT39), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n606), .B(new_n510), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n504), .A2(new_n505), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(KEYINPUT39), .A3(new_n608), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n614), .A2(KEYINPUT40), .A3(new_n510), .A4(new_n606), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n612), .A2(new_n615), .A3(new_n514), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n465), .A2(KEYINPUT30), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n469), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n568), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n587), .B1(new_n604), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n543), .B2(new_n544), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT76), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT76), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n625), .B(new_n622), .C1(new_n543), .C2(new_n544), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n543), .A2(new_n622), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n577), .B2(new_n579), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n621), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n269), .B(new_n372), .C1(new_n586), .C2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n590), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g433(.A1(new_n470), .A2(new_n521), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n631), .A2(KEYINPUT106), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT106), .B1(new_n631), .B2(new_n636), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(G8gat), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT16), .B(G8gat), .Z(new_n640));
  NAND4_X1  g439(.A1(new_n632), .A2(KEYINPUT42), .A3(new_n635), .A4(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n637), .B2(new_n638), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n639), .B(new_n641), .C1(new_n643), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g443(.A(KEYINPUT108), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n629), .A2(new_n627), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n629), .B2(new_n627), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n632), .A2(G15gat), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n651));
  INV_X1    g450(.A(new_n569), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n630), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n545), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n269), .A4(new_n372), .ZN(new_n657));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT107), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(KEYINPUT107), .B(new_n658), .C1(new_n631), .C2(new_n545), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n650), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(KEYINPUT109), .B(new_n650), .C1(new_n659), .C2(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n631), .A2(new_n619), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR3_X1   g468(.A1(new_n646), .A2(new_n647), .A3(new_n621), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n306), .B1(new_n586), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n306), .C1(new_n586), .C2(new_n630), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n371), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n339), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n265), .A2(new_n266), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681), .B2(new_n520), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n677), .A2(new_n305), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n269), .B(new_n683), .C1(new_n586), .C2(new_n630), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n520), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT45), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(G1328gat));
  OAI21_X1  g486(.A(G36gat), .B1(new_n681), .B2(new_n636), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n684), .A2(G36gat), .A3(new_n636), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT46), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1329gat));
  INV_X1    g490(.A(G43gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n648), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n673), .A2(new_n674), .A3(new_n680), .A4(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n684), .B2(new_n545), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g496(.A1(new_n673), .A2(new_n568), .A3(new_n674), .A4(new_n680), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G50gat), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n268), .B1(new_n653), .B2(new_n654), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n619), .A2(G50gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n683), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n699), .A2(KEYINPUT48), .A3(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n700), .A2(KEYINPUT111), .A3(new_n683), .A4(new_n701), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705));
  INV_X1    g504(.A(new_n701), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n684), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(G50gat), .B2(new_n698), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n710));
  OAI21_X1  g509(.A(new_n703), .B1(new_n709), .B2(new_n710), .ZN(G1331gat));
  INV_X1    g510(.A(new_n621), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n648), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n653), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n341), .A2(new_n678), .A3(new_n676), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n590), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n635), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT49), .B(G64gat), .Z(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n716), .A2(new_n723), .A3(new_n656), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n714), .A2(new_n715), .ZN(new_n725));
  OAI21_X1  g524(.A(G71gat), .B1(new_n725), .B2(new_n648), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n716), .A2(new_n568), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  INV_X1    g530(.A(new_n339), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n678), .A3(new_n676), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n675), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734), .B2(new_n520), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n305), .B1(new_n653), .B2(new_n713), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(new_n678), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n306), .B(new_n737), .C1(new_n586), .C2(new_n670), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n744), .A2(new_n272), .A3(new_n590), .A4(new_n371), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n735), .A2(new_n745), .ZN(G1336gat));
  NOR3_X1   g545(.A1(new_n636), .A2(G92gat), .A3(new_n676), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n673), .A2(new_n635), .A3(new_n674), .A4(new_n733), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n714), .A2(KEYINPUT51), .A3(new_n306), .A4(new_n737), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n743), .ZN(new_n754));
  AOI22_X1  g553(.A1(G92gat), .A2(new_n749), .B1(new_n754), .B2(new_n747), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n748), .A2(new_n752), .B1(new_n755), .B2(new_n751), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n734), .B2(new_n648), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n545), .A2(G99gat), .A3(new_n676), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n744), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1338gat));
  NOR3_X1   g559(.A1(new_n619), .A2(G106gat), .A3(new_n676), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n744), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n673), .A2(new_n568), .A3(new_n674), .A4(new_n733), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G106gat), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI22_X1  g565(.A1(G106gat), .A2(new_n763), .B1(new_n754), .B2(new_n761), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n762), .A2(new_n766), .B1(new_n767), .B2(new_n765), .ZN(G1339gat));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n346), .B1(new_n285), .B2(new_n362), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n361), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n769), .B1(new_n367), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n774));
  AOI21_X1  g573(.A(new_n344), .B1(new_n364), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n773), .A2(KEYINPUT114), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n367), .A2(new_n772), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n775), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n769), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n370), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n678), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n252), .A2(new_n253), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n237), .B1(new_n236), .B2(new_n250), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n258), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n266), .A3(new_n371), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n306), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n793), .A2(new_n266), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(new_n786), .A3(new_n306), .A4(new_n787), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n339), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n372), .A2(new_n679), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n545), .A2(new_n568), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n635), .A2(new_n520), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(G113gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n805), .A3(new_n268), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n520), .B1(new_n799), .B2(new_n800), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n582), .A2(new_n584), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n807), .A2(new_n636), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n678), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n806), .B1(new_n810), .B2(new_n805), .ZN(G1340gat));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n804), .A2(new_n812), .A3(new_n676), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n371), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n812), .ZN(G1341gat));
  INV_X1    g614(.A(G127gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n809), .A2(new_n816), .A3(new_n732), .ZN(new_n817));
  OAI21_X1  g616(.A(G127gat), .B1(new_n804), .B2(new_n339), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1342gat));
  INV_X1    g618(.A(G134gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n809), .A2(new_n820), .A3(new_n306), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n821), .A2(KEYINPUT56), .ZN(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n804), .B2(new_n305), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(KEYINPUT56), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(G1343gat));
  AND2_X1   g624(.A1(new_n648), .A2(new_n803), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n568), .A2(KEYINPUT57), .ZN(new_n827));
  INV_X1    g626(.A(new_n800), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n782), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n781), .A2(new_n775), .A3(KEYINPUT117), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n769), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n780), .A2(new_n832), .A3(new_n370), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n780), .A2(new_n832), .A3(KEYINPUT118), .A4(new_n370), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n263), .A3(new_n267), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n306), .B1(new_n837), .B2(new_n794), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n797), .B1(new_n838), .B2(KEYINPUT119), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n840), .B(new_n306), .C1(new_n837), .C2(new_n794), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n339), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n828), .B1(new_n842), .B2(KEYINPUT120), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n339), .C1(new_n839), .C2(new_n841), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n827), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n801), .B2(new_n568), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n269), .B(new_n826), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n646), .A2(new_n647), .A3(new_n619), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n807), .A2(new_n636), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n268), .A2(G141gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n678), .B(new_n826), .C1(new_n846), .C2(new_n847), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n856), .A2(G141gat), .B1(new_n852), .B2(new_n853), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(G1344gat));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n801), .B2(new_n568), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n568), .A2(new_n860), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n305), .B2(new_n784), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n796), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n305), .A2(new_n863), .A3(new_n784), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n339), .B1(new_n867), .B2(new_n838), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n372), .A2(new_n268), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n861), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n371), .A3(new_n826), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G148gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT59), .ZN(new_n874));
  INV_X1    g673(.A(G148gat), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(KEYINPUT59), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n826), .B1(new_n846), .B2(new_n847), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n676), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n852), .A2(new_n875), .A3(new_n371), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1345gat));
  OAI21_X1  g680(.A(new_n485), .B1(new_n877), .B2(new_n339), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n339), .A2(new_n485), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n852), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1346gat));
  OAI21_X1  g684(.A(G162gat), .B1(new_n877), .B2(new_n305), .ZN(new_n886));
  INV_X1    g685(.A(G162gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n852), .A2(new_n887), .A3(new_n306), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1347gat));
  AOI21_X1  g690(.A(new_n590), .B1(new_n799), .B2(new_n800), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n892), .A2(new_n635), .A3(new_n808), .ZN(new_n893));
  AOI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n678), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n636), .A2(new_n590), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n801), .A2(new_n802), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT124), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n269), .A2(G169gat), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G1348gat));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n896), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G176gat), .B1(new_n901), .B2(new_n676), .ZN(new_n902));
  INV_X1    g701(.A(G176gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n893), .A2(new_n903), .A3(new_n371), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1349gat));
  AOI21_X1  g704(.A(new_n401), .B1(new_n897), .B2(new_n732), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n893), .A2(new_n411), .A3(new_n732), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G183gat), .B1(new_n901), .B2(new_n339), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n911), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n901), .B2(new_n305), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n893), .A2(new_n407), .A3(new_n306), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT125), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT61), .B(G190gat), .C1(new_n901), .C2(new_n305), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(G1351gat));
  AND2_X1   g719(.A1(new_n851), .A2(new_n635), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n892), .ZN(new_n922));
  AOI21_X1  g721(.A(G197gat), .B1(new_n922), .B2(new_n678), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n648), .A2(new_n895), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n871), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n269), .A2(G197gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n676), .A2(G204gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n921), .A2(new_n892), .A3(new_n928), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT62), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n861), .A2(new_n676), .A3(new_n870), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n924), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT126), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n935), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n931), .A4(new_n930), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n871), .A2(new_n732), .A3(new_n924), .ZN(new_n941));
  NOR2_X1   g740(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(G211gat), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n922), .A2(new_n381), .A3(new_n732), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n941), .A2(G211gat), .ZN(new_n945));
  XNOR2_X1  g744(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n943), .B(new_n944), .C1(new_n945), .C2(new_n946), .ZN(G1354gat));
  NAND3_X1  g746(.A1(new_n922), .A2(new_n382), .A3(new_n306), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n925), .A2(new_n306), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n382), .ZN(G1355gat));
endmodule


