//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n214), .B1(new_n217), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n209), .A2(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n251), .B1(new_n227), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n215), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n253), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT11), .B1(new_n253), .B2(new_n255), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT74), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT74), .B1(new_n256), .B2(new_n257), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n255), .B1(new_n208), .B2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT12), .B1(new_n263), .B2(G68), .ZN(new_n265));
  AOI22_X1  g0065(.A1(G68), .A2(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n260), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT14), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT13), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT65), .B1(new_n274), .B2(new_n277), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT73), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n222), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT73), .B1(new_n278), .B2(new_n279), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  OAI211_X1 g0086(.A(G232), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  OAI211_X1 g0088(.A(G226), .B(new_n288), .C1(new_n285), .C2(new_n286), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G97), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT72), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT72), .A4(new_n290), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n274), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n269), .B1(new_n284), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n274), .A2(new_n277), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT65), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n277), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n281), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n283), .A2(new_n302), .A3(G238), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n275), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n304), .A2(KEYINPUT13), .A3(new_n295), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n268), .B(G169), .C1(new_n297), .C2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n284), .A2(new_n269), .A3(new_n296), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT13), .B1(new_n304), .B2(new_n295), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n308), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n268), .B1(new_n311), .B2(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n267), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(G223), .B(new_n288), .C1(new_n285), .C2(new_n286), .ZN(new_n314));
  OAI211_X1 g0114(.A(G226), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n315));
  INV_X1    g0115(.A(G33), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(new_n223), .ZN(new_n317));
  INV_X1    g0117(.A(new_n274), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n274), .A2(G232), .A3(new_n277), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n275), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(G200), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT16), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT3), .B(G33), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(G20), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n285), .A2(new_n286), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n221), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G58), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n221), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n335), .B2(new_n201), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n250), .A2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n327), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n331), .B2(new_n209), .ZN(new_n340));
  NOR4_X1   g0140(.A1(new_n285), .A2(new_n286), .A3(new_n328), .A4(G20), .ZN(new_n341));
  OAI21_X1  g0141(.A(G68), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n338), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(KEYINPUT16), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n344), .A3(new_n255), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n334), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT8), .B(G58), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(KEYINPUT66), .ZN(new_n348));
  INV_X1    g0148(.A(new_n263), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n262), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n326), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT17), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n326), .A2(new_n345), .A3(KEYINPUT17), .A4(new_n353), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n356), .A2(KEYINPUT75), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT75), .B1(new_n356), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n267), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n311), .B2(new_n320), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n307), .B2(new_n308), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n255), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n342), .A2(new_n343), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n327), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n352), .B1(new_n368), .B2(new_n344), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n325), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G169), .B2(new_n325), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n369), .A2(KEYINPUT18), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n325), .A2(G169), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n370), .B2(new_n325), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n345), .A2(new_n353), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n313), .A2(new_n360), .A3(new_n365), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n300), .A2(new_n301), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n276), .B1(new_n381), .B2(G226), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n329), .A2(G222), .A3(new_n288), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n329), .A2(G223), .A3(G1698), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n384), .C1(new_n227), .C2(new_n329), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n318), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n370), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n263), .A2(G50), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n262), .B2(G50), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n250), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n252), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n348), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(new_n366), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n389), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n363), .B1(new_n382), .B2(new_n386), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n388), .B2(G190), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT70), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n391), .C1(new_n395), .C2(new_n366), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n348), .A2(new_n394), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n366), .B1(new_n405), .B2(new_n392), .ZN(new_n406));
  INV_X1    g0206(.A(new_n391), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT70), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n409), .B1(new_n404), .B2(new_n408), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n401), .B(new_n402), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n404), .A2(new_n408), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT9), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n410), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n402), .B1(new_n417), .B2(new_n401), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n399), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n329), .A2(G232), .A3(new_n288), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n329), .A2(G238), .A3(G1698), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n229), .C2(new_n329), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n318), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n381), .A2(G244), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n275), .A3(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(new_n320), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(G200), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n347), .B(KEYINPUT67), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n428), .A2(new_n250), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n252), .B1(new_n209), .B2(new_n227), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n255), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n349), .A2(KEYINPUT68), .A3(new_n227), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT68), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n263), .B2(G77), .ZN(new_n435));
  AOI22_X1  g0235(.A1(G77), .A2(new_n262), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n426), .A2(new_n427), .A3(new_n432), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n436), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n423), .A2(new_n370), .A3(new_n424), .A4(new_n275), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n425), .A2(new_n397), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT69), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT69), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT71), .B1(new_n419), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n399), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n401), .B1(new_n411), .B2(new_n412), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT10), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(new_n413), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT71), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n445), .A4(new_n443), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n380), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n208), .B(G45), .C1(new_n270), .C2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G41), .ZN(new_n458));
  OAI211_X1 g0258(.A(G270), .B(new_n274), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT76), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n271), .A2(G1), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n457), .A2(G41), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(KEYINPUT76), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n467));
  AND2_X1   g0267(.A1(G33), .A2(G41), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(G274), .C1(new_n468), .C2(new_n215), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT77), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n469), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT77), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(new_n465), .A4(new_n462), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n460), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g0274(.A1(KEYINPUT3), .A2(G33), .ZN(new_n475));
  INV_X1    g0275(.A(G303), .ZN(new_n476));
  NAND2_X1  g0276(.A1(KEYINPUT3), .A2(G33), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n318), .ZN(new_n479));
  INV_X1    g0279(.A(G257), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n288), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n230), .A2(G1698), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n481), .A2(new_n482), .B1(new_n475), .B2(new_n477), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n474), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n209), .C1(G33), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G20), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n255), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n489), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n263), .A2(G116), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n316), .A2(G1), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n349), .A2(new_n255), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(G116), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G179), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n455), .B1(new_n486), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n460), .B(new_n484), .C1(new_n470), .C2(new_n473), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n370), .B1(new_n496), .B2(new_n500), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(KEYINPUT81), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n501), .A2(G169), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n486), .A2(new_n501), .A3(KEYINPUT21), .A4(G169), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n474), .A2(G190), .A3(new_n485), .ZN(new_n512));
  INV_X1    g0312(.A(new_n501), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n513), .C1(new_n504), .C2(new_n363), .ZN(new_n514));
  AND4_X1   g0314(.A1(new_n507), .A2(new_n510), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n329), .A2(new_n209), .A3(G68), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n209), .B1(new_n290), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G87), .B2(new_n206), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(new_n252), .B2(new_n488), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(new_n255), .B1(new_n349), .B2(new_n430), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n222), .A2(new_n288), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n228), .A2(G1698), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n285), .C2(new_n286), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n316), .A2(new_n490), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n274), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G274), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n463), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n224), .B1(new_n271), .B2(G1), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n274), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(G200), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n499), .A2(G87), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n522), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n528), .A2(new_n533), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT80), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(G190), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n523), .A2(new_n524), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n526), .B1(new_n540), .B2(new_n329), .ZN(new_n541));
  OAI211_X1 g0341(.A(G190), .B(new_n532), .C1(new_n541), .C2(new_n274), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT80), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n536), .A2(KEYINPUT79), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT79), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n522), .A2(new_n534), .A3(new_n545), .A4(new_n535), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n397), .B1(new_n528), .B2(new_n533), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n521), .A2(new_n255), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n430), .A2(new_n349), .ZN(new_n549));
  INV_X1    g0349(.A(new_n430), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n499), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n537), .A2(new_n370), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n544), .A2(new_n546), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n470), .A2(new_n473), .ZN(new_n556));
  OAI211_X1 g0356(.A(G244), .B(new_n288), .C1(new_n285), .C2(new_n286), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n329), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n329), .A2(G250), .A3(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n487), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n318), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(new_n274), .C1(new_n456), .C2(new_n458), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT78), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n556), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n397), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n488), .A2(new_n229), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n205), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n229), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n250), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n340), .B2(new_n341), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n255), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n263), .A2(G97), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n499), .B2(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n556), .A2(new_n563), .A3(new_n566), .A4(new_n370), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n568), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n209), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n229), .A2(KEYINPUT23), .A3(G20), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n585), .B1(new_n526), .B2(new_n209), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n209), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g0390(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n591), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n587), .B(KEYINPUT22), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(new_n586), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n255), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT25), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n263), .A2(new_n597), .A3(G107), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n263), .B2(G107), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n499), .A2(G107), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G264), .B(new_n274), .C1(new_n456), .C2(new_n458), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n224), .A2(new_n288), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n480), .A2(G1698), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n285), .C2(new_n286), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n606), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n318), .A3(new_n610), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n320), .A2(new_n556), .A3(new_n602), .A4(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n602), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n274), .B1(new_n607), .B2(new_n608), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n610), .ZN(new_n615));
  AOI21_X1  g0415(.A(G200), .B1(new_n615), .B2(new_n556), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n596), .B(new_n601), .C1(new_n612), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n556), .A2(new_n611), .A3(new_n602), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n397), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n615), .A2(new_n370), .A3(new_n556), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n590), .A2(new_n591), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n594), .A2(new_n586), .A3(new_n593), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n366), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n601), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n619), .B(new_n620), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n567), .A2(G200), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n556), .A2(new_n563), .A3(new_n566), .A4(G190), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n577), .A3(new_n579), .A4(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n582), .A2(new_n617), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n454), .A2(new_n515), .A3(new_n555), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n441), .ZN(new_n631));
  OAI21_X1  g0431(.A(G169), .B1(new_n297), .B2(new_n305), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n309), .A3(new_n306), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n634), .B2(new_n267), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n360), .A2(new_n365), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n379), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n450), .A2(new_n413), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n448), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n454), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n552), .A2(new_n553), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT84), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n643), .B(new_n274), .C1(new_n525), .C2(new_n527), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n532), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n397), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n641), .B1(new_n646), .B2(KEYINPUT85), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT85), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n648), .A3(new_n397), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n548), .A2(new_n549), .A3(new_n535), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n522), .A2(KEYINPUT86), .A3(new_n535), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n539), .A2(new_n543), .B1(new_n645), .B2(G200), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n647), .A2(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(new_n582), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n643), .B1(new_n541), .B2(new_n274), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n533), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT85), .B1(new_n662), .B2(G169), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n649), .A3(new_n554), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n536), .A2(KEYINPUT79), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n539), .A2(new_n543), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n546), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n554), .A2(new_n547), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT26), .B1(new_n669), .B2(new_n582), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n659), .A2(new_n664), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n486), .A2(new_n502), .A3(new_n455), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT81), .B1(new_n504), .B2(new_n505), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n511), .A2(new_n510), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n507), .A2(KEYINPUT87), .A3(new_n510), .A4(new_n511), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n625), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n617), .A2(new_n628), .A3(new_n582), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n655), .A2(new_n654), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n664), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n671), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n639), .B1(new_n640), .B2(new_n685), .ZN(G369));
  AND2_X1   g0486(.A1(new_n677), .A2(new_n678), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n501), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT88), .Z(new_n695));
  MUX2_X1   g0495(.A(new_n515), .B(new_n687), .S(new_n695), .Z(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n617), .A2(new_n625), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n693), .B1(new_n623), .B2(new_n624), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n693), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n625), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n701), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(new_n698), .ZN(new_n706));
  INV_X1    g0506(.A(new_n625), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n701), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(G399));
  NAND2_X1  g0509(.A1(new_n212), .A2(new_n270), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n205), .A2(new_n223), .A3(new_n490), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT89), .Z(new_n713));
  NOR3_X1   g0513(.A1(new_n711), .A2(new_n713), .A3(new_n208), .ZN(new_n714));
  INV_X1    g0514(.A(new_n219), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n711), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT28), .Z(new_n717));
  NAND4_X1  g0517(.A1(new_n629), .A2(new_n515), .A3(new_n555), .A4(new_n701), .ZN(new_n718));
  XNOR2_X1  g0518(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n719));
  OAI21_X1  g0519(.A(G179), .B1(new_n479), .B2(new_n483), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n720), .A2(new_n528), .A3(new_n533), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n615), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n556), .A2(new_n563), .A3(new_n566), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT90), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n474), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n615), .A2(new_n474), .A3(new_n721), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT90), .B1(new_n726), .B2(new_n567), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n719), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n662), .A2(G179), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n486), .A3(new_n567), .A4(new_n618), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT30), .A4(new_n474), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n693), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT31), .B(new_n693), .C1(new_n728), .C2(new_n732), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n718), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n685), .B2(new_n693), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n628), .A2(new_n582), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n617), .A3(new_n656), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n704), .A2(new_n707), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT26), .B1(new_n683), .B2(new_n582), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n555), .A2(new_n658), .A3(new_n657), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n664), .A3(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT29), .B(new_n701), .C1(new_n745), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n739), .B1(new_n741), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n717), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(G13), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n208), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n711), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n212), .A2(new_n329), .ZN(new_n757));
  INV_X1    g0557(.A(G355), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n212), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n245), .A2(new_n271), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n212), .A2(new_n331), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n271), .B2(new_n715), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n215), .B1(G20), .B2(new_n397), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n756), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n209), .A2(new_n370), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n209), .A2(G179), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n320), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n774), .A2(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n320), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n209), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n779), .B1(G294), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n771), .A2(new_n320), .A3(G200), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT33), .B(G317), .Z(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n771), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n784), .A2(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n776), .A2(new_n786), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n329), .B(new_n789), .C1(G329), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n772), .A2(new_n363), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(G326), .B1(new_n795), .B2(G303), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n783), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n781), .A2(new_n488), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT32), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n774), .A2(new_n334), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n798), .B(new_n802), .C1(G50), .C2(new_n793), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n799), .ZN(new_n804));
  INV_X1    g0604(.A(new_n784), .ZN(new_n805));
  INV_X1    g0605(.A(new_n787), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n805), .A2(G68), .B1(new_n806), .B2(G77), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n777), .A2(new_n229), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n331), .B(new_n809), .C1(G87), .C2(new_n795), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT93), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n797), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n770), .B1(new_n812), .B2(new_n767), .ZN(new_n813));
  INV_X1    g0613(.A(new_n766), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n696), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n697), .B(KEYINPUT92), .ZN(new_n816));
  INV_X1    g0616(.A(new_n756), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n696), .B2(G330), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT94), .ZN(G396));
  AOI21_X1  g0620(.A(new_n743), .B1(new_n679), .B2(new_n625), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n701), .B1(new_n821), .B2(new_n671), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n441), .B(KEYINPUT95), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n438), .A2(new_n693), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n823), .A2(new_n437), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n631), .A2(new_n693), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n823), .A2(new_n437), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n701), .B(new_n830), .C1(new_n821), .C2(new_n671), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n829), .A2(new_n832), .A3(new_n738), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT96), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n738), .B1(new_n829), .B2(new_n832), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT97), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n756), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(new_n837), .C1(new_n836), .C2(new_n835), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n767), .A2(new_n764), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n756), .B1(G77), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G294), .ZN(new_n842));
  INV_X1    g0642(.A(new_n793), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n774), .A2(new_n842), .B1(new_n843), .B2(new_n476), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G107), .B2(new_n795), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n787), .A2(new_n490), .B1(new_n790), .B2(new_n788), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n329), .B(new_n846), .C1(G283), .C2(new_n805), .ZN(new_n847));
  INV_X1    g0647(.A(new_n777), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n798), .B1(G87), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n329), .B1(new_n790), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G68), .B2(new_n848), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n782), .A2(G58), .B1(new_n795), .B2(G50), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n805), .A2(G150), .B1(new_n806), .B2(G159), .ZN(new_n855));
  INV_X1    g0655(.A(G143), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n855), .B1(new_n774), .B2(new_n856), .C1(new_n857), .C2(new_n843), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n853), .B(new_n854), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n850), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n841), .B1(new_n862), .B2(new_n767), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n827), .B2(new_n765), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n838), .A2(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n753), .A2(new_n208), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n823), .A2(new_n693), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n831), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n267), .A2(new_n693), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n313), .A2(new_n365), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n362), .A2(new_n364), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n267), .B(new_n693), .C1(new_n634), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n356), .A2(new_n357), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT75), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n356), .A2(KEYINPUT75), .A3(new_n357), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n379), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n369), .A2(new_n691), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n691), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n377), .B1(new_n376), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n354), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n372), .A2(new_n691), .B1(new_n345), .B2(new_n353), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n326), .A2(new_n345), .A3(new_n353), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n882), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n882), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT18), .B1(new_n369), .B2(new_n372), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n376), .A2(new_n377), .A3(new_n374), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n875), .A2(new_n898), .B1(new_n901), .B2(new_n691), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n882), .B2(new_n893), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n895), .B(new_n892), .C1(new_n880), .C2(new_n881), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT39), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n881), .B1(new_n901), .B2(new_n876), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n884), .A2(new_n354), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n886), .B1(new_n889), .B2(KEYINPUT101), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n907), .A2(new_n908), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n895), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n897), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n905), .A2(KEYINPUT100), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n634), .A2(new_n267), .A3(new_n701), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT100), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(KEYINPUT39), .C1(new_n903), .C2(new_n904), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n902), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n741), .A2(new_n749), .A3(new_n454), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n639), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(G330), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n897), .A2(new_n912), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n873), .A2(new_n737), .A3(new_n827), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n870), .A2(new_n872), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n737), .A2(new_n827), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT102), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT102), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n873), .A2(new_n933), .A3(new_n737), .A4(new_n827), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n898), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n454), .A2(new_n737), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n925), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n866), .B1(new_n924), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n924), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n217), .A2(new_n490), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(KEYINPUT35), .B2(new_n573), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT98), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT36), .Z(new_n949));
  NOR3_X1   g0749(.A1(new_n219), .A2(new_n227), .A3(new_n335), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n221), .A2(G50), .ZN(new_n951));
  OAI211_X1 g0751(.A(G1), .B(new_n752), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n942), .A2(new_n949), .A3(new_n952), .ZN(G367));
  OAI221_X1 g0753(.A(new_n768), .B1(new_n212), .B2(new_n430), .C1(new_n241), .C2(new_n761), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(new_n756), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n656), .B1(new_n654), .B2(new_n701), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n664), .A2(new_n654), .A3(new_n701), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n787), .A2(new_n202), .B1(new_n790), .B2(new_n857), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n331), .B(new_n959), .C1(G159), .C2(new_n805), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n795), .A2(G58), .B1(new_n848), .B2(G77), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G68), .A2(new_n782), .B1(new_n793), .B2(G143), .ZN(new_n962));
  INV_X1    g0762(.A(G150), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(new_n774), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT107), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n960), .B(new_n961), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n777), .A2(new_n488), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G311), .B2(new_n793), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n229), .B2(new_n781), .C1(new_n476), .C2(new_n774), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n805), .A2(G294), .B1(new_n791), .B2(G317), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT46), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n794), .B2(new_n490), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n795), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n329), .B1(new_n806), .B2(G283), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n973), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n966), .A2(new_n967), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT47), .Z(new_n978));
  INV_X1    g0778(.A(new_n767), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n955), .B1(new_n958), .B2(new_n814), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n710), .B(KEYINPUT41), .ZN(new_n981));
  INV_X1    g0781(.A(new_n703), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n580), .A2(new_n693), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n742), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n582), .B2(new_n701), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n708), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n708), .A2(new_n985), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(KEYINPUT104), .B(new_n982), .C1(new_n989), .C2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n697), .ZN(new_n996));
  INV_X1    g0796(.A(new_n706), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(KEYINPUT105), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n997), .A2(KEYINPUT105), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n702), .A2(new_n705), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  MUX2_X1   g0801(.A(new_n996), .B(new_n816), .S(new_n1001), .Z(new_n1002));
  AOI22_X1  g0802(.A1(new_n987), .A2(new_n988), .B1(new_n993), .B2(new_n992), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT104), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n703), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n995), .A2(new_n1002), .A3(new_n1005), .A4(new_n750), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n981), .B1(new_n1006), .B2(new_n750), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n754), .B(KEYINPUT106), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n982), .A2(new_n985), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n706), .A2(new_n985), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT103), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT42), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n582), .B1(new_n984), .B2(new_n625), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1013), .A2(KEYINPUT42), .B1(new_n701), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1014), .A2(new_n1016), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1011), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1021), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1023), .A2(new_n1019), .A3(new_n1010), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n980), .B1(new_n1009), .B2(new_n1025), .ZN(G387));
  OR2_X1    g0826(.A1(new_n702), .A2(new_n814), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n713), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1028), .A2(new_n757), .B1(G107), .B2(new_n212), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n428), .A2(new_n202), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI21_X1  g0833(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1032), .A2(new_n1028), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n761), .B1(new_n238), .B2(G45), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1029), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n756), .B1(new_n1037), .B2(new_n769), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n348), .A2(new_n805), .B1(new_n806), .B2(G68), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT109), .Z(new_n1040));
  AOI211_X1 g0840(.A(new_n331), .B(new_n968), .C1(G150), .C2(new_n791), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n781), .A2(new_n430), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G50), .B2(new_n773), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n793), .A2(G159), .B1(new_n795), .B2(G77), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n329), .B1(new_n791), .B2(G326), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n781), .A2(new_n778), .B1(new_n794), .B2(new_n842), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n805), .A2(G311), .B1(new_n806), .B2(G303), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n773), .A2(G317), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n775), .C2(new_n843), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1046), .B1(new_n490), .B2(new_n777), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1045), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1038), .B1(new_n1057), .B2(new_n767), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1002), .A2(new_n1008), .B1(new_n1027), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1002), .A2(new_n750), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n711), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1002), .A2(new_n750), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  AND2_X1   g0863(.A1(new_n1002), .A2(new_n750), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1003), .B(new_n982), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1006), .B(new_n711), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n985), .A2(new_n814), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n768), .B1(new_n488), .B2(new_n212), .C1(new_n248), .C2(new_n761), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n756), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G150), .A2(new_n793), .B1(new_n773), .B2(G159), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  AOI22_X1  g0871(.A1(new_n428), .A2(new_n806), .B1(G50), .B2(new_n805), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT110), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n781), .A2(new_n227), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n329), .B1(new_n790), .B2(new_n856), .C1(new_n223), .C2(new_n777), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(G68), .C2(new_n795), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1071), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G311), .A2(new_n773), .B1(new_n793), .B2(G317), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT52), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n787), .A2(new_n842), .B1(new_n790), .B2(new_n775), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n329), .B(new_n1080), .C1(G303), .C2(new_n805), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n794), .A2(new_n778), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n809), .B(new_n1082), .C1(G116), .C2(new_n782), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1069), .B1(new_n1085), .B2(new_n767), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1065), .A2(new_n1008), .B1(new_n1067), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1066), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(KEYINPUT111), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT111), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1066), .A2(new_n1090), .A3(new_n1087), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(G390));
  INV_X1    g0892(.A(KEYINPUT114), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n701), .B(new_n830), .C1(new_n745), .C2(new_n748), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n867), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n737), .A2(G330), .A3(new_n827), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1095), .B1(new_n1097), .B2(new_n873), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n737), .A2(KEYINPUT113), .A3(G330), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT113), .B1(new_n737), .B2(G330), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n828), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1098), .B1(new_n1101), .B2(new_n873), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1096), .A2(new_n930), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n873), .A2(G330), .A3(new_n737), .A4(new_n827), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT112), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1096), .A2(new_n930), .A3(KEYINPUT112), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n868), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n739), .A2(new_n454), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n922), .A2(new_n639), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1093), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(KEYINPUT114), .B(new_n1111), .C1(new_n1102), .C2(new_n1108), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n915), .A2(new_n919), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n874), .A2(new_n916), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1094), .A2(new_n867), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n916), .B(new_n926), .C1(new_n1119), .C2(new_n930), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n1104), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1104), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n915), .A2(new_n919), .B1(new_n874), .B2(new_n916), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1120), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n710), .B1(new_n1115), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1126), .B2(new_n1115), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1121), .A2(new_n1125), .A3(new_n1008), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n756), .B1(new_n348), .B2(new_n840), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n793), .A2(G128), .B1(new_n848), .B2(G50), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n851), .B2(new_n774), .C1(new_n800), .C2(new_n781), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n805), .A2(G137), .B1(new_n806), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n795), .A2(new_n1136), .A3(G150), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n794), .B2(new_n963), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n331), .B1(new_n791), .B2(G125), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1135), .A2(new_n1137), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1074), .B1(G116), .B2(new_n773), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n778), .B2(new_n843), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n795), .A2(G87), .B1(new_n848), .B2(G68), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G97), .A2(new_n806), .B1(new_n791), .B2(G294), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n329), .B1(new_n805), .B2(G107), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1132), .A2(new_n1141), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT116), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n979), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1130), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1116), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n765), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1128), .A2(new_n1129), .A3(new_n1154), .ZN(G378));
  INV_X1    g0955(.A(new_n921), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n928), .A2(KEYINPUT102), .B1(new_n897), .B2(new_n896), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT40), .B1(new_n1157), .B2(new_n934), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT55), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n415), .B2(new_n883), .ZN(new_n1162));
  AOI211_X1 g0962(.A(KEYINPUT55), .B(new_n691), .C1(new_n404), .C2(new_n408), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n451), .A2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n448), .B(new_n1164), .C1(new_n450), .C2(new_n413), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n419), .A2(new_n1164), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n451), .A2(new_n1165), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n1170), .A3(new_n1159), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT118), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1168), .A2(KEYINPUT118), .A3(new_n1171), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(KEYINPUT119), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1158), .A2(new_n1174), .A3(new_n925), .A4(new_n929), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1168), .A2(KEYINPUT119), .A3(new_n1171), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n937), .B2(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1156), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1174), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n937), .A2(new_n1179), .A3(G330), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1158), .A2(new_n925), .A3(new_n929), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n921), .C1(new_n1181), .C2(new_n1176), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1109), .A2(new_n1093), .A3(new_n1112), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1106), .A2(new_n868), .A3(new_n1107), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1119), .A2(new_n1104), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1100), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n737), .A2(KEYINPUT113), .A3(G330), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n827), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1186), .B1(new_n1189), .B2(new_n930), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1112), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT114), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1126), .B1(new_n1184), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1193), .B2(new_n1111), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n710), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1183), .B(KEYINPUT57), .C1(new_n1193), .C2(new_n1111), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT120), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1112), .B1(new_n1115), .B2(new_n1126), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT120), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT57), .A4(new_n1183), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1196), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n784), .A2(new_n851), .B1(new_n787), .B2(new_n857), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G150), .A2(new_n782), .B1(new_n793), .B2(G125), .ZN(new_n1204));
  INV_X1    g1004(.A(G128), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n774), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1203), .B(new_n1206), .C1(new_n795), .C2(new_n1134), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n848), .A2(G159), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n331), .B2(new_n270), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n774), .A2(new_n229), .B1(new_n777), .B2(new_n334), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G116), .B2(new_n793), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G41), .B(new_n329), .C1(new_n805), .C2(G97), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n550), .A2(new_n806), .B1(new_n791), .B2(G283), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n782), .A2(G68), .B1(new_n795), .B2(G77), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1215), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1213), .B(new_n1223), .C1(new_n1222), .C2(new_n1221), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n767), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n756), .C1(G50), .C2(new_n840), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1173), .A2(new_n1172), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n764), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1183), .B2(new_n1008), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1202), .A2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1109), .A2(new_n1008), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n930), .A2(new_n764), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT122), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n817), .B1(new_n221), .B2(new_n839), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1042), .B1(G283), .B2(new_n773), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT123), .Z(new_n1236));
  AOI22_X1  g1036(.A1(new_n795), .A2(G97), .B1(new_n848), .B2(G77), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n842), .B2(new_n843), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n331), .B1(new_n784), .B2(new_n490), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n787), .A2(new_n229), .B1(new_n790), .B2(new_n476), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n774), .A2(new_n857), .B1(new_n202), .B2(new_n781), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G159), .B2(new_n795), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n843), .A2(new_n851), .B1(new_n777), .B2(new_n334), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n329), .B1(new_n784), .B2(new_n1133), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n787), .A2(new_n963), .B1(new_n790), .B2(new_n1205), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1236), .A2(new_n1241), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1233), .B(new_n1234), .C1(new_n979), .C2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1231), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n981), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1115), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1102), .A2(new_n1111), .A3(new_n1108), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT121), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1102), .A2(new_n1108), .A3(KEYINPUT121), .A4(new_n1111), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1251), .B1(new_n1253), .B2(new_n1258), .ZN(G381));
  NOR2_X1   g1059(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1089), .A2(new_n1261), .A3(new_n980), .A4(new_n1091), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1262), .A2(G384), .A3(G381), .A4(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(G375), .A2(G378), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(G407));
  NAND2_X1  g1067(.A1(new_n692), .A2(G213), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1270), .ZN(G409));
  NAND3_X1  g1071(.A1(new_n1202), .A2(G378), .A3(new_n1229), .ZN(new_n1272));
  INV_X1    g1072(.A(G378), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1229), .A2(KEYINPUT124), .B1(new_n1194), .B2(new_n981), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1229), .A2(KEYINPUT124), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1268), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1269), .A2(G2897), .ZN(new_n1279));
  INV_X1    g1079(.A(G384), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n711), .B1(new_n1254), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1192), .A2(KEYINPUT60), .A3(new_n1184), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1280), .B1(new_n1285), .B2(new_n1250), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1258), .B1(new_n1115), .B2(KEYINPUT60), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G384), .B(new_n1251), .C1(new_n1287), .C2(new_n1282), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1279), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n1288), .A3(KEYINPUT125), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1289), .B1(new_n1293), .B2(new_n1279), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1277), .A2(new_n1268), .A3(new_n1293), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G393), .A2(G396), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1264), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G390), .A2(G387), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n1299), .B(new_n1301), .C1(new_n1302), .C2(new_n1262), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1300), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1300), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1299), .B1(new_n1305), .B2(new_n1263), .ZN(new_n1306));
  AND4_X1   g1106(.A1(new_n1262), .A2(new_n1302), .A3(new_n1304), .A4(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1269), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1293), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1295), .A2(new_n1298), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1286), .A2(new_n1288), .A3(KEYINPUT125), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1279), .B1(new_n1313), .B2(new_n1290), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1289), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1312), .B1(new_n1309), .B2(new_n1316), .ZN(new_n1317));
  XOR2_X1   g1117(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1318));
  NAND2_X1  g1118(.A1(new_n1296), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1309), .A2(KEYINPUT62), .A3(new_n1293), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1311), .B1(new_n1321), .B2(new_n1308), .ZN(G405));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1273), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1272), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1293), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1323), .A2(new_n1326), .A3(new_n1272), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1302), .A2(new_n1262), .A3(new_n1306), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1304), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1329), .B(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1328), .B(new_n1331), .ZN(G402));
endmodule


