//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(G224), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT7), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n188), .ZN(new_n191));
  XNOR2_X1  g005(.A(G143), .B(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT0), .B(G128), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n195), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n205), .B1(new_n192), .B2(new_n201), .ZN(new_n206));
  AND4_X1   g020(.A1(new_n205), .A2(new_n197), .A3(new_n199), .A4(new_n201), .ZN(new_n207));
  OAI22_X1  g021(.A1(new_n194), .A2(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n200), .A2(new_n210), .A3(G128), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n197), .B(new_n199), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(G125), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n191), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT64), .B1(new_n192), .B2(new_n193), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n203), .A3(new_n195), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n197), .A2(new_n199), .A3(new_n201), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n192), .A2(new_n205), .A3(new_n201), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n217), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n225), .A2(new_n188), .A3(new_n214), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n190), .B1(new_n216), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n209), .A2(new_n215), .ZN(new_n228));
  XNOR2_X1  g042(.A(G110), .B(G122), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n229), .B(KEYINPUT8), .ZN(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n233), .A2(KEYINPUT5), .A3(G119), .ZN(new_n234));
  INV_X1    g048(.A(G113), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT2), .A2(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT2), .A2(G113), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n237), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n232), .A2(new_n236), .B1(new_n242), .B2(new_n231), .ZN(new_n243));
  INV_X1    g057(.A(G104), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT3), .B1(new_n244), .B2(G107), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n246));
  INV_X1    g060(.A(G107), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G104), .ZN(new_n248));
  INV_X1    g062(.A(G101), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(G107), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n245), .A2(new_n248), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n244), .A2(G107), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n247), .A2(G104), .ZN(new_n253));
  OAI21_X1  g067(.A(G101), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n254), .A3(KEYINPUT85), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n230), .B1(new_n243), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n254), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT85), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n243), .A3(new_n255), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n228), .A2(new_n189), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n227), .A2(KEYINPUT86), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n188), .B1(new_n225), .B2(new_n214), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n218), .A2(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n215), .B(new_n191), .C1(new_n266), .C2(new_n217), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n189), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n214), .B1(new_n208), .B2(G125), .ZN(new_n269));
  INV_X1    g083(.A(new_n261), .ZN(new_n270));
  OAI22_X1  g084(.A1(new_n269), .A2(new_n190), .B1(new_n270), .B2(new_n256), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n264), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n245), .A2(new_n248), .A3(new_n250), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G101), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT4), .A3(new_n251), .ZN(new_n275));
  INV_X1    g089(.A(new_n231), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n242), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n242), .A2(new_n276), .A3(new_n277), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n282), .A3(G101), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n275), .A2(new_n280), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n251), .A2(new_n254), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n251), .B2(new_n254), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n243), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n288), .A3(new_n229), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n263), .A2(new_n272), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n265), .A2(new_n267), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n284), .A2(new_n288), .A3(KEYINPUT82), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT82), .B1(new_n284), .B2(new_n288), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(new_n229), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n289), .A2(KEYINPUT6), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT83), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n284), .A2(new_n288), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n284), .A2(new_n288), .A3(KEYINPUT82), .ZN(new_n302));
  INV_X1    g116(.A(new_n229), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n305));
  INV_X1    g119(.A(new_n297), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT6), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n301), .A2(new_n308), .A3(new_n302), .A4(new_n303), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT84), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n295), .A2(new_n229), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT84), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n311), .A2(new_n312), .A3(new_n308), .A4(new_n302), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n298), .A2(new_n307), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n292), .B1(new_n293), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G210), .B1(G237), .B2(G902), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT87), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n310), .A2(new_n313), .ZN(new_n318));
  INV_X1    g132(.A(new_n307), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n305), .B1(new_n304), .B2(new_n306), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n318), .B(new_n293), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n289), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n268), .A2(new_n271), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(KEYINPUT86), .ZN(new_n324));
  AOI21_X1  g138(.A(G902), .B1(new_n324), .B2(new_n272), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n325), .A3(new_n316), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n321), .A2(new_n325), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n328));
  INV_X1    g142(.A(new_n316), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT9), .B(G234), .ZN(new_n332));
  OAI21_X1  g146(.A(G221), .B1(new_n332), .B2(G902), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT78), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT79), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n211), .A2(new_n213), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n258), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(G137), .ZN(new_n341));
  INV_X1    g155(.A(G137), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT11), .A3(G134), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(G137), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G131), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n347));
  INV_X1    g161(.A(G131), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n341), .A2(new_n343), .A3(new_n348), .A4(new_n344), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n345), .A2(KEYINPUT66), .A3(G131), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n338), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT12), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n338), .A2(new_n353), .A3(KEYINPUT12), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G140), .ZN(new_n359));
  INV_X1    g173(.A(G953), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n360), .A2(G227), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n359), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n266), .A2(new_n283), .A3(new_n275), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n286), .B2(new_n287), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n337), .B2(new_n258), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n364), .A2(new_n366), .A3(new_n352), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n369), .A2(new_n370), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n358), .B(new_n363), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n364), .A2(new_n368), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(KEYINPUT81), .A3(new_n352), .A4(new_n366), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n369), .A2(new_n370), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n375), .A2(new_n376), .B1(new_n353), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n378), .B2(new_n363), .ZN(new_n379));
  INV_X1    g193(.A(G469), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n379), .A2(new_n380), .A3(new_n291), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n353), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n363), .C1(new_n371), .C2(new_n372), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n375), .A2(new_n376), .B1(new_n357), .B2(new_n356), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n383), .B(G469), .C1(new_n384), .C2(new_n363), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(new_n291), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n336), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(G475), .A2(G902), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(G237), .A2(G953), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n393), .A2(G143), .A3(G214), .ZN(new_n394));
  AOI21_X1  g208(.A(G143), .B1(new_n393), .B2(G214), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(G214), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n198), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(G143), .A3(G214), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n348), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n217), .A2(KEYINPUT16), .A3(G140), .ZN(new_n402));
  XNOR2_X1  g216(.A(G125), .B(G140), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G146), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT19), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n403), .B(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n401), .B(new_n405), .C1(G146), .C2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n394), .A2(new_n395), .ZN(new_n409));
  NAND2_X1  g223(.A1(KEYINPUT18), .A2(G131), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n196), .ZN(new_n411));
  INV_X1    g225(.A(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n217), .A2(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G146), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n409), .A2(new_n410), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT18), .B(G131), .C1(new_n394), .C2(new_n395), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n408), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G113), .B(G122), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(new_n244), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n401), .A2(KEYINPUT17), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n196), .B1(new_n427), .B2(new_n402), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT17), .B(G131), .C1(new_n394), .C2(new_n395), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n405), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n419), .B(new_n422), .C1(new_n425), .C2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n392), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n433));
  INV_X1    g247(.A(new_n431), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n422), .B1(new_n408), .B2(new_n419), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n424), .A2(KEYINPUT88), .A3(new_n431), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n390), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n432), .B1(new_n438), .B2(KEYINPUT20), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(G902), .A3(G953), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G898), .ZN(new_n443));
  INV_X1    g257(.A(G952), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(G953), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n442), .A2(new_n443), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G475), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n419), .B1(new_n425), .B2(new_n430), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n423), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n431), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n450), .B2(new_n291), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n439), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G478), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n454));
  INV_X1    g268(.A(G217), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n332), .A2(new_n455), .A3(G953), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT89), .B1(new_n458), .B2(G116), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n233), .A3(G122), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT14), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(G116), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n459), .A2(new_n461), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT93), .B1(new_n466), .B2(KEYINPUT14), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n468), .B(new_n462), .C1(new_n459), .C2(new_n461), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G107), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n198), .A2(G128), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n212), .A2(G143), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G134), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n340), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n466), .A2(new_n247), .A3(new_n464), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n466), .A2(new_n247), .A3(new_n464), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n247), .B1(new_n466), .B2(new_n464), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n476), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT13), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(new_n487), .C1(new_n212), .C2(G143), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n473), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT13), .B1(new_n198), .B2(G128), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n486), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n198), .A2(KEYINPUT13), .A3(G128), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n487), .B1(new_n212), .B2(G143), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT90), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(KEYINPUT91), .A3(new_n473), .A4(new_n488), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n484), .B1(G134), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n481), .B1(new_n498), .B2(KEYINPUT92), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n493), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n488), .A2(new_n473), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT91), .B1(new_n501), .B2(new_n495), .ZN(new_n502));
  OAI21_X1  g316(.A(G134), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n476), .ZN(new_n504));
  INV_X1    g318(.A(new_n483), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(new_n478), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT92), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n457), .B1(new_n499), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n479), .B1(new_n470), .B2(G107), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n498), .A2(KEYINPUT92), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n456), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT94), .B1(new_n515), .B2(new_n291), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n517), .B(G902), .C1(new_n510), .C2(new_n514), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n454), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n499), .A2(new_n509), .A3(new_n457), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n456), .B1(new_n512), .B2(new_n513), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n291), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n454), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n452), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n389), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(G214), .B1(G237), .B2(G902), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n331), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n455), .B1(G234), .B2(new_n291), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G119), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G128), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n212), .A2(G119), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT72), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT72), .B1(new_n534), .B2(new_n535), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT24), .B(G110), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT73), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n533), .A2(G128), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT74), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT23), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(KEYINPUT74), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n534), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n428), .A2(new_n405), .B1(new_n546), .B2(G110), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n411), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n404), .B2(G146), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT75), .B(G110), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n543), .A2(new_n534), .A3(new_n545), .A4(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT24), .B(G110), .Z(new_n553));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n212), .A2(G119), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n541), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT72), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n552), .B1(new_n558), .B2(KEYINPUT76), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT76), .B(new_n538), .C1(new_n536), .C2(new_n537), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT77), .B(new_n550), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n538), .B1(new_n536), .B2(new_n537), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n560), .A3(new_n552), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT77), .B1(new_n567), .B2(new_n550), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n548), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n360), .A2(G221), .A3(G234), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n548), .B(new_n572), .C1(new_n563), .C2(new_n568), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n291), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT25), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n574), .A2(KEYINPUT25), .A3(new_n291), .A4(new_n575), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n532), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n531), .A2(G902), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n575), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(G472), .A2(G902), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n350), .A2(new_n220), .A3(new_n351), .A4(new_n224), .ZN(new_n587));
  INV_X1    g401(.A(new_n337), .ZN(new_n588));
  INV_X1    g402(.A(new_n344), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n340), .A2(G137), .ZN(new_n590));
  OAI21_X1  g404(.A(G131), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n349), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT30), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n280), .A2(new_n281), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n592), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n587), .A2(KEYINPUT67), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT67), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n266), .A2(new_n599), .A3(new_n351), .A4(new_n350), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n594), .B(new_n596), .C1(new_n601), .C2(KEYINPUT30), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n393), .A2(G210), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(KEYINPUT27), .Z(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT26), .B(G101), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n593), .B2(new_n595), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT31), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n602), .B2(new_n607), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n593), .A2(new_n595), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n601), .B2(new_n595), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT28), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n587), .A2(new_n592), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n616), .A2(KEYINPUT71), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n596), .B1(new_n616), .B2(KEYINPUT71), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT28), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n606), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n586), .B1(new_n612), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n606), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n602), .A2(new_n613), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n606), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT29), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT28), .B1(new_n617), .B2(new_n618), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n616), .A2(new_n596), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n620), .B1(new_n613), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n606), .A2(new_n629), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(KEYINPUT32), .A2(new_n624), .B1(new_n637), .B2(G472), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT32), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n625), .B1(new_n615), .B2(new_n621), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n640), .A2(new_n609), .A3(new_n611), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n639), .B1(new_n641), .B2(new_n586), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n584), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n331), .A2(new_n526), .A3(KEYINPUT95), .A4(new_n527), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n530), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  INV_X1    g460(.A(new_n527), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n327), .A2(new_n329), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(new_n326), .ZN(new_n649));
  INV_X1    g463(.A(new_n446), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n439), .A2(new_n451), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n515), .A2(KEYINPUT33), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n515), .A2(KEYINPUT33), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(G478), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n453), .A2(new_n291), .ZN(new_n655));
  AOI21_X1  g469(.A(G902), .B1(new_n510), .B2(new_n514), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n453), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n649), .A2(new_n650), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n612), .A2(new_n623), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n585), .ZN(new_n662));
  INV_X1    g476(.A(G472), .ZN(new_n663));
  AOI21_X1  g477(.A(G902), .B1(new_n612), .B2(new_n623), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n584), .A3(new_n389), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NAND2_X1  g483(.A1(new_n519), .A2(new_n524), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n438), .A2(KEYINPUT20), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n436), .A2(new_n391), .A3(new_n437), .A4(new_n390), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n451), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(new_n649), .A3(new_n650), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n666), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT96), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  OR2_X1    g493(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n569), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n569), .A2(new_n680), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n681), .A2(new_n582), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n578), .A2(new_n579), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n683), .B1(new_n684), .B2(new_n531), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n665), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n530), .A2(new_n644), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  AOI21_X1  g503(.A(new_n685), .B1(new_n638), .B2(new_n642), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n445), .A2(new_n440), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT97), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(new_n442), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n451), .B(new_n695), .C1(new_n671), .C2(new_n672), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n697));
  INV_X1    g511(.A(new_n454), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n522), .A2(new_n517), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n656), .A2(KEYINPUT94), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n696), .B(new_n697), .C1(new_n701), .C2(new_n523), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n697), .B1(new_n670), .B2(new_n696), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n385), .A2(new_n387), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n379), .A2(new_n380), .A3(new_n291), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n335), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n690), .A2(new_n705), .A3(new_n708), .A4(new_n649), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XOR2_X1   g524(.A(new_n695), .B(KEYINPUT39), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(KEYINPUT40), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n627), .A2(new_n625), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n613), .A2(new_n632), .ZN(new_n715));
  AOI21_X1  g529(.A(G902), .B1(new_n715), .B2(new_n606), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n663), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n662), .B2(new_n639), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n624), .A2(KEYINPUT32), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n699), .A2(new_n700), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n523), .B1(new_n721), .B2(new_n454), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n439), .A2(new_n451), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n685), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n647), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n713), .A2(new_n720), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n331), .B(KEYINPUT38), .Z(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n198), .ZN(G45));
  NOR2_X1   g544(.A1(new_n658), .A2(new_n695), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n690), .A2(new_n708), .A3(new_n649), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  OAI21_X1  g547(.A(new_n382), .B1(new_n371), .B2(new_n372), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n362), .B1(new_n375), .B2(new_n376), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n734), .A2(new_n362), .B1(new_n735), .B2(new_n358), .ZN(new_n736));
  OAI21_X1  g550(.A(G469), .B1(new_n736), .B2(G902), .ZN(new_n737));
  INV_X1    g551(.A(new_n334), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n707), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT99), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT99), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n737), .A2(new_n741), .A3(new_n738), .A4(new_n707), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n660), .A2(new_n643), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND3_X1  g560(.A1(new_n675), .A2(new_n643), .A3(new_n743), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT100), .B(G116), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G18));
  AND3_X1   g563(.A1(new_n649), .A2(new_n740), .A3(new_n742), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n722), .A3(new_n452), .A4(new_n690), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  XNOR2_X1  g566(.A(new_n584), .B(KEYINPUT103), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT104), .B1(new_n722), .B2(new_n723), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n670), .A2(new_n755), .A3(new_n651), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n754), .A2(new_n650), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT101), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n634), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT101), .B1(new_n631), .B2(new_n633), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n606), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n586), .B1(new_n761), .B2(new_n612), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n664), .B2(new_n663), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT102), .B(G472), .C1(new_n641), .C2(G902), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n753), .A2(new_n757), .A3(new_n750), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  AOI211_X1 g582(.A(new_n685), .B(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n750), .A3(new_n731), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n642), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n662), .A2(KEYINPUT106), .A3(new_n639), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n638), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n753), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n647), .B1(new_n315), .B2(new_n316), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n334), .B1(new_n706), .B2(new_n707), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n317), .A2(new_n778), .A3(new_n779), .A4(new_n330), .ZN(new_n780));
  INV_X1    g594(.A(new_n731), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n780), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n643), .A3(new_n731), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n782), .B1(new_n786), .B2(KEYINPUT105), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n637), .A2(G472), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n719), .A2(new_n642), .A3(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n581), .A2(new_n583), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n781), .A3(new_n780), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT105), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n784), .B1(new_n787), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G131), .ZN(G33));
  INV_X1    g610(.A(KEYINPUT107), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n705), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT107), .B1(new_n703), .B2(new_n704), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n643), .A3(new_n785), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G134), .ZN(G36));
  OAI21_X1  g615(.A(new_n383), .B1(new_n384), .B2(new_n363), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(G469), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n804), .A2(KEYINPUT108), .A3(G469), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT46), .B1(new_n810), .B2(new_n387), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n381), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(KEYINPUT46), .A3(new_n387), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n334), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n711), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n665), .A2(new_n725), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n654), .A2(new_n723), .A3(new_n657), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT43), .Z(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(KEYINPUT44), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n317), .A2(new_n330), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(new_n778), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT44), .B1(new_n818), .B2(new_n820), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n815), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(new_n342), .ZN(G39));
  INV_X1    g641(.A(new_n823), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n828), .A2(new_n789), .A3(new_n790), .A4(new_n781), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n814), .A2(KEYINPUT47), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n814), .A2(KEYINPUT47), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(new_n412), .ZN(G42));
  AND2_X1   g648(.A1(new_n737), .A2(new_n707), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT49), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n819), .A2(new_n647), .A3(new_n335), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n753), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n728), .A2(new_n838), .A3(new_n719), .A4(new_n718), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n754), .A2(new_n649), .A3(new_n756), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n707), .A2(new_n387), .A3(new_n385), .ZN(new_n842));
  INV_X1    g656(.A(new_n695), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n685), .A2(new_n842), .A3(new_n738), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n719), .B2(new_n718), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n754), .A2(new_n649), .A3(new_n756), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n580), .A2(new_n683), .A3(new_n695), .ZN(new_n849));
  INV_X1    g663(.A(new_n717), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n624), .B2(KEYINPUT32), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n641), .A2(new_n639), .A3(new_n586), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n779), .B(new_n849), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT112), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n770), .A2(new_n709), .A3(new_n732), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n840), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n847), .A2(new_n854), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n789), .A2(new_n708), .A3(new_n725), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n649), .C1(new_n705), .C2(new_n731), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n858), .A2(new_n861), .A3(KEYINPUT52), .A4(new_n770), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n643), .B(new_n743), .C1(new_n675), .C2(new_n660), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n767), .A3(new_n751), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n792), .A2(new_n793), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n786), .A2(KEYINPUT105), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n782), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n865), .B1(new_n868), .B2(new_n784), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n658), .A2(new_n446), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n331), .A2(new_n527), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT110), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT110), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n331), .A2(new_n873), .A3(new_n870), .A4(new_n527), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n666), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n331), .A2(new_n527), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n670), .A2(new_n723), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT111), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n878), .A3(new_n650), .A4(new_n666), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n645), .A2(new_n687), .A3(new_n875), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n860), .A2(new_n823), .A3(new_n722), .A4(new_n696), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n769), .A2(new_n731), .A3(new_n785), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n800), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n863), .A2(new_n869), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(KEYINPUT53), .B2(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n884), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n767), .A2(new_n751), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n795), .A2(new_n864), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT115), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT115), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n869), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n885), .A2(new_n899), .A3(new_n886), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n885), .B2(new_n886), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n891), .B(new_n898), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n728), .A2(new_n647), .A3(new_n743), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n820), .A2(new_n693), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n753), .A3(new_n766), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n904), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT50), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n823), .A2(new_n743), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(new_n906), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n720), .A2(new_n584), .A3(new_n691), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n651), .B1(new_n654), .B2(new_n657), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n769), .A2(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n835), .A2(new_n335), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n831), .A2(new_n832), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n907), .A2(new_n828), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n908), .A2(new_n909), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n914), .A2(new_n659), .ZN(new_n927));
  INV_X1    g741(.A(new_n750), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n927), .B(new_n445), .C1(new_n928), .C2(new_n907), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n912), .A2(new_n777), .ZN(new_n930));
  NOR2_X1   g744(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n931));
  AND2_X1   g745(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n929), .B(new_n933), .C1(new_n930), .C2(new_n932), .ZN(new_n934));
  AND4_X1   g748(.A1(new_n903), .A2(new_n925), .A3(new_n926), .A4(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(G952), .A2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n839), .B1(new_n935), .B2(new_n936), .ZN(G75));
  NOR2_X1   g751(.A1(new_n360), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(G210), .A3(G902), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT119), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n314), .B(new_n293), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT56), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n942), .B1(new_n941), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n939), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n885), .A2(new_n886), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT114), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n885), .A2(new_n899), .A3(new_n886), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n895), .A2(new_n897), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n951), .A2(new_n952), .B1(new_n892), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n291), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(KEYINPUT118), .A3(G210), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT56), .B1(new_n941), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n944), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n949), .A2(new_n959), .ZN(G51));
  NAND2_X1  g774(.A1(new_n951), .A2(new_n952), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n891), .B1(new_n961), .B2(new_n898), .ZN(new_n962));
  INV_X1    g776(.A(new_n902), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n386), .B(KEYINPUT57), .Z(new_n965));
  OAI21_X1  g779(.A(new_n379), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n810), .B(KEYINPUT120), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n955), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n938), .B1(new_n966), .B2(new_n968), .ZN(G54));
  NAND3_X1  g783(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n436), .A2(new_n437), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n938), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .A4(new_n971), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(G60));
  AND2_X1   g789(.A1(new_n652), .A2(new_n653), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n655), .B(KEYINPUT59), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n962), .B2(new_n963), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(KEYINPUT121), .A3(new_n939), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT121), .ZN(new_n981));
  INV_X1    g795(.A(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n940), .A2(KEYINPUT54), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n902), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n984), .B2(new_n938), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n976), .B1(new_n903), .B2(new_n977), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n980), .A2(new_n985), .A3(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(new_n574), .A2(new_n575), .ZN(new_n988));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT60), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n954), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n940), .A2(new_n681), .A3(new_n682), .A4(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n939), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT122), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n940), .A2(new_n992), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n938), .B1(new_n1000), .B2(new_n988), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n996), .A3(new_n997), .A4(new_n993), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n999), .A2(new_n1002), .ZN(G66));
  NOR2_X1   g817(.A1(new_n880), .A2(new_n865), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1004), .A2(G953), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n443), .B2(new_n187), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n314), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(G898), .B2(new_n360), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1008), .B(new_n1010), .ZN(G69));
  OAI21_X1  g825(.A(new_n594), .B1(new_n601), .B2(KEYINPUT30), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT124), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(new_n407), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n833), .A2(new_n826), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n814), .A2(new_n711), .A3(new_n777), .A4(new_n841), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n861), .A2(new_n770), .A3(new_n800), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1016), .A2(new_n795), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(G953), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT125), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n360), .A2(G900), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(KEYINPUT125), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1014), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n360), .B1(G227), .B2(G900), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1014), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n729), .A2(KEYINPUT62), .A3(new_n856), .ZN(new_n1029));
  OR2_X1    g843(.A1(new_n878), .A2(new_n659), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n828), .A2(new_n791), .A3(new_n712), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(KEYINPUT62), .B1(new_n729), .B2(new_n856), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1015), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1028), .B1(new_n1034), .B2(new_n360), .ZN(new_n1035));
  OR3_X1    g849(.A1(new_n1026), .A2(new_n1027), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1027), .B1(new_n1026), .B2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(G72));
  INV_X1    g852(.A(new_n1004), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT126), .ZN(new_n1041));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  AND3_X1   g857(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1041), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n1044), .A2(new_n1045), .A3(new_n714), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n627), .A2(new_n625), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1015), .A2(new_n1004), .A3(new_n1018), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n1043), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1048), .B1(new_n1050), .B2(KEYINPUT127), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1051), .B1(KEYINPUT127), .B2(new_n1050), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n889), .A2(new_n714), .A3(new_n1043), .A4(new_n1048), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1052), .A2(new_n939), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1046), .A2(new_n1054), .ZN(G57));
endmodule


