//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G221), .A2(G219), .A3(G218), .A4(G220), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT69), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(new_n456), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT71), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n470), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  AND4_X1   g056(.A1(new_n467), .A2(new_n471), .A3(new_n472), .A4(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n477), .A2(new_n470), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n470), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n483), .A2(G124), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OR3_X1    g062(.A1(new_n477), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n468), .A2(new_n470), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT72), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G136), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n474), .A2(new_n476), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT73), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n468), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n474), .A2(new_n476), .A3(G138), .A4(new_n470), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n506), .A2(new_n470), .A3(G114), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT74), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .A4(new_n470), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n500), .A2(new_n503), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(new_n517), .B1(G75), .B2(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n515), .A2(KEYINPUT75), .A3(G62), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(new_n515), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI21_X1  g101(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n520), .A2(new_n528), .ZN(G166));
  XOR2_X1   g104(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(new_n531), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n527), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT5), .B(G543), .Z(new_n540));
  NAND2_X1  g115(.A1(new_n523), .A2(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G168));
  XOR2_X1   g119(.A(KEYINPUT77), .B(G52), .Z(new_n545));
  NAND2_X1  g120(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n547), .B2(new_n524), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n514), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(G171));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n524), .A2(new_n552), .B1(new_n553), .B2(new_n527), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n514), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n540), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n521), .A2(new_n522), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n540), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n566), .A2(G651), .B1(new_n568), .B2(G91), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT78), .B(KEYINPUT9), .Z(new_n570));
  NAND3_X1  g145(.A1(new_n537), .A2(G53), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n527), .A2(new_n572), .B1(new_n573), .B2(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n571), .B2(new_n574), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n569), .B1(new_n576), .B2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n568), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n537), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n540), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n537), .B2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n568), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n568), .A2(G85), .B1(new_n537), .B2(G47), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT80), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n514), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n568), .A2(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n527), .B2(KEYINPUT81), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n540), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n602), .A2(new_n604), .B1(new_n607), .B2(G651), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G284));
  XOR2_X1   g185(.A(G284), .B(KEYINPUT82), .Z(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  INV_X1    g192(.A(new_n557), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n601), .A2(new_n608), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n622), .B2(new_n619), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT83), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g200(.A(new_n491), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G123), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT85), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n627), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n489), .A2(new_n465), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT13), .B(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n635), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT87), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT17), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT88), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT90), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n662), .A2(new_n665), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT89), .ZN(new_n669));
  INV_X1    g244(.A(new_n661), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n663), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n667), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n680), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(KEYINPUT34), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(G23), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G288), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  OAI21_X1  g280(.A(G1976), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n701), .A2(new_n702), .ZN(new_n707));
  INV_X1    g282(.A(G1976), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(new_n708), .A3(new_n703), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G22), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G166), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n699), .A2(G6), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G305), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n722), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n724), .A2(new_n720), .A3(new_n715), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n710), .A2(new_n714), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(KEYINPUT95), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(KEYINPUT95), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n698), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n710), .A2(new_n714), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n723), .A2(new_n725), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n726), .A2(KEYINPUT95), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n699), .A2(G24), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT93), .Z(new_n737));
  INV_X1    g312(.A(G290), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n699), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1986), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G25), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G107), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT91), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n483), .A2(G119), .ZN(new_n747));
  INV_X1    g322(.A(G131), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n746), .B(new_n747), .C1(new_n491), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n742), .B1(new_n754), .B2(new_n741), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT35), .B(G1991), .Z(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n740), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n729), .A2(new_n735), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(KEYINPUT36), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n729), .A2(new_n762), .A3(new_n735), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n699), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n613), .B2(new_n699), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT101), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(KEYINPUT101), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT100), .B(G1956), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n741), .A2(G35), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n493), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n741), .A2(G33), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  AOI22_X1  g355(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G139), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n780), .B1(new_n470), .B2(new_n781), .C1(new_n491), .C2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(new_n741), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n785), .A2(G2072), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n699), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n699), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT99), .B(G1966), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(G164), .A2(G29), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G27), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2078), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n777), .A2(new_n786), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n741), .A2(G32), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n626), .A2(G141), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n466), .A2(G105), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT26), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n798), .B(new_n800), .C1(G129), .C2(new_n483), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT27), .B(G1996), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT97), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n776), .A2(G2090), .ZN(new_n808));
  AND4_X1   g383(.A1(new_n772), .A2(new_n795), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n741), .A2(G26), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT28), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n483), .A2(G128), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n470), .A2(G116), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(G140), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n812), .B1(new_n813), .B2(new_n814), .C1(new_n491), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G29), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT96), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(KEYINPUT96), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n811), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n699), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n557), .B2(new_n699), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1341), .Z(new_n825));
  NOR2_X1   g400(.A1(G171), .A2(new_n699), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G5), .B2(new_n699), .ZN(new_n827));
  INV_X1    g402(.A(G1961), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n632), .A2(G29), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n825), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G4), .A2(G16), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n609), .B2(G16), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n831), .B1(G1348), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(G1348), .ZN(new_n835));
  AND2_X1   g410(.A1(KEYINPUT24), .A2(G34), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n741), .B1(KEYINPUT24), .B2(G34), .ZN(new_n837));
  OAI22_X1  g412(.A1(G160), .A2(new_n741), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(G2084), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(G2084), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n835), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT30), .B(G28), .ZN(new_n842));
  OR2_X1    g417(.A1(KEYINPUT31), .A2(G11), .ZN(new_n843));
  NAND2_X1  g418(.A1(KEYINPUT31), .A2(G11), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n842), .A2(new_n741), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI221_X1 g420(.A(new_n845), .B1(new_n803), .B2(new_n805), .C1(new_n827), .C2(new_n828), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n785), .A2(G2072), .B1(new_n793), .B2(new_n792), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g423(.A1(new_n822), .A2(new_n834), .A3(new_n841), .A4(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n770), .A2(new_n771), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n809), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT102), .B1(new_n764), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  AOI211_X1 g429(.A(new_n854), .B(new_n851), .C1(new_n761), .C2(new_n763), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(G311));
  NAND2_X1  g431(.A1(new_n764), .A2(new_n852), .ZN(G150));
  NAND2_X1  g432(.A1(new_n609), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  INV_X1    g435(.A(G55), .ZN(new_n861));
  OAI22_X1  g436(.A1(new_n524), .A2(new_n860), .B1(new_n861), .B2(new_n527), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n514), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n557), .A2(new_n865), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n556), .A2(new_n554), .B1(new_n862), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n859), .B(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n865), .A2(new_n872), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT103), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(G145));
  XNOR2_X1  g453(.A(G160), .B(new_n493), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n632), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n816), .B(new_n512), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(new_n784), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n784), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n882), .A2(new_n883), .A3(new_n802), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n802), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n638), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n626), .A2(G142), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n470), .A2(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n483), .A2(G130), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n753), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n753), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n888), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n638), .A3(new_n896), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n901), .A3(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n887), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n902), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(new_n886), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n880), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n880), .B1(new_n887), .B2(new_n903), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n886), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT40), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G395));
  XNOR2_X1  g490(.A(G166), .B(G288), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n594), .A2(G305), .A3(new_n596), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G305), .B1(new_n594), .B2(new_n596), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  INV_X1    g496(.A(G288), .ZN(new_n922));
  XNOR2_X1  g497(.A(G166), .B(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n923), .A3(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n869), .B1(G559), .B2(new_n621), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n622), .A2(new_n868), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n575), .B(KEYINPUT79), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(new_n569), .A3(new_n601), .A4(new_n608), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n621), .A2(G299), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR3_X1    g508(.A1(new_n929), .A2(KEYINPUT105), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT41), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n929), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT105), .B1(new_n929), .B2(new_n933), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n934), .A2(new_n942), .A3(new_n938), .A4(new_n939), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n926), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(new_n619), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n926), .A3(new_n943), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT107), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n865), .B2(G868), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n945), .B2(new_n946), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(G295));
  NOR2_X1   g526(.A1(new_n948), .A2(new_n950), .ZN(G331));
  OAI22_X1  g527(.A1(new_n543), .A2(new_n539), .B1(new_n548), .B2(new_n550), .ZN(new_n953));
  INV_X1    g528(.A(new_n543), .ZN(new_n954));
  INV_X1    g529(.A(new_n550), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n568), .A2(G90), .B1(new_n537), .B2(new_n545), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n532), .A2(new_n535), .B1(new_n537), .B2(G51), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n868), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n866), .A2(new_n953), .A3(new_n958), .A4(new_n867), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(KEYINPUT108), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n869), .A2(new_n963), .A3(new_n953), .A4(new_n958), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n933), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n960), .A2(new_n961), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n936), .A2(new_n937), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n969), .A3(new_n925), .ZN(new_n970));
  INV_X1    g545(.A(G37), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n925), .B1(new_n967), .B2(new_n969), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n936), .A2(new_n937), .ZN(new_n975));
  OAI22_X1  g550(.A1(new_n975), .A2(new_n965), .B1(new_n933), .B2(new_n968), .ZN(new_n976));
  INV_X1    g551(.A(new_n925), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n971), .A4(new_n970), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n980), .A3(KEYINPUT109), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(KEYINPUT43), .C1(new_n972), .C2(new_n973), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n972), .A2(KEYINPUT43), .A3(new_n973), .ZN(new_n989));
  INV_X1    g564(.A(new_n978), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT43), .B1(new_n990), .B2(new_n972), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT44), .ZN(new_n992));
  OAI22_X1  g567(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n992), .ZN(G397));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n498), .B1(new_n468), .B2(new_n495), .ZN(new_n996));
  AND4_X1   g571(.A1(new_n498), .A2(new_n474), .A3(new_n476), .A4(new_n495), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n511), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n503), .A2(new_n510), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n472), .A2(G40), .A3(new_n467), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n471), .A3(new_n481), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT56), .B(G2072), .Z(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n512), .A2(new_n1012), .A3(new_n995), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1006), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1956), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT113), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1010), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n569), .A2(new_n575), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n613), .A2(KEYINPUT57), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n994), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1010), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1019), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1018), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT116), .A3(new_n1023), .ZN(new_n1030));
  INV_X1    g605(.A(G1348), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1014), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1005), .A2(new_n1000), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n821), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n609), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1025), .A2(new_n1030), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT115), .B1(new_n1029), .B2(new_n1023), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1020), .A2(new_n1039), .A3(new_n1024), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1008), .A2(G1996), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT58), .B(G1341), .Z(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1005), .B2(new_n1000), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n618), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT59), .Z(new_n1047));
  INV_X1    g622(.A(KEYINPUT61), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1025), .A2(new_n1049), .A3(new_n1030), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n1035), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1032), .A2(new_n1053), .A3(KEYINPUT60), .A4(new_n1034), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n609), .A3(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT117), .B(new_n621), .C1(new_n1035), .C2(new_n1051), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1035), .A2(new_n1051), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1047), .A2(new_n1050), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1029), .A2(new_n1023), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT61), .B1(new_n1041), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1042), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1033), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  INV_X1    g640(.A(G1981), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n590), .A2(new_n1066), .A3(new_n591), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT112), .B(G86), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n568), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1066), .B1(new_n590), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1065), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n590), .A2(new_n1070), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT49), .B(new_n1067), .C1(new_n1073), .C2(new_n1066), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1064), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n922), .A2(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n708), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1064), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1076), .B(G8), .C1(new_n1005), .C2(new_n1000), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT52), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1075), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1014), .A2(G2090), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1008), .A2(new_n713), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1063), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G303), .A2(G8), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(G303), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1081), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1008), .B2(G2078), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1014), .A2(new_n828), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OR3_X1    g674(.A1(new_n1008), .A2(new_n1096), .A3(G2078), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n793), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n479), .A2(KEYINPUT121), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n470), .B1(new_n479), .B2(KEYINPUT121), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(new_n1098), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G171), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1095), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1099), .A2(G301), .A3(new_n1100), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(G171), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(KEYINPUT54), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1094), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1966), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1008), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G2084), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1011), .A2(new_n1006), .A3(new_n1116), .A4(new_n1013), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(G168), .A2(new_n1063), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1011), .A2(new_n1006), .A3(new_n1013), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1121), .A2(new_n1116), .B1(new_n1008), .B2(new_n1114), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1063), .B1(new_n1122), .B2(G168), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT51), .B1(new_n1123), .B2(KEYINPUT118), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT118), .B(G8), .C1(new_n1118), .C2(G286), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT119), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1063), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT118), .B(KEYINPUT51), .C1(new_n1131), .C2(new_n1119), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n1120), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1113), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1062), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1129), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1134), .B1(new_n1133), .B2(new_n1120), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1120), .ZN(new_n1141));
  AOI211_X1 g716(.A(KEYINPUT119), .B(new_n1141), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT62), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1093), .A2(new_n1081), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1075), .A2(new_n708), .A3(new_n922), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1064), .B1(new_n1147), .B2(new_n1068), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1122), .A2(new_n1063), .A3(G286), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1094), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1094), .A2(KEYINPUT63), .A3(new_n1150), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1137), .A2(new_n1145), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n754), .A2(new_n756), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n754), .A2(new_n756), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n816), .B(new_n821), .ZN(new_n1160));
  INV_X1    g735(.A(G1996), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n802), .B(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(G290), .B(G1986), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1157), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1156), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1167));
  AND2_X1   g742(.A1(KEYINPUT123), .A2(KEYINPUT46), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1160), .A2(new_n797), .A3(new_n801), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1157), .ZN(new_n1171));
  OAI221_X1 g746(.A(new_n1169), .B1(KEYINPUT123), .B2(KEYINPUT46), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT47), .Z(new_n1173));
  NAND3_X1  g748(.A1(new_n1163), .A2(KEYINPUT124), .A3(new_n1157), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1171), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT126), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1175), .B(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT124), .B1(new_n1163), .B2(new_n1157), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n816), .A2(G2067), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1162), .A2(new_n1160), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(new_n1159), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n754), .A2(KEYINPUT122), .A3(new_n756), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1181), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1179), .A2(new_n1180), .B1(new_n1171), .B2(new_n1186), .ZN(new_n1187));
  OR3_X1    g762(.A1(new_n1173), .A2(new_n1187), .A3(KEYINPUT127), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT127), .B1(new_n1173), .B2(new_n1187), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1166), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g766(.A1(G227), .A2(new_n463), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n696), .A2(new_n658), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n1194), .B1(new_n909), .B2(new_n912), .ZN(new_n1195));
  AND2_X1   g769(.A1(new_n981), .A2(new_n984), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1196), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


