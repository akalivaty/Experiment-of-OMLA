//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n522, new_n523, new_n524, new_n525, new_n526, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n538, new_n539, new_n540, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n461), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n461), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  MUX2_X1   g050(.A(G100), .B(G112), .S(G2105), .Z(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G124), .B1(G2104), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(new_n463), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT68), .Z(G162));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  OAI211_X1 g057(.A(G138), .B(new_n462), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n461), .A2(new_n485), .A3(G138), .A4(new_n462), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n481), .C2(new_n482), .ZN(new_n489));
  OR2_X1    g064(.A1(KEYINPUT69), .A2(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT69), .A2(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n462), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n488), .A2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  INV_X1    g078(.A(G88), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n501), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n509), .A2(new_n499), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT72), .B(G89), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n513), .B(new_n514), .C1(new_n507), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n505), .A2(G543), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT71), .B(G51), .Z(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n516), .A2(new_n519), .ZN(G286));
  INV_X1    g095(.A(G286), .ZN(G168));
  NAND2_X1  g096(.A1(new_n502), .A2(G52), .ZN(new_n522));
  INV_X1    g097(.A(G90), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(new_n507), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n499), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(G171));
  AOI22_X1  g102(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n499), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n502), .A2(G43), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(new_n507), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(G153));
  AND3_X1   g110(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G36), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT73), .Z(G188));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n506), .B(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(G78), .A2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(G651), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G53), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT9), .B1(new_n517), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n502), .A2(new_n550), .A3(G53), .ZN(new_n551));
  INV_X1    g126(.A(new_n507), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n549), .A2(new_n551), .B1(G91), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n547), .A2(new_n553), .ZN(G299));
  INV_X1    g129(.A(G171), .ZN(G301));
  INV_X1    g130(.A(G166), .ZN(G303));
  NAND2_X1  g131(.A1(new_n552), .A2(G87), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n502), .A2(G49), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(G288));
  NAND2_X1  g135(.A1(new_n506), .A2(G61), .ZN(new_n561));
  INV_X1    g136(.A(G73), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n562), .B2(new_n496), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n562), .A2(new_n496), .A3(KEYINPUT75), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  INV_X1    g142(.A(G86), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n507), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n505), .A2(KEYINPUT76), .A3(G86), .A4(new_n506), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n502), .A2(G48), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n499), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n552), .A2(G85), .B1(G47), .B2(new_n502), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G290));
  AND3_X1   g152(.A1(new_n505), .A2(G92), .A3(new_n506), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(KEYINPUT10), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(new_n580), .B1(G54), .B2(new_n502), .ZN(new_n581));
  INV_X1    g156(.A(G66), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n543), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT78), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G171), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT79), .Z(G284));
  INV_X1    g167(.A(new_n591), .ZN(G321));
  MUX2_X1   g168(.A(G286), .B(G299), .S(new_n588), .Z(G297));
  MUX2_X1   g169(.A(G286), .B(G299), .S(new_n588), .Z(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n587), .B1(new_n596), .B2(G860), .ZN(G148));
  INV_X1    g172(.A(new_n534), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(new_n587), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(G559), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n599), .B1(new_n601), .B2(G868), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g178(.A1(new_n464), .A2(G2104), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT13), .Z(new_n606));
  INV_X1    g181(.A(G2100), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n464), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n475), .A2(G123), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(KEYINPUT80), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(KEYINPUT80), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(G111), .C2(new_n462), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n610), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND3_X1  g192(.A1(new_n608), .A2(new_n609), .A3(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(G2443), .B(G2446), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT82), .ZN(new_n620));
  XOR2_X1   g195(.A(G2451), .B(G2454), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2427), .ZN(new_n630));
  INV_X1    g205(.A(G2430), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n626), .A2(new_n633), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n634), .A2(G14), .A3(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT18), .ZN(new_n643));
  INV_X1    g218(.A(new_n639), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .A3(new_n637), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n637), .B1(new_n644), .B2(KEYINPUT17), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(new_n641), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n638), .A2(new_n641), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n648), .B2(KEYINPUT17), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n643), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT83), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(G227));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n656), .C2(new_n662), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G29), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G25), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  MUX2_X1   g248(.A(G95), .B(G107), .S(G2105), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G2104), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT86), .Z(new_n676));
  INV_X1    g251(.A(G119), .ZN(new_n677));
  INV_X1    g252(.A(G131), .ZN(new_n678));
  OAI22_X1  g253(.A1(new_n677), .A2(new_n474), .B1(new_n463), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n673), .B1(new_n680), .B2(new_n671), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT87), .Z(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT35), .B(G1991), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G24), .B(G290), .S(G16), .Z(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G1986), .Z(new_n686));
  MUX2_X1   g261(.A(G6), .B(G305), .S(G16), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G166), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G1971), .Z(new_n698));
  NAND3_X1  g273(.A1(new_n689), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n684), .B(new_n686), .C1(KEYINPUT34), .C2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(KEYINPUT34), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT36), .Z(new_n702));
  NOR2_X1   g277(.A1(G171), .A2(new_n690), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G5), .B2(new_n690), .ZN(new_n704));
  INV_X1    g279(.A(G1961), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G2078), .ZN(new_n707));
  NAND2_X1  g282(.A1(G164), .A2(G29), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G27), .B2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n706), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n475), .A2(G129), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT88), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n465), .A2(G105), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT26), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n713), .B(new_n715), .C1(new_n464), .C2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(new_n671), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n671), .B2(G32), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n690), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n690), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G1966), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(new_n721), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n671), .A2(G26), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n464), .A2(G140), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n475), .A2(G128), .ZN(new_n730));
  MUX2_X1   g305(.A(G104), .B(G116), .S(G2105), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G2104), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(new_n671), .ZN(new_n735));
  INV_X1    g310(.A(G2067), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n722), .A2(new_n725), .A3(new_n726), .A4(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n710), .B(new_n738), .C1(new_n707), .C2(new_n709), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n724), .A2(G1966), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT89), .Z(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n587), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G4), .B2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n741), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n742), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n616), .A2(new_n671), .ZN(new_n747));
  OR2_X1    g322(.A1(KEYINPUT30), .A2(G28), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT30), .A2(G28), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  NOR3_X1   g326(.A1(new_n747), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n671), .A2(G33), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n465), .A2(G103), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT25), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(KEYINPUT25), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(new_n756), .B1(G139), .B2(new_n464), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n462), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2072), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n752), .B1(new_n760), .B2(new_n761), .C1(new_n704), .C2(new_n705), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g338(.A1(KEYINPUT24), .A2(G34), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  AOI21_X1  g341(.A(G29), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G160), .B2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(G2084), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n534), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1341), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n768), .A2(G2084), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n762), .A2(new_n769), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n739), .A2(new_n746), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n671), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n671), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT29), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(G2090), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(G2090), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT90), .B(KEYINPUT23), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n690), .A2(G20), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1956), .Z(new_n785));
  NOR4_X1   g360(.A1(new_n775), .A2(new_n779), .A3(new_n780), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n702), .A2(new_n786), .ZN(G150));
  INV_X1    g362(.A(G150), .ZN(G311));
  NAND2_X1  g363(.A1(new_n502), .A2(G55), .ZN(new_n789));
  INV_X1    g364(.A(G93), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n507), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(new_n499), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G860), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT93), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT37), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n795), .B(new_n598), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n600), .A2(new_n596), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(KEYINPUT39), .ZN(new_n805));
  INV_X1    g380(.A(G860), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n804), .B2(KEYINPUT39), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n798), .B1(new_n805), .B2(new_n807), .ZN(G145));
  XNOR2_X1  g383(.A(new_n680), .B(KEYINPUT96), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(new_n605), .ZN(new_n810));
  MUX2_X1   g385(.A(G106), .B(G118), .S(G2105), .Z(new_n811));
  AOI22_X1  g386(.A1(new_n475), .A2(G130), .B1(G2104), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G142), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n463), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT97), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n810), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n717), .B(new_n759), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n494), .A2(KEYINPUT95), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT95), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n489), .B(new_n821), .C1(new_n492), .C2(new_n493), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n487), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n734), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n819), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n818), .A2(new_n825), .ZN(new_n827));
  XNOR2_X1  g402(.A(G162), .B(new_n616), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n472), .B(KEYINPUT94), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G37), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n831), .B1(new_n816), .B2(new_n825), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n825), .B2(new_n816), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(G395));
  NOR2_X1   g413(.A1(new_n795), .A2(G868), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n799), .B(new_n601), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n587), .A2(G299), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n587), .A2(G299), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(KEYINPUT41), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(new_n846), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n842), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n845), .B1(new_n849), .B2(KEYINPUT41), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n844), .B1(new_n850), .B2(new_n840), .ZN(new_n851));
  XNOR2_X1  g426(.A(G290), .B(G288), .ZN(new_n852));
  XNOR2_X1  g427(.A(G305), .B(G166), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT42), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n851), .B(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n839), .B1(new_n856), .B2(G868), .ZN(G295));
  AOI21_X1  g432(.A(new_n839), .B1(new_n856), .B2(G868), .ZN(G331));
  XNOR2_X1  g433(.A(G301), .B(G286), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n799), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n843), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n860), .B(new_n845), .C1(new_n849), .C2(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n854), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(G37), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n860), .A2(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n849), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(new_n854), .C1(new_n843), .C2(new_n867), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT101), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT101), .B1(new_n862), .B2(new_n863), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n854), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n866), .A2(new_n875), .A3(KEYINPUT43), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT44), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n870), .A2(KEYINPUT43), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n866), .A2(new_n875), .A3(new_n871), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(KEYINPUT44), .B2(new_n880), .ZN(G397));
  INV_X1    g456(.A(G1384), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n487), .A2(new_n822), .ZN(new_n883));
  INV_X1    g458(.A(new_n491), .ZN(new_n884));
  NOR2_X1   g459(.A1(KEYINPUT69), .A2(G114), .ZN(new_n885));
  OAI21_X1  g460(.A(G2105), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n493), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n821), .B1(new_n888), .B2(new_n489), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n882), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n466), .A2(new_n471), .A3(G40), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(G290), .A2(G1986), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT103), .Z(new_n898));
  NAND2_X1  g473(.A1(G290), .A2(G1986), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G1996), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT104), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n718), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n733), .B(new_n736), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(G1996), .B2(new_n717), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n896), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n680), .B(new_n683), .Z(new_n909));
  AOI211_X1 g484(.A(new_n900), .B(new_n908), .C1(new_n895), .C2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n882), .B1(new_n488), .B2(new_n494), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT50), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n893), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n890), .A2(KEYINPUT106), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n916), .B(new_n882), .C1(new_n883), .C2(new_n889), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n913), .A4(new_n917), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n891), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n894), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  INV_X1    g500(.A(new_n917), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n916), .B1(new_n823), .B2(new_n882), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n707), .A2(KEYINPUT53), .ZN(new_n930));
  OAI22_X1  g505(.A1(new_n922), .A2(G1961), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT124), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT124), .ZN(new_n933));
  OAI221_X1 g508(.A(new_n933), .B1(new_n929), .B2(new_n930), .C1(new_n922), .C2(G1961), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n911), .A2(new_n891), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n823), .A2(KEYINPUT45), .A3(new_n882), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n893), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT105), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n707), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT53), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n932), .A2(new_n934), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G171), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n466), .A2(KEYINPUT53), .A3(G40), .A4(new_n707), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n470), .B(KEYINPUT125), .Z(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(G2105), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n892), .A3(new_n936), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n941), .B(new_n947), .C1(G1961), .C2(new_n922), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n943), .B1(G171), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT113), .B(G2084), .Z(new_n952));
  AOI211_X1 g527(.A(new_n914), .B(new_n952), .C1(new_n920), .C2(new_n921), .ZN(new_n953));
  AOI21_X1  g528(.A(G1966), .B1(new_n924), .B2(new_n928), .ZN(new_n954));
  OAI21_X1  g529(.A(G8), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G286), .A2(G8), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n955), .A2(KEYINPUT122), .A3(KEYINPUT51), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G168), .B2(new_n955), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n960), .A2(KEYINPUT51), .B1(new_n955), .B2(new_n956), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G303), .A2(G8), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT55), .Z(new_n965));
  INV_X1    g540(.A(G2090), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n922), .A2(KEYINPUT108), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G1971), .B2(new_n938), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT108), .B1(new_n922), .B2(new_n966), .ZN(new_n969));
  OAI211_X1 g544(.A(G8), .B(new_n965), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n926), .A2(new_n927), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(new_n893), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n692), .A2(G1976), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(G1976), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(G288), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n915), .A2(new_n893), .A3(new_n917), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(G8), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT52), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n565), .A2(G651), .B1(G48), .B2(new_n502), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n570), .A4(new_n569), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n552), .A2(G86), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n984), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n982), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n983), .A2(new_n987), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT49), .B(new_n985), .C1(new_n990), .C2(new_n984), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n989), .A2(new_n978), .A3(new_n991), .A4(G8), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT110), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n981), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n915), .A2(KEYINPUT50), .A3(new_n917), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n911), .A2(new_n913), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n894), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n966), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n938), .B2(G1971), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n965), .B1(new_n999), .B2(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n994), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n970), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n942), .A2(G171), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n948), .B2(G171), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n951), .A2(new_n963), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT121), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n978), .A2(G2067), .ZN(new_n1009));
  INV_X1    g584(.A(new_n914), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT107), .B1(new_n972), .B2(new_n913), .ZN(new_n1011));
  INV_X1    g586(.A(new_n921), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1009), .B1(new_n1013), .B2(new_n742), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1014), .A2(KEYINPUT120), .A3(KEYINPUT60), .A4(new_n600), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1009), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT60), .B(new_n1017), .C1(new_n922), .C2(G1348), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1018), .B2(new_n587), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n587), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1014), .A2(KEYINPUT60), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT56), .B(G2072), .Z(new_n1024));
  OR2_X1    g599(.A1(new_n937), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n997), .B2(G1956), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT115), .B(new_n1025), .C1(new_n997), .C2(G1956), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G299), .A2(KEYINPUT114), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(G299), .A2(KEYINPUT114), .A3(KEYINPUT57), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1030), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1035), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(new_n1025), .C1(G1956), .C2(new_n997), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1038), .A2(KEYINPUT61), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT117), .B(G1996), .Z(new_n1041));
  NOR2_X1   g616(.A1(new_n937), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT58), .B(G1341), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n978), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n978), .A2(KEYINPUT118), .A3(new_n1043), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT119), .B1(new_n1048), .B2(new_n598), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n978), .A2(KEYINPUT118), .A3(new_n1043), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT118), .B1(new_n978), .B2(new_n1043), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1050), .A2(new_n1051), .B1(new_n937), .B2(new_n1041), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n534), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(KEYINPUT59), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1048), .A2(KEYINPUT119), .A3(new_n598), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1053), .B1(new_n1052), .B2(new_n534), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT61), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1038), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1026), .A2(new_n1035), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1040), .A2(new_n1055), .A3(new_n1059), .A4(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1023), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1014), .A2(new_n600), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1037), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1038), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT116), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1070), .B(new_n1038), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1008), .B1(new_n1065), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1063), .A2(new_n1055), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1059), .A4(new_n1040), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1076), .A2(KEYINPUT121), .A3(new_n1071), .A4(new_n1069), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1007), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT62), .B1(new_n958), .B2(new_n961), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT126), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT126), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(KEYINPUT62), .C1(new_n958), .C2(new_n961), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n962), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1002), .A2(new_n943), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G288), .A2(G1976), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n993), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n973), .B1(new_n1088), .B2(new_n986), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n981), .A2(new_n993), .A3(KEYINPUT111), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT111), .B1(new_n981), .B2(new_n993), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1092), .B2(new_n970), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1089), .B(KEYINPUT112), .C1(new_n1092), .C2(new_n970), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  OAI211_X1 g672(.A(G8), .B(G168), .C1(new_n953), .C2(new_n954), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1002), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(G8), .B1(new_n968), .B2(new_n969), .ZN(new_n1100));
  INV_X1    g675(.A(new_n965), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n994), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n981), .A2(new_n993), .A3(KEYINPUT111), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1098), .A2(new_n1097), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1102), .A2(new_n1106), .A3(new_n970), .A4(new_n1107), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1095), .A2(new_n1096), .B1(new_n1099), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1086), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n910), .B1(new_n1078), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n896), .B1(new_n718), .B2(new_n905), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n903), .B2(KEYINPUT46), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(KEYINPUT46), .B2(new_n903), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  OR4_X1    g691(.A1(new_n676), .A2(new_n908), .A3(new_n679), .A4(new_n683), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n734), .A2(new_n736), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n896), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n908), .B1(new_n895), .B2(new_n909), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n898), .A2(new_n896), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT48), .Z(new_n1122));
  AOI211_X1 g697(.A(new_n1116), .B(new_n1119), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1111), .A2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g699(.A1(new_n872), .A2(new_n876), .ZN(new_n1126));
  OR3_X1    g700(.A1(G229), .A2(G401), .A3(new_n459), .ZN(new_n1127));
  NOR3_X1   g701(.A1(new_n836), .A2(G227), .A3(new_n1127), .ZN(new_n1128));
  AND2_X1   g702(.A1(new_n1126), .A2(new_n1128), .ZN(G308));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(G225));
endmodule


