//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n442, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(new_n442), .A2(G57), .A3(G69), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT67), .A4(G125), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT68), .Z(G160));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n466), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n473), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n473), .A3(new_n483), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  NOR2_X1   g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n486), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n463), .A2(new_n465), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n497));
  NOR2_X1   g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(new_n473), .B2(G114), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n463), .A2(new_n465), .A3(new_n473), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n501), .A2(KEYINPUT72), .A3(new_n502), .A4(G138), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n473), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT4), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n505), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT71), .B1(new_n505), .B2(KEYINPUT4), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n500), .B1(new_n507), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(G50), .A2(new_n519), .B1(new_n524), .B2(G88), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OR3_X1    g101(.A1(new_n523), .A2(KEYINPUT74), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT74), .B1(new_n523), .B2(new_n526), .ZN(new_n528));
  INV_X1    g103(.A(G75), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT75), .B1(new_n529), .B2(new_n518), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n529), .A2(new_n518), .A3(KEYINPUT75), .ZN(new_n532));
  OAI21_X1  g107(.A(G651), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n519), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(new_n517), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT76), .B(G89), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(new_n540), .B1(G63), .B2(G651), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n536), .B(new_n538), .C1(new_n541), .C2(new_n523), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(new_n523), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT77), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(G52), .A2(new_n519), .B1(new_n524), .B2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n524), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n519), .A2(G43), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n544), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n515), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n514), .A2(G53), .A3(G543), .A4(new_n516), .ZN(new_n563));
  XOR2_X1   g138(.A(KEYINPUT78), .B(KEYINPUT9), .Z(new_n564));
  OR2_X1    g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n524), .A2(G91), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT79), .B(G65), .Z(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n570), .B2(new_n523), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n565), .A2(new_n566), .A3(new_n568), .A4(new_n572), .ZN(G299));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n514), .A2(G49), .A3(G543), .A4(new_n516), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n514), .A2(G87), .A3(new_n544), .A4(new_n516), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n515), .B1(new_n523), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  AND4_X1   g159(.A1(new_n574), .A2(new_n578), .A3(new_n581), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n583), .B1(new_n576), .B2(new_n577), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n574), .B1(new_n586), .B2(new_n581), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n585), .A2(new_n587), .ZN(G288));
  NAND4_X1  g163(.A1(new_n514), .A2(G86), .A3(new_n544), .A4(new_n516), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n514), .A2(G48), .A3(G543), .A4(new_n516), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n523), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n524), .A2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n519), .A2(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n544), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(new_n515), .C2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n601));
  NAND3_X1  g176(.A1(new_n524), .A2(G92), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n519), .A2(G54), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n544), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n515), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n524), .A2(G92), .ZN(new_n607));
  INV_X1    g182(.A(new_n601), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n604), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G284));
  XOR2_X1   g187(.A(G284), .B(KEYINPUT84), .Z(G321));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G299), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n555), .A2(new_n614), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n610), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n485), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n488), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n466), .A2(new_n476), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT85), .B(G2100), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT87), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2443), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n657), .B(KEYINPUT88), .Z(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  OAI221_X1 g240(.A(new_n659), .B1(new_n660), .B2(new_n661), .C1(new_n663), .C2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n629), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2100), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT89), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT19), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT90), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(KEYINPUT20), .A3(new_n675), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n672), .A2(new_n677), .ZN(new_n681));
  OAI221_X1 g256(.A(new_n678), .B1(new_n680), .B2(new_n672), .C1(new_n681), .C2(KEYINPUT20), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1991), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1996), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n687), .B(new_n689), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G11), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT29), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(G2090), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT99), .ZN(new_n698));
  NAND2_X1  g273(.A1(G299), .A2(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT23), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G20), .ZN(new_n702));
  MUX2_X1   g277(.A(KEYINPUT23), .B(new_n700), .S(new_n702), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G1956), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n697), .A2(KEYINPUT99), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n703), .A2(G1956), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n698), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n701), .A2(G21), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G168), .B2(new_n701), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT97), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1966), .ZN(new_n711));
  INV_X1    g286(.A(G2084), .ZN(new_n712));
  NAND2_X1  g287(.A1(G160), .A2(G29), .ZN(new_n713));
  NOR2_X1   g288(.A1(KEYINPUT24), .A2(G34), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  AOI21_X1  g291(.A(G29), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT96), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n713), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n711), .B1(new_n712), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n701), .A2(G4), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n611), .B2(new_n701), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1348), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n693), .A2(G27), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G164), .B2(new_n693), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2078), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n701), .A2(G19), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n556), .B2(new_n701), .ZN(new_n731));
  OR2_X1    g306(.A1(G29), .A2(G32), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n485), .A2(G129), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n488), .A2(G141), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n733), .A2(new_n734), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(new_n693), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n731), .A2(G1341), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(G171), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G5), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n731), .A2(G1341), .B1(new_n739), .B2(new_n740), .ZN(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(KEYINPUT30), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n628), .B2(new_n693), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n693), .A2(G33), .ZN(new_n751));
  NAND2_X1  g326(.A1(G115), .A2(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G127), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n466), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2105), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT25), .Z(new_n757));
  INV_X1    g332(.A(G139), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n757), .C1(new_n487), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2072), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n750), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n729), .A2(new_n745), .A3(new_n746), .A4(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n742), .B(G1961), .C1(G5), .C2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n693), .A2(G26), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n485), .A2(G128), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n488), .A2(G140), .ZN(new_n770));
  NOR2_X1   g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(new_n473), .B2(G116), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n769), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G29), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n768), .B(new_n774), .S(KEYINPUT28), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n696), .A2(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n721), .A2(new_n712), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n767), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n707), .A2(new_n722), .A3(new_n765), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G25), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT93), .B1(new_n781), .B2(G29), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n781), .A2(KEYINPUT93), .A3(G29), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n485), .A2(G119), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n488), .A2(G131), .ZN(new_n785));
  NOR2_X1   g360(.A1(G95), .A2(G2105), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n782), .B(new_n783), .C1(new_n792), .C2(new_n693), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT35), .B(G1991), .Z(new_n794));
  XOR2_X1   g369(.A(new_n793), .B(new_n794), .Z(new_n795));
  AND3_X1   g370(.A1(new_n578), .A2(new_n581), .A3(new_n584), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(new_n701), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n701), .B2(G23), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT33), .B(G1976), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT95), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n701), .A2(G6), .ZN(new_n802));
  INV_X1    g377(.A(G305), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n701), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n798), .A2(new_n800), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n701), .A2(G22), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G303), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1971), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n801), .A2(new_n806), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n795), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n816));
  MUX2_X1   g391(.A(G24), .B(G290), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1986), .Z(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n816), .B1(new_n815), .B2(new_n818), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n692), .B(new_n780), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n813), .A2(new_n814), .ZN(new_n825));
  INV_X1    g400(.A(new_n795), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(new_n818), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n819), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n829), .A2(KEYINPUT100), .A3(new_n692), .A4(new_n780), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n824), .A2(new_n830), .ZN(G311));
  NAND2_X1  g406(.A1(new_n822), .A2(KEYINPUT101), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n829), .A2(new_n833), .A3(new_n692), .A4(new_n780), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(G150));
  NAND2_X1  g410(.A1(new_n524), .A2(G93), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n519), .A2(G55), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n544), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(new_n515), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NOR2_X1   g417(.A1(new_n610), .A2(new_n618), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n840), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n555), .B1(new_n846), .B2(KEYINPUT102), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n845), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n851), .B2(G860), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT71), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n505), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n856), .A2(new_n503), .A3(new_n506), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n499), .A2(new_n498), .ZN(new_n859));
  INV_X1    g434(.A(new_n497), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n759), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n738), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n773), .B(KEYINPUT103), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G142), .ZN(new_n868));
  NOR2_X1   g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n487), .A2(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(G130), .B2(new_n485), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n632), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n791), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n867), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G160), .B(new_n628), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G162), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n867), .A2(new_n874), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT104), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n875), .A2(new_n879), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(KEYINPUT105), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n879), .B1(new_n875), .B2(new_n876), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n889), .B2(new_n882), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n890), .B2(new_n885), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n853), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(KEYINPUT105), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n888), .A3(new_n885), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(G395));
  XNOR2_X1  g471(.A(new_n850), .B(KEYINPUT106), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n621), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n610), .B(G299), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n899), .B(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT107), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT107), .B1(new_n899), .B2(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(new_n803), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n796), .B(G290), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n586), .A2(new_n581), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G290), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT108), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(KEYINPUT108), .A3(new_n907), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  AND4_X1   g496(.A1(new_n901), .A2(new_n906), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n901), .A2(new_n906), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G868), .B2(new_n846), .ZN(G295));
  OAI21_X1  g500(.A(new_n924), .B1(G868), .B2(new_n846), .ZN(G331));
  XNOR2_X1  g501(.A(G301), .B(G168), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n850), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n903), .B2(new_n905), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n900), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n932), .B2(new_n918), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n899), .B(new_n934), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n930), .B(KEYINPUT110), .C1(new_n935), .C2(new_n928), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n916), .B(KEYINPUT109), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n928), .A2(new_n935), .A3(KEYINPUT110), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n933), .A2(KEYINPUT43), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n931), .B2(new_n929), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT43), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n933), .A2(new_n945), .A3(new_n939), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n933), .B2(new_n941), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(G397));
  NOR2_X1   g524(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n858), .B2(new_n862), .ZN(new_n951));
  INV_X1    g526(.A(G40), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n952), .B(new_n477), .C1(new_n471), .C2(G2105), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT58), .B(G1341), .Z(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G164), .B2(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n951), .A2(KEYINPUT45), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n953), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n960), .B2(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n556), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT59), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT59), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n964), .A3(new_n556), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n950), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n953), .B1(new_n951), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n863), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT117), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n951), .A2(KEYINPUT117), .A3(new_n967), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(G2072), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n974), .A2(G1956), .B1(new_n960), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(G299), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n979));
  NOR2_X1   g554(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n980));
  NAND2_X1  g555(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(G299), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n978), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n863), .B2(new_n969), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n957), .B(G1384), .C1(new_n858), .C2(new_n862), .ZN(new_n988));
  INV_X1    g563(.A(new_n953), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n976), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n984), .B(new_n991), .C1(G1956), .C2(new_n974), .ZN(new_n992));
  NAND2_X1  g567(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n986), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n986), .B2(new_n992), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n966), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT122), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n954), .A2(G2067), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n999), .A2(KEYINPUT120), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT120), .ZN(new_n1001));
  INV_X1    g576(.A(new_n970), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(new_n968), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1000), .B(new_n1001), .C1(G1348), .C2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(new_n611), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT60), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT122), .B(new_n966), .C1(new_n994), .C2(new_n995), .ZN(new_n1007));
  OR3_X1    g582(.A1(new_n1004), .A2(KEYINPUT60), .A3(new_n610), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n998), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n992), .A3(new_n611), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n986), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n1012));
  INV_X1    g587(.A(G2090), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1003), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n960), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n958), .A2(KEYINPUT111), .A3(new_n959), .A4(new_n953), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1012), .B(new_n1014), .C1(new_n1018), .C2(G1971), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1971), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1014), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT112), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1019), .A2(G8), .A3(new_n1022), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n954), .A2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n954), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n585), .B2(new_n587), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n796), .A2(G1976), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n1028), .B(new_n1038), .C1(new_n951), .C2(new_n953), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT113), .B1(new_n954), .B2(G8), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT114), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  XNOR2_X1  g620(.A(G305), .B(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n594), .A2(KEYINPUT115), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G1981), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1046), .B(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1031), .A2(new_n1049), .A3(KEYINPUT116), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT116), .B1(new_n1031), .B2(new_n1049), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n974), .A2(new_n1013), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1020), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1024), .ZN(new_n1058));
  AND4_X1   g633(.A1(new_n1026), .A2(new_n1044), .A3(new_n1054), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2078), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1016), .A2(new_n1060), .A3(new_n1017), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1003), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n744), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n990), .A2(KEYINPUT53), .A3(new_n1060), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1063), .A2(G301), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT126), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n990), .A2(new_n1069), .A3(new_n1060), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT125), .B1(new_n960), .B2(G2078), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(KEYINPUT53), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1063), .A2(new_n1065), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1061), .A2(new_n1062), .B1(new_n744), .B2(new_n1064), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(G301), .A4(new_n1066), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1068), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n960), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(new_n712), .A3(new_n953), .A4(new_n970), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1038), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G286), .A2(G8), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1085), .A2(KEYINPUT51), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(KEYINPUT123), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  NAND3_X1  g666(.A1(G286), .A2(new_n1091), .A3(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1003), .A2(new_n712), .B1(new_n960), .B2(new_n1081), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(new_n1038), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT124), .B1(new_n1096), .B2(KEYINPUT51), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1084), .B1(new_n990), .B2(G1966), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1093), .B1(new_n1098), .B2(G8), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1089), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1095), .A2(new_n1086), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1073), .B2(G171), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1075), .A2(new_n1066), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1075), .A2(KEYINPUT127), .A3(G301), .A4(new_n1072), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(KEYINPUT54), .A4(new_n1111), .ZN(new_n1112));
  AND4_X1   g687(.A1(new_n1059), .A2(new_n1080), .A3(new_n1106), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1011), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1115), .A3(new_n1105), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1100), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT124), .B(KEYINPUT51), .C1(new_n1085), .C2(new_n1093), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1088), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT62), .B1(new_n1119), .B2(new_n1104), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1074), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1116), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1085), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1123), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1059), .ZN(new_n1126));
  NOR4_X1   g701(.A1(new_n1026), .A2(new_n1053), .A3(new_n1043), .A4(new_n1037), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1054), .A2(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(G305), .A2(G1981), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1053), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1019), .A2(G8), .A3(new_n1022), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1024), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1123), .A2(G286), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1132), .A2(new_n1134), .A3(new_n1026), .A4(new_n1135), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1127), .B(new_n1131), .C1(KEYINPUT63), .C2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1114), .A2(new_n1126), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n958), .A2(new_n989), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n792), .A2(new_n794), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n773), .B(G2067), .Z(new_n1141));
  INV_X1    g716(.A(G1996), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n738), .B(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n792), .A2(new_n794), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(G290), .B(G1986), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1139), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1139), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n792), .A2(new_n794), .A3(new_n1141), .A4(new_n1143), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n773), .A2(G2067), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1141), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1139), .B1(new_n1153), .B2(new_n738), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT46), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1149), .B2(G1996), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1139), .A2(KEYINPUT46), .A3(new_n1142), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT47), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1145), .A2(new_n1139), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1149), .A2(G290), .A3(G1986), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT48), .Z(new_n1162));
  AOI211_X1 g737(.A(new_n1152), .B(new_n1159), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1148), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(new_n929), .ZN(new_n1166));
  NAND3_X1  g740(.A1(new_n1166), .A2(new_n918), .A3(new_n930), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n1167), .A2(new_n941), .A3(new_n884), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n1168), .A2(KEYINPUT43), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n933), .A2(new_n945), .A3(new_n939), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n651), .A2(G319), .ZN(new_n1172));
  AOI211_X1 g746(.A(G227), .B(new_n1172), .C1(new_n890), .C2(new_n885), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n1171), .A2(new_n1173), .A3(new_n690), .ZN(G308));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1173), .A3(new_n690), .ZN(G225));
endmodule


