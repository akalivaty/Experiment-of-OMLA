//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(KEYINPUT73), .A3(G128), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n193), .B(new_n194), .C1(new_n190), .C2(G128), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n190), .A2(G128), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n191), .B(new_n199), .C1(new_n200), .C2(KEYINPUT23), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n197), .B1(G110), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G146), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n208), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n201), .A2(G110), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n216), .B(new_n217), .C1(new_n196), .C2(new_n195), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n220), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n223), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n213), .A2(new_n218), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n188), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n227), .A2(new_n228), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n189), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n226), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n189), .A2(G902), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n232), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n190), .A2(G116), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT2), .B(G113), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n237), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n242), .A2(new_n243), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(G137), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n257), .A2(G137), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n259), .A2(G134), .ZN(new_n265));
  OAI21_X1  g079(.A(G131), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT65), .B1(new_n211), .B2(G143), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G146), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT64), .A2(G143), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT64), .A2(G143), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n211), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n211), .A2(G143), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT1), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n273), .A2(new_n276), .B1(G128), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT64), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n271), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT64), .A2(G143), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(G146), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n211), .A2(KEYINPUT66), .A3(G143), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n287));
  AND4_X1   g101(.A1(new_n283), .A2(new_n285), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n268), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G131), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n263), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G146), .B1(new_n281), .B2(new_n282), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n269), .A2(new_n272), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n283), .A2(new_n293), .A3(new_n285), .A4(new_n286), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n255), .A2(new_n289), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G237), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n221), .A3(G210), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT27), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT26), .B(G101), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT69), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n301), .A2(new_n309), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n312));
  AND3_X1   g126(.A1(new_n292), .A2(new_n298), .A3(new_n299), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n278), .A2(G128), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n296), .B2(new_n297), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n283), .A2(new_n285), .A3(new_n286), .A4(new_n287), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n267), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT30), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n289), .A2(new_n300), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n255), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT68), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n324));
  AOI211_X1 g138(.A(new_n324), .B(new_n255), .C1(new_n318), .C2(new_n320), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n311), .B(new_n312), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n301), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n301), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n255), .B1(new_n289), .B2(new_n300), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n328), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n306), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n320), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n319), .B1(new_n289), .B2(new_n300), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n322), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n324), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n321), .A2(KEYINPUT68), .A3(new_n322), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n340), .A2(new_n341), .B1(new_n308), .B2(new_n310), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n326), .B(new_n336), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(G472), .A2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT32), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT32), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n328), .B1(new_n331), .B2(new_n327), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n306), .A2(KEYINPUT29), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n188), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT72), .B(new_n188), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n329), .B1(new_n340), .B2(new_n341), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n306), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n334), .B2(new_n335), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n355), .B(new_n356), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G472), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n236), .B1(new_n350), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n364));
  INV_X1    g178(.A(G475), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n188), .ZN(new_n366));
  XNOR2_X1  g180(.A(G113), .B(G122), .ZN(new_n367));
  INV_X1    g181(.A(G104), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G214), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n370), .A2(G237), .A3(G953), .ZN(new_n371));
  AOI21_X1  g185(.A(G143), .B1(KEYINPUT64), .B2(KEYINPUT81), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT81), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n204), .A2(new_n206), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G146), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n375), .A2(new_n376), .B1(new_n212), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n281), .A2(new_n380), .A3(new_n282), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n302), .A2(new_n221), .A3(G214), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n383), .A2(KEYINPUT18), .A3(G131), .A4(new_n373), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n383), .A2(G131), .A3(new_n373), .ZN(new_n386));
  AOI21_X1  g200(.A(G131), .B1(new_n383), .B2(new_n373), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT17), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(G131), .A3(new_n373), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n209), .B(new_n215), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n369), .B(new_n385), .C1(new_n388), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT83), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n375), .A2(new_n261), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n390), .A3(new_n389), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n395), .A2(new_n396), .A3(new_n209), .A4(new_n215), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n369), .A4(new_n385), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n401));
  INV_X1    g215(.A(new_n369), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n389), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT19), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n377), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n406));
  AOI21_X1  g220(.A(G146), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n209), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n379), .A2(new_n384), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n401), .B(new_n402), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n403), .A2(new_n409), .B1(new_n379), .B2(new_n384), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT82), .B1(new_n413), .B2(new_n369), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n366), .B1(new_n400), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n364), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n399), .A2(new_n393), .B1(new_n412), .B2(new_n414), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT84), .B(KEYINPUT20), .C1(new_n419), .C2(new_n366), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n417), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n397), .A2(new_n385), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n402), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n426), .A3(new_n402), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n400), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n365), .B1(new_n428), .B2(new_n188), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n422), .A2(KEYINPUT86), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT86), .B1(new_n422), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n274), .A2(new_n275), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G128), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n271), .A2(G128), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n257), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G122), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G116), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n246), .A2(G122), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G107), .ZN(new_n442));
  INV_X1    g256(.A(G107), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n437), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n434), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n274), .A2(new_n275), .A3(new_n198), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(KEYINPUT88), .A3(KEYINPUT13), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n435), .A2(new_n448), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT87), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n449), .A2(new_n452), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n446), .B1(new_n457), .B2(G134), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n246), .A2(KEYINPUT14), .A3(G122), .ZN(new_n459));
  OAI211_X1 g273(.A(G107), .B(new_n459), .C1(new_n441), .C2(KEYINPUT14), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n459), .A2(G107), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(KEYINPUT89), .C1(KEYINPUT14), .C2(new_n441), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n444), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G134), .B1(new_n453), .B2(new_n435), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n437), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT9), .B(G234), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n470), .A2(new_n187), .A3(G953), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n469), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n472), .A2(new_n473), .A3(new_n188), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n469), .A2(new_n471), .ZN(new_n481));
  INV_X1    g295(.A(new_n471), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n458), .A2(new_n468), .A3(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n473), .B(new_n188), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n478), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G952), .ZN(new_n488));
  AOI211_X1 g302(.A(G953), .B(new_n488), .C1(G234), .C2(G237), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n188), .B(new_n221), .C1(G234), .C2(G237), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT21), .B(G898), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n431), .A2(new_n432), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n315), .A2(new_n316), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(G125), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G224), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G953), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n298), .A2(new_n299), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n500), .B(new_n504), .C1(new_n505), .C2(new_n205), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT3), .B1(new_n368), .B2(G107), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT3), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n443), .A3(G104), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n368), .A2(G107), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G101), .ZN(new_n512));
  INV_X1    g326(.A(G101), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n507), .A2(new_n509), .A3(new_n513), .A4(new_n510), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n516), .A3(G101), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n251), .A2(new_n515), .A3(new_n517), .A4(new_n254), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n238), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n250), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n368), .A2(G107), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n443), .A2(G104), .ZN(new_n524));
  OAI21_X1  g338(.A(G101), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n514), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G110), .B(G122), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n518), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n505), .A2(new_n205), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n531), .A2(new_n499), .B1(new_n503), .B2(new_n502), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n506), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n534), .B(new_n535), .C1(new_n527), .C2(new_n522), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n529), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n502), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n500), .B(new_n541), .C1(new_n505), .C2(new_n205), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n502), .B1(new_n531), .B2(new_n499), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n529), .B(KEYINPUT77), .Z(new_n546));
  INV_X1    g360(.A(KEYINPUT76), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n518), .A2(new_n547), .A3(new_n528), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n518), .B2(new_n528), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n530), .A2(KEYINPUT6), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(KEYINPUT6), .B(new_n546), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n545), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n540), .B1(new_n554), .B2(KEYINPUT78), .ZN(new_n555));
  INV_X1    g369(.A(new_n546), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n518), .A2(new_n528), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT76), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n518), .A2(new_n547), .A3(new_n528), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n551), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n553), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n562), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n497), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n544), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n554), .A2(KEYINPUT78), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n496), .A4(new_n540), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT75), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G221), .ZN(new_n574));
  INV_X1    g388(.A(new_n470), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n188), .ZN(new_n576));
  INV_X1    g390(.A(G469), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n188), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n198), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n316), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n527), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n292), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n498), .A2(KEYINPUT10), .A3(new_n527), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n515), .A2(new_n517), .A3(new_n298), .A4(new_n299), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT1), .ZN(new_n590));
  OAI21_X1  g404(.A(G128), .B1(new_n296), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n579), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n526), .B1(new_n592), .B2(new_n316), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n587), .B(new_n588), .C1(new_n593), .C2(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n292), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(G110), .B(G140), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n221), .A2(G227), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n315), .A2(new_n526), .A3(new_n316), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n586), .B1(new_n583), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT12), .ZN(new_n604));
  INV_X1    g418(.A(new_n602), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n292), .B1(new_n593), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT12), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n601), .B(new_n589), .C1(new_n604), .C2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n578), .B1(new_n610), .B2(new_n577), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n589), .B1(new_n604), .B2(new_n608), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n599), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n601), .B1(new_n594), .B2(new_n292), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT74), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT74), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n589), .A2(new_n616), .A3(new_n601), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n617), .A3(new_n595), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n613), .A2(new_n618), .A3(G469), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n576), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n570), .A2(new_n573), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n363), .A2(new_n495), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  NAND2_X1  g437(.A1(new_n344), .A2(new_n188), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(G472), .ZN(new_n625));
  INV_X1    g439(.A(new_n236), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(new_n620), .A3(new_n626), .A4(new_n346), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n481), .A2(new_n483), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT33), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G478), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n474), .A2(new_n188), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n629), .A2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n474), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n422), .A2(new_n430), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT86), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n422), .A2(KEYINPUT86), .A3(new_n430), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n572), .B(new_n492), .C1(new_n564), .C2(new_n569), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n628), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n430), .A2(new_n486), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n418), .A2(new_n420), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT92), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT92), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n418), .A2(new_n648), .A3(new_n420), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n645), .B1(new_n650), .B2(new_n421), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n628), .A2(new_n641), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n625), .A2(new_n346), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n223), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n219), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n234), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n232), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT93), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n232), .A2(KEYINPUT93), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n495), .A2(new_n621), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT94), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(G12));
  AOI21_X1  g482(.A(new_n663), .B1(new_n350), .B2(new_n362), .ZN(new_n669));
  INV_X1    g483(.A(new_n489), .ZN(new_n670));
  INV_X1    g484(.A(new_n490), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(G900), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n669), .A2(new_n621), .A3(new_n651), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XNOR2_X1  g488(.A(new_n570), .B(KEYINPUT38), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n638), .A2(new_n639), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n331), .A2(new_n306), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n188), .B1(new_n342), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G472), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n350), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n659), .A2(new_n487), .A3(new_n572), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n675), .A2(new_n676), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT95), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(KEYINPUT95), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n603), .A2(KEYINPUT12), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n606), .A2(new_n607), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n614), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n601), .B1(new_n589), .B2(new_n595), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n577), .B(new_n188), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n578), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n619), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n576), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n672), .B(KEYINPUT39), .Z(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT40), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n683), .A2(new_n684), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(new_n433), .Z(G45));
  INV_X1    g512(.A(new_n635), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n699), .B(new_n672), .C1(new_n431), .C2(new_n432), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(KEYINPUT96), .A3(new_n621), .A4(new_n669), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT96), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n344), .A2(new_n348), .A3(new_n345), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n348), .B1(new_n344), .B2(new_n345), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n362), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n661), .A2(new_n662), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n572), .B1(new_n564), .B2(new_n569), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n620), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n703), .B1(new_n709), .B2(new_n700), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n702), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NOR2_X1   g526(.A1(new_n687), .A2(new_n688), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n713), .B2(G902), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n714), .A2(new_n692), .A3(new_n689), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n363), .A2(new_n640), .A3(new_n641), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n363), .A2(new_n641), .A3(new_n651), .A4(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  INV_X1    g534(.A(KEYINPUT97), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n721), .A2(new_n570), .A3(new_n573), .A4(new_n715), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n708), .B2(new_n715), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n495), .B(new_n669), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND2_X1  g539(.A1(new_n351), .A2(new_n335), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n326), .B(new_n726), .C1(new_n342), .C2(new_n343), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n345), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n625), .A2(new_n626), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT98), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n624), .A2(G472), .B1(new_n727), .B2(new_n345), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(KEYINPUT98), .A3(new_n626), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n431), .A2(new_n432), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n570), .A2(new_n573), .A3(new_n486), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n715), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n492), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  AND3_X1   g555(.A1(new_n625), .A2(new_n659), .A3(new_n728), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n701), .B(new_n742), .C1(new_n722), .C2(new_n723), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  NAND2_X1  g558(.A1(new_n706), .A2(new_n626), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n564), .A2(new_n573), .A3(new_n569), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT99), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n693), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n691), .A2(KEYINPUT99), .A3(new_n692), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n747), .A2(new_n701), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT100), .ZN(new_n754));
  INV_X1    g568(.A(new_n746), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n706), .A3(new_n755), .A4(new_n626), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n754), .B(KEYINPUT42), .C1(new_n756), .C2(new_n700), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n261), .ZN(G33));
  NAND2_X1  g573(.A1(new_n651), .A2(new_n672), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n257), .ZN(G36));
  NAND2_X1  g576(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n676), .A2(new_n635), .ZN(new_n765));
  MUX2_X1   g579(.A(new_n763), .B(new_n764), .S(new_n765), .Z(new_n766));
  NAND2_X1  g580(.A1(new_n655), .A2(new_n659), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT102), .Z(new_n768));
  AOI21_X1  g582(.A(KEYINPUT44), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(KEYINPUT44), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n755), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT103), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT45), .B1(new_n613), .B2(new_n618), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n577), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n613), .A2(new_n618), .A3(KEYINPUT45), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n578), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n689), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n692), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(new_n694), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n773), .A2(KEYINPUT103), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n771), .A2(new_n774), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT105), .B(G137), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G39));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n781), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n706), .A2(new_n626), .A3(new_n746), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n701), .A3(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(KEYINPUT106), .B(G140), .Z(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(G42));
  AND2_X1   g609(.A1(new_n714), .A2(new_n689), .ZN(new_n796));
  NAND2_X1  g610(.A1(KEYINPUT107), .A2(KEYINPUT49), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(KEYINPUT107), .B2(KEYINPUT49), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n573), .A3(new_n692), .A4(new_n626), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n798), .A2(KEYINPUT107), .A3(KEYINPUT49), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n680), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n675), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n765), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n699), .B1(new_n431), .B2(new_n432), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n638), .A2(new_n639), .A3(new_n486), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n708), .A2(new_n493), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n627), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n740), .A2(new_n724), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n716), .A2(new_n719), .A3(new_n622), .A4(new_n665), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n758), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n649), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n648), .B1(new_n418), .B2(new_n420), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n421), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n487), .A2(new_n430), .A3(new_n672), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n693), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n706), .A2(new_n707), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n742), .A2(new_n751), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n820), .B2(new_n700), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n755), .ZN(new_n822));
  INV_X1    g636(.A(new_n761), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT108), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT108), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n640), .A2(new_n672), .A3(new_n742), .A4(new_n751), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n746), .B1(new_n826), .B2(new_n819), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n827), .B2(new_n761), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n813), .A2(KEYINPUT53), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n672), .B(KEYINPUT111), .Z(new_n831));
  OR2_X1    g645(.A1(new_n659), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT112), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n737), .A2(new_n833), .A3(new_n620), .A4(new_n680), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n711), .A2(new_n673), .A3(new_n743), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n722), .A2(new_n723), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n640), .A2(new_n672), .A3(new_n742), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n673), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n743), .A2(KEYINPUT110), .A3(new_n673), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n711), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n837), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n837), .B2(new_n845), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n830), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n811), .A2(new_n812), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n753), .A2(new_n757), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n828), .A4(new_n824), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT109), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n813), .A2(KEYINPUT109), .A3(new_n824), .A4(new_n828), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n835), .A2(new_n836), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n855), .A2(new_n856), .B1(new_n837), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n849), .B(new_n850), .C1(new_n858), .C2(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n856), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n847), .A2(new_n848), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n862), .A2(new_n863), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n859), .B1(new_n864), .B2(new_n850), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n766), .A2(new_n489), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(new_n734), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(KEYINPUT115), .A3(new_n755), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n734), .A3(new_n755), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n796), .A2(new_n576), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n789), .A2(new_n790), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n876), .A2(KEYINPUT51), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n738), .A2(new_n746), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n742), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n626), .A2(new_n489), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n680), .A2(new_n738), .A3(new_n746), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n735), .A3(new_n635), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n675), .A2(new_n573), .A3(new_n738), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n868), .A2(new_n734), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n889), .A2(KEYINPUT118), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(KEYINPUT118), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n877), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT114), .B(new_n859), .C1(new_n864), .C2(new_n850), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n791), .A2(KEYINPUT116), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n791), .A2(KEYINPUT116), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n874), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n870), .B(new_n873), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT51), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n868), .A2(new_n363), .A3(new_n878), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT48), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n869), .B1(new_n722), .B2(new_n723), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n488), .B(G953), .C1(new_n881), .C2(new_n640), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n867), .A2(new_n892), .A3(new_n893), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT119), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n804), .B1(new_n905), .B2(new_n907), .ZN(G75));
  OAI21_X1  g722(.A(new_n849), .B1(new_n858), .B2(KEYINPUT53), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(G210), .A3(G902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n562), .B(new_n544), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n221), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  XOR2_X1   g732(.A(new_n713), .B(KEYINPUT120), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n859), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n578), .B(KEYINPUT57), .Z(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n909), .A2(G902), .A3(new_n777), .A4(new_n776), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT121), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n917), .B1(new_n924), .B2(new_n926), .ZN(G54));
  INV_X1    g741(.A(new_n917), .ZN(new_n928));
  AND4_X1   g742(.A1(KEYINPUT58), .A2(new_n909), .A3(G475), .A4(G902), .ZN(new_n929));
  INV_X1    g743(.A(new_n419), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n930), .B2(new_n929), .ZN(G60));
  INV_X1    g746(.A(new_n630), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n867), .A2(new_n893), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n632), .B(KEYINPUT59), .Z(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n935), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n921), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g754(.A(KEYINPUT122), .B(new_n938), .C1(new_n920), .C2(new_n859), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n928), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n936), .A2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT60), .Z(new_n945));
  AND3_X1   g759(.A1(new_n909), .A2(KEYINPUT123), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT123), .B1(new_n909), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n657), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n857), .A2(new_n837), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT53), .B1(new_n860), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n848), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n837), .A2(new_n845), .A3(new_n846), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n829), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n945), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n909), .A2(KEYINPUT123), .A3(new_n945), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n233), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n948), .A2(new_n928), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n948), .A2(new_n958), .A3(KEYINPUT61), .A4(new_n928), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G66));
  INV_X1    g777(.A(new_n851), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n221), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n491), .B2(new_n501), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(KEYINPUT124), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(KEYINPUT124), .B2(new_n965), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n552), .B(new_n553), .C1(G898), .C2(new_n221), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(G69));
  AND3_X1   g784(.A1(new_n842), .A2(new_n711), .A3(new_n844), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n697), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n747), .A2(new_n695), .A3(new_n807), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT125), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n793), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n785), .A2(new_n973), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n221), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n405), .A2(new_n406), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n321), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(G900), .B2(G953), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n745), .A2(new_n735), .A3(new_n736), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n761), .B1(new_n783), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n793), .A2(new_n986), .A3(new_n852), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n785), .A2(new_n971), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n984), .B1(new_n988), .B2(G953), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n221), .B1(G227), .B2(G900), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n983), .A2(new_n992), .A3(new_n991), .A4(new_n989), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n988), .B2(new_n964), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n357), .A2(new_n335), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n917), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n999), .B1(new_n358), .B2(new_n342), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n864), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n999), .B1(new_n978), .B2(new_n964), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n357), .A2(new_n335), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(G57));
endmodule


