//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G116), .C2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  OAI21_X1  g0017(.A(KEYINPUT64), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OR3_X1    g0018(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT64), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n222), .A2(new_n217), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(new_n218), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NOR3_X1   g0028(.A1(new_n221), .A2(new_n224), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G222), .A2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G223), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G77), .B2(new_n250), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT66), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n216), .A2(new_n266), .B1(new_n267), .B2(new_n257), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n268), .B2(G226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G190), .ZN(new_n272));
  XOR2_X1   g0072(.A(KEYINPUT8), .B(G58), .Z(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT68), .B1(new_n247), .B2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(new_n217), .A3(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n273), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n203), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n279), .B(new_n280), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT67), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(new_n223), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n285), .A3(new_n223), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n286), .A2(new_n285), .A3(new_n223), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n216), .A2(G20), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n216), .A2(G13), .A3(G20), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n291), .B(new_n296), .C1(G50), .C2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n270), .A2(G200), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n272), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n272), .A2(new_n301), .A3(KEYINPUT70), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(G190), .A2(new_n271), .B1(new_n299), .B2(new_n300), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n302), .C1(KEYINPUT70), .C2(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n270), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(new_n298), .C1(G179), .C2(new_n270), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G238), .A2(G1698), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n250), .B(new_n314), .C1(new_n213), .C2(G1698), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n259), .C1(G107), .C2(new_n250), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n266), .A2(new_n216), .A3(G274), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n268), .A2(G244), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G20), .A2(G77), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n217), .A2(G33), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  INV_X1    g0125(.A(new_n273), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n282), .B(KEYINPUT69), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n323), .B1(new_n324), .B2(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n290), .B1(new_n295), .B2(G77), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(G77), .B2(new_n297), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n319), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(G190), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n319), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n334), .B2(new_n330), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n310), .A2(new_n313), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n211), .A2(G1698), .ZN(new_n338));
  AND2_X1   g0138(.A1(G232), .A2(G1698), .ZN(new_n339));
  AND2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NOR2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n258), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n258), .A2(G238), .A3(new_n261), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n317), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT13), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n252), .A2(G226), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G232), .A2(G1698), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n248), .A2(new_n249), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n343), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n259), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n263), .B1(new_n268), .B2(G238), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT72), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n347), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT72), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G179), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n354), .B1(new_n352), .B2(new_n353), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT13), .ZN(new_n362));
  OAI21_X1  g0162(.A(G169), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(new_n355), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(G169), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n360), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n288), .A2(G68), .A3(new_n289), .A4(new_n294), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT74), .B1(new_n297), .B2(G68), .ZN(new_n370));
  INV_X1    g0170(.A(G13), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(G1), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT74), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(G20), .A4(new_n207), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n374), .A3(KEYINPUT12), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT12), .ZN(new_n376));
  OAI211_X1 g0176(.A(KEYINPUT74), .B(new_n376), .C1(new_n297), .C2(G68), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n369), .A2(new_n375), .A3(KEYINPUT75), .A4(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n369), .A2(new_n375), .A3(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g0181(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G77), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n274), .B2(new_n277), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n283), .A2(new_n202), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n217), .A2(G68), .ZN(new_n387));
  OR3_X1    g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n383), .B1(new_n388), .B2(new_n290), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n390), .A2(new_n293), .A3(new_n382), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n378), .B(new_n381), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(G190), .B2(new_n359), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n347), .B2(new_n355), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT71), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n368), .A2(new_n392), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n248), .A2(new_n217), .A3(new_n249), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n249), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n207), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n212), .A2(new_n207), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n404), .B2(new_n201), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n282), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n398), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n340), .A2(new_n341), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(new_n217), .ZN(new_n410));
  INV_X1    g0210(.A(new_n402), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n407), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n414), .A3(new_n290), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n326), .A2(new_n297), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n295), .B2(new_n326), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(G223), .A2(G1698), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n211), .A2(G1698), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n340), .C2(new_n341), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G87), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n259), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n263), .B1(new_n268), .B2(G232), .ZN(new_n425));
  AOI21_X1  g0225(.A(G169), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n321), .A3(new_n425), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n424), .A2(KEYINPUT76), .A3(new_n321), .A4(new_n425), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n418), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT77), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n418), .A2(new_n431), .A3(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(KEYINPUT77), .A3(new_n433), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n424), .A2(G190), .A3(new_n425), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n424), .A2(new_n425), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G200), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n415), .A2(new_n417), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT17), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n397), .A2(new_n437), .A3(new_n438), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n337), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n208), .A2(new_n252), .ZN(new_n446));
  INV_X1    g0246(.A(G244), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G1698), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n448), .C1(new_n340), .C2(new_n341), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n247), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n258), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n216), .A2(G45), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n262), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n258), .A2(G250), .A3(new_n454), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n453), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G179), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n458), .B2(new_n311), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT79), .ZN(new_n461));
  INV_X1    g0261(.A(G87), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  INV_X1    g0263(.A(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n343), .A2(new_n217), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT19), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n217), .B(G68), .C1(new_n340), .C2(new_n341), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT19), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n324), .B2(new_n463), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n297), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n471), .A2(new_n290), .B1(new_n472), .B2(new_n325), .ZN(new_n473));
  INV_X1    g0273(.A(new_n325), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n216), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n293), .A2(new_n297), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n461), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n461), .A3(new_n476), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n460), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n453), .ZN(new_n481));
  INV_X1    g0281(.A(new_n455), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n456), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G200), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n458), .A2(G190), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n293), .A2(G87), .A3(new_n297), .A4(new_n475), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n473), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n217), .B2(G107), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n464), .A2(KEYINPUT23), .A3(G20), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n491), .B1(new_n451), .B2(new_n217), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n217), .B(G87), .C1(new_n340), .C2(new_n341), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT24), .B(new_n492), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n290), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT83), .A4(new_n290), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n293), .A2(new_n297), .A3(new_n475), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(new_n464), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n372), .A2(G20), .A3(new_n464), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT25), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(G257), .B(G1698), .C1(new_n340), .C2(new_n341), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT84), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n250), .A2(new_n514), .A3(G257), .A4(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G294), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n250), .A2(G250), .A3(new_n252), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n259), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G41), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n455), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n522), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n258), .B1(new_n525), .B2(new_n454), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n527), .B2(G264), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G169), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n321), .B2(new_n529), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n488), .B1(new_n511), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n472), .A2(new_n463), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n506), .B2(new_n463), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n283), .A2(new_n384), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n464), .A2(KEYINPUT6), .A3(G97), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  XNOR2_X1  g0339(.A(G97), .B(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(KEYINPUT78), .B(new_n536), .C1(new_n541), .C2(new_n217), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT78), .ZN(new_n543));
  AND2_X1   g0343(.A1(G97), .A2(G107), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n217), .B1(new_n546), .B2(new_n537), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n535), .ZN(new_n548));
  OAI21_X1  g0348(.A(G107), .B1(new_n410), .B2(new_n411), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n534), .B1(new_n550), .B2(new_n290), .ZN(new_n551));
  OAI21_X1  g0351(.A(G244), .B1(new_n340), .B2(new_n341), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G283), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n553), .A2(G1698), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(G244), .C1(new_n341), .C2(new_n340), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(G250), .B1(new_n340), .B2(new_n341), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n252), .B1(new_n559), .B2(KEYINPUT4), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n259), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G257), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n523), .B1(new_n526), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n559), .A2(KEYINPUT4), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G1698), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n552), .A2(new_n553), .B1(G33), .B2(G283), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n557), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n563), .B1(new_n570), .B2(new_n259), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G190), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n551), .A2(new_n566), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n565), .A2(new_n311), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n321), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n573), .B1(new_n576), .B2(new_n551), .ZN(new_n577));
  INV_X1    g0377(.A(new_n510), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n503), .B2(new_n504), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n529), .A2(new_n394), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G190), .B2(new_n529), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n577), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n562), .A2(new_n252), .ZN(new_n583));
  INV_X1    g0383(.A(G264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G1698), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n585), .C1(new_n340), .C2(new_n341), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n248), .A2(G303), .A3(new_n249), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT80), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT80), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n259), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n527), .A2(G270), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n523), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n286), .A2(new_n223), .B1(G20), .B2(new_n450), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n555), .B(new_n217), .C1(G33), .C2(new_n463), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(KEYINPUT81), .B2(KEYINPUT20), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(KEYINPUT81), .B2(KEYINPUT20), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n293), .A2(G116), .A3(new_n297), .A4(new_n475), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n372), .A2(G20), .A3(new_n450), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT81), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n595), .A2(new_n601), .A3(new_n596), .A4(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n594), .A2(G169), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n594), .A2(new_n607), .A3(G169), .A4(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n592), .A2(new_n593), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(G179), .A3(new_n523), .A4(new_n604), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n594), .A2(G200), .ZN(new_n612));
  INV_X1    g0412(.A(new_n604), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n333), .C2(new_n594), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n609), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n445), .A2(new_n532), .A3(new_n582), .A4(new_n615), .ZN(G372));
  AND2_X1   g0416(.A1(new_n434), .A2(new_n436), .ZN(new_n617));
  INV_X1    g0417(.A(new_n392), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n359), .A2(G190), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n395), .A2(KEYINPUT71), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n395), .A2(KEYINPUT71), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n331), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n364), .A2(new_n367), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n321), .B1(new_n357), .B2(new_n358), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n392), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n617), .B1(new_n628), .B2(new_n443), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n313), .B1(new_n309), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT86), .Z(new_n631));
  NOR2_X1   g0431(.A1(new_n529), .A2(new_n321), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(G169), .B2(new_n529), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n609), .B(new_n611), .C1(new_n579), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n579), .A2(new_n581), .ZN(new_n635));
  INV_X1    g0435(.A(new_n577), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n473), .A2(new_n476), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n458), .A2(new_n311), .ZN(new_n638));
  NOR4_X1   g0438(.A1(new_n453), .A2(new_n457), .A3(new_n321), .A4(new_n455), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n487), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT85), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n561), .A2(new_n321), .A3(new_n564), .ZN(new_n644));
  AOI21_X1  g0444(.A(G169), .B1(new_n561), .B2(new_n564), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n550), .A2(new_n290), .ZN(new_n647));
  INV_X1    g0447(.A(new_n534), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n646), .A2(new_n649), .A3(new_n487), .A4(new_n640), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n640), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n473), .A2(new_n461), .A3(new_n476), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n477), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n458), .A2(new_n394), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n473), .A2(new_n486), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n654), .A2(new_n460), .B1(new_n657), .B2(new_n485), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n551), .A2(new_n644), .A3(new_n645), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n643), .B1(new_n651), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n646), .A2(new_n649), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT26), .B1(new_n488), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n641), .A2(new_n659), .A3(new_n652), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(KEYINPUT85), .A3(new_n664), .A4(new_n640), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n642), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n445), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n631), .A2(new_n667), .ZN(G369));
  NOR2_X1   g0468(.A1(new_n371), .A2(G20), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n216), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n615), .B1(new_n613), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n609), .A2(new_n611), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n613), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n511), .A2(new_n531), .A3(new_n675), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT88), .Z(new_n685));
  NAND2_X1  g0485(.A1(new_n511), .A2(new_n531), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n686), .B(new_n635), .C1(new_n579), .C2(new_n676), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n675), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n675), .B1(new_n609), .B2(new_n611), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n226), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n465), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n222), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n666), .A2(new_n676), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n666), .A2(KEYINPUT91), .A3(new_n676), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT92), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n634), .A2(new_n487), .A3(new_n635), .A4(new_n636), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n659), .A2(new_n652), .A3(new_n487), .A4(new_n480), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n640), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n708), .B1(new_n713), .B2(new_n676), .ZN(new_n714));
  AOI211_X1 g0514(.A(KEYINPUT92), .B(new_n675), .C1(new_n709), .C2(new_n712), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT29), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n565), .A2(new_n459), .ZN(new_n717));
  INV_X1    g0517(.A(new_n529), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n610), .A3(KEYINPUT30), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n571), .A2(new_n639), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n519), .A2(new_n592), .A3(new_n528), .A4(new_n593), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n483), .A2(KEYINPUT89), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT89), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n458), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n321), .A3(new_n565), .A4(new_n594), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n719), .B(new_n723), .C1(new_n728), .C2(new_n718), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n675), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT90), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n582), .A2(new_n532), .A3(new_n615), .A4(new_n676), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT90), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n730), .A2(new_n735), .A3(new_n731), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n733), .A2(new_n734), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n707), .A2(new_n716), .B1(G330), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n701), .B1(new_n739), .B2(G1), .ZN(G364));
  INV_X1    g0540(.A(new_n683), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n216), .B1(new_n669), .B2(G45), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n697), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n741), .B(new_n743), .C1(G330), .C2(new_n681), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n743), .B(KEYINPUT93), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n695), .A2(new_n409), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G355), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n695), .A2(new_n250), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G45), .B2(new_n222), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n241), .A2(new_n265), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n748), .B1(G116), .B2(new_n226), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n223), .B1(G20), .B2(new_n311), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n217), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(G20), .A2(G179), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT95), .Z(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n250), .B1(new_n462), .B2(new_n761), .C1(new_n765), .C2(new_n384), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n760), .A2(new_n764), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n770));
  XNOR2_X1  g0570(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n394), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n760), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n464), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n333), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n217), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n463), .ZN(new_n777));
  OR3_X1    g0577(.A1(new_n771), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n763), .A2(G190), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n394), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n766), .B(new_n778), .C1(G50), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n779), .A2(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT97), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n763), .A2(new_n784), .A3(new_n772), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(new_n763), .B2(new_n772), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n781), .B1(new_n212), .B2(new_n783), .C1(new_n207), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n776), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G329), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n409), .B1(new_n767), .B2(new_n792), .C1(new_n793), .C2(new_n773), .ZN(new_n794));
  INV_X1    g0594(.A(new_n765), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n791), .B(new_n794), .C1(new_n795), .C2(G311), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G322), .A2(new_n782), .B1(new_n780), .B2(G326), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  OAI221_X1 g0600(.A(new_n798), .B1(new_n799), .B2(new_n761), .C1(new_n788), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n789), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n756), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n746), .B(new_n759), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT98), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  INV_X1    g0607(.A(new_n755), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n807), .C1(new_n681), .C2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n744), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  XOR2_X1   g0611(.A(KEYINPUT100), .B(G143), .Z(new_n812));
  AOI22_X1  g0612(.A1(G137), .A2(new_n780), .B1(new_n782), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n813), .B1(new_n281), .B2(new_n788), .C1(new_n768), .C2(new_n765), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n250), .B1(new_n761), .B2(new_n202), .ZN(new_n817));
  INV_X1    g0617(.A(new_n767), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G132), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n816), .B(new_n819), .C1(new_n212), .C2(new_n776), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n773), .A2(new_n207), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n814), .A2(new_n815), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n409), .B1(new_n767), .B2(new_n824), .C1(new_n462), .C2(new_n773), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n777), .B(new_n825), .C1(new_n795), .C2(G116), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G294), .A2(new_n782), .B1(new_n780), .B2(G303), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(new_n793), .C2(new_n788), .ZN(new_n828));
  INV_X1    g0628(.A(new_n761), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(G107), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n756), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n756), .A2(new_n753), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n745), .B1(new_n384), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT99), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n623), .A2(KEYINPUT101), .A3(new_n675), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n330), .A2(new_n675), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n331), .B(new_n836), .C1(new_n334), .C2(new_n330), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT101), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n331), .B2(new_n676), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n835), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n831), .B(new_n834), .C1(new_n754), .C2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT102), .Z(new_n842));
  INV_X1    g0642(.A(new_n840), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n704), .A2(new_n706), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n666), .A2(new_n676), .A3(new_n840), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n738), .A2(G330), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n842), .B1(new_n851), .B2(new_n743), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  INV_X1    g0653(.A(KEYINPUT35), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n217), .B(new_n223), .C1(new_n541), .C2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n855), .B(G116), .C1(new_n854), .C2(new_n541), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  OAI21_X1  g0657(.A(G77), .B1(new_n212), .B2(new_n207), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n858), .A2(new_n222), .B1(G50), .B2(new_n207), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(G1), .A3(new_n371), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n734), .A2(new_n732), .A3(new_n737), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n368), .A2(new_n392), .A3(new_n675), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n392), .A2(new_n675), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n397), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n627), .A2(new_n622), .A3(new_n863), .A4(new_n864), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n862), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n868), .A3(new_n840), .ZN(new_n869));
  INV_X1    g0669(.A(new_n673), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n418), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n673), .B1(new_n415), .B2(new_n417), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n872), .A2(new_n432), .A3(new_n442), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n873), .B(KEYINPUT105), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n432), .A2(new_n442), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n878), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n442), .B(KEYINPUT17), .Z(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(new_n617), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n437), .A2(new_n443), .A3(new_n438), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n873), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n880), .B2(new_n873), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n869), .A2(KEYINPUT106), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n888), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n898), .A2(new_n896), .A3(new_n894), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n627), .A2(new_n622), .A3(new_n864), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT104), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n866), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n843), .B1(new_n902), .B2(new_n862), .ZN(new_n903));
  NAND2_X1  g0703(.A1(KEYINPUT106), .A2(KEYINPUT40), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n861), .A3(new_n904), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n895), .A2(new_n896), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT107), .Z(new_n907));
  NAND2_X1  g0707(.A1(new_n445), .A2(new_n861), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(G330), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n707), .A2(new_n445), .A3(new_n716), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n631), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n894), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n627), .A2(new_n675), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n617), .A2(new_n673), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n331), .A2(new_n675), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n846), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n898), .A2(new_n894), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n868), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n912), .B(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n910), .A2(new_n927), .B1(new_n216), .B2(new_n669), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT108), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n910), .A2(new_n927), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n857), .B(new_n860), .C1(new_n929), .C2(new_n930), .ZN(G367));
  OAI21_X1  g0731(.A(new_n636), .B1(new_n551), .B2(new_n676), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n659), .A2(new_n675), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n688), .A2(new_n692), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n662), .B1(new_n932), .B2(new_n686), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n676), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n656), .A2(new_n675), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n641), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n640), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n689), .A3(new_n934), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n689), .A2(new_n934), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n940), .A3(new_n944), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n947), .B1(new_n946), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n696), .B(KEYINPUT41), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT45), .B1(new_n693), .B2(new_n934), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT44), .ZN(new_n959));
  INV_X1    g0759(.A(new_n934), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n688), .A2(new_n692), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n691), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT44), .B1(new_n693), .B2(new_n934), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n689), .B1(new_n958), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n957), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n955), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n967), .A2(new_n690), .A3(new_n963), .A4(new_n962), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n688), .B(new_n692), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(new_n683), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n965), .A2(new_n968), .A3(new_n739), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n954), .B1(new_n971), .B2(new_n739), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n742), .B(KEYINPUT109), .Z(new_n973));
  OAI21_X1  g0773(.A(new_n952), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(G137), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n250), .B1(new_n767), .B2(new_n975), .C1(new_n212), .C2(new_n761), .ZN(new_n976));
  INV_X1    g0776(.A(new_n776), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(G68), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n765), .B2(new_n202), .ZN(new_n979));
  INV_X1    g0779(.A(new_n773), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n976), .B(new_n979), .C1(G77), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n780), .A2(new_n812), .ZN(new_n982));
  INV_X1    g0782(.A(new_n788), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(G159), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n782), .A2(G150), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n981), .A2(new_n982), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n780), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n799), .A2(new_n783), .B1(new_n987), .B2(new_n824), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n829), .A2(KEYINPUT46), .A3(G116), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n761), .B2(new_n450), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(new_n464), .C2(new_n776), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n818), .A2(G317), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n765), .B2(new_n793), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n988), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n463), .B2(new_n773), .C1(new_n790), .C2(new_n788), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n986), .B1(new_n996), .B2(new_n250), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n745), .B1(new_n998), .B2(new_n756), .ZN(new_n999));
  INV_X1    g0799(.A(new_n749), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n757), .B1(new_n226), .B2(new_n325), .C1(new_n1000), .C2(new_n237), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(new_n808), .C2(new_n943), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n974), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT110), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT110), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n974), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(G387));
  NAND2_X1  g0807(.A1(new_n829), .A2(G77), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n281), .B2(new_n767), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n250), .B1(new_n1009), .B2(KEYINPUT111), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1009), .A2(KEYINPUT111), .B1(G97), .B2(new_n980), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n325), .B2(new_n776), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G159), .C2(new_n780), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n788), .A2(new_n326), .B1(new_n207), .B2(new_n765), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT112), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(new_n202), .C2(new_n783), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT113), .Z(new_n1017));
  AOI22_X1  g0817(.A1(G317), .A2(new_n782), .B1(new_n780), .B2(G322), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n799), .B2(new_n765), .C1(new_n824), .C2(new_n788), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n793), .B2(new_n776), .C1(new_n790), .C2(new_n761), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n250), .B1(new_n818), .B2(G326), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n773), .A2(new_n450), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1017), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n745), .B1(new_n1028), .B2(new_n756), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n688), .B2(new_n808), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n234), .A2(new_n265), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n698), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1031), .A2(new_n749), .B1(new_n1032), .B2(new_n747), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n273), .A2(new_n202), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1032), .B1(new_n1034), .B2(KEYINPUT50), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n265), .C1(KEYINPUT50), .C2(new_n1034), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G68), .B2(G77), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1033), .A2(new_n1037), .B1(G107), .B2(new_n226), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1030), .B1(new_n758), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n970), .B2(new_n973), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n970), .A2(new_n739), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n696), .B1(new_n970), .B2(new_n739), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(G393));
  NAND2_X1  g0844(.A1(new_n965), .A2(new_n968), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n1041), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n971), .A3(new_n696), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n965), .A2(new_n968), .A3(new_n973), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n788), .A2(new_n202), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n250), .B1(new_n773), .B2(new_n462), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n818), .B2(new_n812), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n384), .B2(new_n776), .C1(new_n326), .C2(new_n765), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT51), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n281), .A2(new_n987), .B1(new_n783), .B2(new_n768), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1049), .B(new_n1052), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n1053), .B2(new_n1054), .C1(new_n207), .C2(new_n761), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G311), .A2(new_n782), .B1(new_n780), .B2(G317), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  AOI211_X1 g0858(.A(new_n250), .B(new_n774), .C1(G322), .C2(new_n818), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n450), .B2(new_n776), .C1(new_n790), .C2(new_n765), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G303), .B2(new_n983), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1058), .B(new_n1061), .C1(new_n793), .C2(new_n761), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n745), .B1(new_n1063), .B2(new_n756), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n757), .B1(new_n463), .B2(new_n226), .C1(new_n1000), .C2(new_n244), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n808), .C2(new_n934), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1048), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT115), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n1047), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1047), .B2(new_n1067), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(G390));
  NAND3_X1  g0872(.A1(new_n445), .A2(G330), .A3(new_n861), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n911), .A2(new_n631), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n713), .A2(new_n676), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(KEYINPUT92), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n713), .A2(new_n708), .A3(new_n676), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n921), .B1(new_n1078), .B2(new_n840), .ZN(new_n1079));
  INV_X1    g0879(.A(G330), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n843), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n868), .B1(new_n861), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n738), .A2(new_n1081), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1082), .B1(new_n1083), .B2(new_n868), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n861), .A2(new_n1081), .A3(new_n868), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1083), .B2(new_n868), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n923), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1074), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n918), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n914), .B2(new_n915), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n868), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n1079), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n923), .A2(new_n868), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1091), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n916), .A2(new_n917), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1095), .A2(new_n868), .A3(new_n1099), .A4(new_n1083), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n840), .B1(new_n714), .B2(new_n715), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n922), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1092), .B1(new_n1102), .B2(new_n868), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1096), .A2(new_n1091), .B1(new_n916), .B2(new_n917), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1086), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1090), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1079), .A2(new_n1084), .B1(new_n1087), .B2(new_n923), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n911), .A2(new_n631), .A3(new_n1073), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1086), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n738), .A2(new_n868), .A3(new_n1081), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1103), .A2(new_n1104), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1109), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1106), .A2(new_n696), .A3(new_n1114), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n273), .A2(new_n756), .A3(new_n753), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n450), .A2(new_n783), .B1(new_n987), .B2(new_n793), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G77), .B2(new_n977), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n409), .B1(new_n767), .B2(new_n790), .C1(new_n462), .C2(new_n761), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n821), .B(new_n1119), .C1(new_n795), .C2(G97), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(new_n464), .C2(new_n788), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n409), .B1(new_n980), .B2(G50), .ZN(new_n1122));
  INV_X1    g0922(.A(G125), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n767), .C1(new_n768), .C2(new_n776), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT54), .B(G143), .Z(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n795), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n983), .A2(G137), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G128), .A2(new_n780), .B1(new_n782), .B2(G132), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n761), .A2(new_n281), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1121), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n746), .B1(new_n1132), .B2(new_n803), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1116), .B(new_n1133), .C1(new_n1098), .C2(new_n753), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n973), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1115), .A2(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(KEYINPUT120), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n313), .ZN(new_n1139));
  OR3_X1    g0939(.A1(new_n309), .A2(KEYINPUT55), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT55), .B1(new_n309), .B2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n298), .A2(new_n870), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT56), .Z(new_n1143));
  AND3_X1   g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n926), .A2(G330), .A3(new_n906), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT106), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n903), .B2(new_n861), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n914), .A2(new_n915), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT40), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n898), .A2(new_n896), .A3(new_n894), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n869), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n904), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1080), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(new_n926), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1147), .B1(new_n1148), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n906), .A2(G330), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n926), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1156), .A2(new_n926), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n1146), .A3(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1074), .A2(new_n1114), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1138), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n697), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1108), .B1(new_n1135), .B2(new_n1109), .ZN(new_n1169));
  OAI211_X1 g0969(.A(KEYINPUT120), .B(new_n1167), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1146), .A2(new_n753), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n832), .A2(new_n202), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G58), .A2(new_n980), .B1(new_n818), .B2(G283), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n978), .A3(new_n1008), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n782), .A2(G107), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT116), .Z(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G116), .C2(new_n780), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n788), .A2(new_n463), .B1(new_n325), .B2(new_n765), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT117), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1178), .A2(new_n264), .A3(new_n409), .A4(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n202), .B1(new_n340), .B2(G41), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n776), .A2(new_n281), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n795), .A2(G137), .B1(new_n829), .B2(new_n1125), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n782), .A2(G128), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n1123), .C2(new_n987), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1185), .B(new_n1188), .C1(G132), .C2(new_n983), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT59), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G41), .B1(new_n818), .B2(G124), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G33), .B1(new_n980), .B2(G159), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1183), .A2(new_n1184), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n743), .B1(new_n1194), .B2(new_n756), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1172), .A2(new_n1173), .A3(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT119), .Z(new_n1197));
  INV_X1    g0997(.A(new_n1168), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n973), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1171), .A2(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n832), .A2(new_n207), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n868), .A2(new_n754), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n776), .A2(new_n325), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n409), .B1(new_n773), .B2(new_n384), .C1(new_n463), .C2(new_n761), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G107), .C2(new_n795), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G283), .A2(new_n782), .B1(new_n780), .B2(G294), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n450), .B2(new_n788), .C1(new_n799), .C2(new_n767), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n983), .A2(new_n1125), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n818), .A2(G128), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G132), .A2(new_n780), .B1(new_n782), .B2(G137), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n776), .A2(new_n202), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n250), .B1(new_n773), .B2(new_n212), .C1(new_n768), .C2(new_n761), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G150), .C2(new_n795), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n803), .B1(new_n1208), .B2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1202), .A2(new_n745), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1089), .A2(new_n973), .B1(new_n1201), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n953), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1220), .B2(new_n1109), .ZN(G381));
  NAND3_X1  g1021(.A1(new_n1004), .A2(new_n1071), .A3(new_n1006), .ZN(new_n1222));
  OR2_X1    g1022(.A1(G393), .A2(G396), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1222), .A2(G384), .A3(G381), .A4(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(G378), .A2(KEYINPUT121), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT121), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1115), .B2(new_n1136), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G375), .A2(new_n1229), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1225), .A2(new_n1230), .ZN(G407));
  NOR2_X1   g1031(.A1(new_n1224), .A2(new_n674), .ZN(new_n1232));
  OAI21_X1  g1032(.A(G213), .B1(new_n1232), .B2(new_n1230), .ZN(G409));
  NAND3_X1  g1033(.A1(new_n1171), .A2(G378), .A3(new_n1199), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1090), .B1(new_n1105), .B2(new_n1100), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n953), .B1(new_n1235), .B2(new_n1108), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n973), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1168), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1196), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1226), .A2(new_n1228), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G213), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(G343), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT60), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1090), .B(new_n696), .C1(new_n1219), .C2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT60), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1218), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT122), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n852), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1249), .B2(new_n852), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1249), .A2(new_n852), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1243), .A2(G2897), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1249), .A2(new_n852), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT122), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1249), .A2(new_n1250), .A3(new_n852), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1254), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1255), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT61), .B1(new_n1245), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1243), .B1(new_n1234), .B2(new_n1240), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1261), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1265), .A2(KEYINPUT62), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT62), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1264), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(new_n810), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1003), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1222), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1070), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1047), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1002), .A3(new_n974), .A4(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1273), .A3(new_n1272), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1274), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1264), .B(KEYINPUT125), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1271), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT63), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1256), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1286));
  AND4_X1   g1086(.A1(new_n1254), .A2(new_n1259), .A3(new_n1260), .A4(new_n1256), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT124), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1257), .A2(new_n1262), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1265), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1285), .A2(new_n1280), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT123), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT123), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1283), .A2(new_n1295), .A3(new_n1284), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1292), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1282), .A2(new_n1299), .ZN(G405));
  INV_X1    g1100(.A(new_n1234), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1229), .B1(new_n1199), .B2(new_n1171), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT126), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1301), .A2(new_n1302), .A3(KEYINPUT126), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n1261), .ZN(new_n1305));
  OAI211_X1 g1105(.A(KEYINPUT126), .B(new_n1266), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1305), .A2(new_n1306), .B1(KEYINPUT127), .B2(new_n1280), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1280), .B(KEYINPUT127), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(G402));
endmodule


