//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  NAND2_X1  g0011(.A1(new_n206), .A2(G50), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  NAND4_X1  g0013(.A1(new_n213), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT66), .B(G77), .Z(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n218), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n214), .B(new_n221), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n216), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n216), .A2(G33), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n250), .B1(new_n251), .B2(new_n253), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n215), .B2(G20), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G50), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(KEYINPUT70), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n264), .A2(KEYINPUT70), .A3(new_n268), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT9), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n270), .B2(new_n271), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n280), .A2(G223), .B1(new_n223), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(G222), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n279), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n262), .B1(G33), .B2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n292), .A3(G274), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n286), .A2(new_n290), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(G226), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n287), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G200), .ZN(new_n298));
  INV_X1    g0098(.A(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G190), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n273), .A2(new_n275), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n298), .A2(KEYINPUT71), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n303), .A2(KEYINPUT10), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n298), .A2(KEYINPUT71), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n273), .A2(new_n306), .A3(new_n275), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n269), .B1(new_n310), .B2(new_n297), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n299), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n265), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n203), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT12), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n203), .A2(G20), .ZN(new_n320));
  INV_X1    g0120(.A(G77), .ZN(new_n321));
  INV_X1    g0121(.A(G50), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n320), .B1(new_n259), .B2(new_n321), .C1(new_n322), .C2(new_n253), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(KEYINPUT11), .A3(new_n263), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n261), .A2(new_n262), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G1), .B2(new_n216), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n319), .B(new_n324), .C1(new_n203), .C2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT11), .B1(new_n323), .B2(new_n263), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n294), .B1(G238), .B2(new_n295), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  INV_X1    g0131(.A(G226), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n284), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G232), .B2(new_n280), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n334), .B2(new_n292), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT13), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(G169), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n335), .B(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G179), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n337), .B1(new_n336), .B2(G169), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n329), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT72), .B1(new_n336), .B2(new_n304), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT72), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n340), .A2(new_n346), .A3(G190), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n329), .B1(new_n336), .B2(G200), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n222), .A2(new_n216), .B1(new_n351), .B2(new_n259), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n254), .A2(new_n253), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n263), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n267), .A2(G77), .B1(new_n222), .B2(new_n317), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n295), .A2(G244), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n293), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n280), .A2(G238), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n283), .A2(G232), .A3(new_n279), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n278), .A2(G107), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT69), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n292), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT69), .A4(new_n361), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n358), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n356), .B1(new_n366), .B2(G190), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(new_n366), .ZN(new_n369));
  INV_X1    g0169(.A(new_n366), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(G179), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n356), .B1(new_n366), .B2(G169), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n344), .A2(new_n350), .A3(new_n369), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n253), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G58), .A2(G68), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n204), .A2(new_n205), .A3(new_n379), .ZN(new_n380));
  AOI211_X1 g0180(.A(new_n376), .B(new_n378), .C1(new_n380), .C2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n252), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n216), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n384), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n387), .A2(KEYINPUT73), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n390), .A3(new_n386), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n381), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n203), .B1(new_n387), .B2(new_n388), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n380), .A2(G20), .ZN(new_n395));
  INV_X1    g0195(.A(new_n378), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n376), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(new_n263), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n258), .A2(new_n267), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n317), .B1(new_n255), .B2(new_n257), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n326), .A2(new_n257), .A3(new_n255), .ZN(new_n404));
  INV_X1    g0204(.A(new_n258), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(KEYINPUT74), .C1(new_n405), .C2(new_n317), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G223), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n279), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n332), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n276), .C2(new_n277), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n292), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI211_X1 g0216(.A(KEYINPUT75), .B(new_n292), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n292), .A2(G232), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n293), .A2(new_n419), .A3(new_n312), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n293), .A2(new_n419), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n310), .B1(new_n414), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT76), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G223), .A2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n332), .B2(G1698), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n283), .B1(G33), .B2(G87), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT75), .B1(new_n429), .B2(new_n292), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n414), .A2(new_n415), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n426), .B(new_n423), .C1(new_n432), .C2(new_n420), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n408), .A2(new_n425), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n408), .A2(new_n425), .A3(KEYINPUT18), .A4(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n422), .A2(G190), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n431), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n368), .B1(new_n414), .B2(new_n422), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n399), .A2(new_n442), .A3(new_n407), .ZN(new_n443));
  XOR2_X1   g0243(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n399), .A2(new_n442), .A3(new_n407), .A4(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n446), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n438), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n316), .A2(new_n375), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G257), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n454));
  OAI211_X1 g0254(.A(G250), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G294), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n286), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n289), .A2(G1), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  NAND2_X1  g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n286), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G264), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT83), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n462), .A2(G274), .A3(new_n292), .A4(new_n459), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT83), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n458), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(G179), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n467), .ZN(new_n471));
  OAI21_X1  g0271(.A(G169), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n216), .B(G87), .C1(new_n276), .C2(new_n277), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT22), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT22), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n283), .A2(new_n476), .A3(new_n216), .A4(G87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G116), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G20), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n216), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n209), .A2(KEYINPUT23), .A3(G20), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n478), .A2(new_n479), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n479), .B1(new_n478), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n263), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n215), .A2(G33), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n325), .A2(new_n265), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G107), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT25), .ZN(new_n494));
  AOI211_X1 g0294(.A(G107), .B(new_n265), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n488), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n473), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n368), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n458), .A2(new_n464), .A3(new_n304), .A4(new_n467), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G274), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n286), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n215), .A2(G45), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n460), .B2(new_n461), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n463), .A2(G270), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G264), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n511));
  OAI211_X1 g0311(.A(G257), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n512));
  INV_X1    g0312(.A(G303), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(new_n283), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n286), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n310), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n317), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n325), .A2(G116), .A3(new_n265), .A4(new_n489), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n261), .A2(new_n262), .B1(G20), .B2(new_n517), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n216), .C1(G33), .C2(new_n208), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n520), .A2(KEYINPUT20), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT20), .B1(new_n520), .B2(new_n522), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n518), .B(new_n519), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n516), .A2(KEYINPUT21), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT21), .B1(new_n516), .B2(new_n525), .ZN(new_n527));
  AND4_X1   g0327(.A1(G179), .A2(new_n525), .A3(new_n515), .A4(new_n510), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n510), .A2(new_n515), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n525), .B1(new_n530), .B2(G200), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n510), .A2(new_n515), .A3(G190), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n265), .A2(G97), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n491), .B2(G97), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n216), .A2(new_n252), .A3(G77), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT79), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT6), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT79), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n209), .A2(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n210), .A2(new_n540), .A3(new_n542), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(G20), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n387), .A2(new_n388), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n538), .B(new_n548), .C1(new_n549), .C2(new_n209), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n537), .B1(new_n550), .B2(new_n263), .ZN(new_n551));
  INV_X1    g0351(.A(new_n461), .ZN(new_n552));
  NOR2_X1   g0352(.A1(KEYINPUT5), .A2(G41), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n459), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(G257), .A3(new_n292), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n467), .ZN(new_n556));
  OAI211_X1 g0356(.A(G244), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n557));
  NOR2_X1   g0357(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n558), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n283), .A2(G244), .A3(new_n279), .A4(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n559), .A2(new_n561), .A3(new_n521), .A4(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n563), .B2(new_n286), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(KEYINPUT81), .B(new_n556), .C1(new_n563), .C2(new_n286), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n551), .B(new_n565), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n216), .B1(new_n331), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(G87), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n208), .A3(new_n209), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n216), .B(G68), .C1(new_n276), .C2(new_n277), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n570), .B1(new_n259), .B2(new_n208), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n263), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n351), .A2(new_n317), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n351), .C2(new_n490), .ZN(new_n580));
  INV_X1    g0380(.A(G250), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n289), .B2(G1), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n215), .A2(new_n506), .A3(G45), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n292), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G238), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n586));
  OAI211_X1 g0386(.A(G244), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n480), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n588), .B2(new_n286), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(G169), .ZN(new_n590));
  AOI211_X1 g0390(.A(G179), .B(new_n585), .C1(new_n588), .C2(new_n286), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n286), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n368), .B1(new_n593), .B2(new_n584), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n325), .A2(G87), .A3(new_n265), .A4(new_n489), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n578), .A2(new_n579), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n589), .A2(G190), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n580), .A2(new_n592), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n563), .A2(new_n286), .ZN(new_n600));
  INV_X1    g0400(.A(new_n556), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n310), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n548), .A2(new_n538), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n209), .B1(new_n387), .B2(new_n388), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n263), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n536), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n564), .A2(new_n312), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n603), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n569), .A2(new_n599), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n505), .A2(new_n534), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n453), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g0412(.A(new_n612), .B(KEYINPUT84), .Z(G372));
  AOI22_X1  g0413(.A1(new_n602), .A2(new_n310), .B1(new_n606), .B2(new_n536), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n597), .A2(new_n598), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n589), .A2(new_n312), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n580), .B(new_n616), .C1(G169), .C2(new_n589), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n614), .A2(new_n615), .A3(new_n608), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT85), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n609), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n621), .A2(new_n599), .A3(new_n622), .A4(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n619), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n499), .A2(new_n529), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n502), .A2(new_n503), .ZN(new_n627));
  INV_X1    g0427(.A(new_n498), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n610), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n630), .A3(new_n617), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n453), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n421), .A2(new_n424), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n408), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(new_n435), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n342), .A2(new_n343), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(new_n329), .B1(new_n350), .B2(new_n373), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n450), .A2(new_n451), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n314), .B1(new_n639), .B2(new_n309), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n632), .A2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(G330), .ZN(new_n642));
  XOR2_X1   g0442(.A(new_n534), .B(KEYINPUT86), .Z(new_n643));
  NAND3_X1  g0443(.A1(new_n215), .A2(new_n216), .A3(G13), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n525), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n529), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT87), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT87), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n642), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n498), .A2(new_n649), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n505), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT88), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT88), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n505), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n649), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n499), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n529), .A2(new_n649), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n659), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n500), .A2(new_n663), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT89), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n671), .A3(new_n668), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n665), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n219), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n573), .A2(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n213), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n677), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  INV_X1    g0482(.A(new_n617), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n569), .A2(new_n599), .A3(new_n609), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n504), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n685), .B2(new_n626), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n649), .B1(new_n686), .B2(new_n625), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n618), .B(new_n619), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n649), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n611), .A2(new_n663), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n466), .A2(new_n469), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n530), .A2(new_n312), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n564), .A4(new_n589), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI211_X1 g0498(.A(G179), .B(new_n589), .C1(new_n515), .C2(new_n510), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n501), .A3(new_n602), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n649), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n693), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n692), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n682), .B1(new_n710), .B2(G1), .ZN(G364));
  INV_X1    g0511(.A(new_n656), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n216), .A2(G13), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n215), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n676), .A2(KEYINPUT90), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT90), .B1(new_n676), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n654), .A2(new_n642), .A3(new_n655), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n712), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n262), .B1(G20), .B2(new_n310), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n248), .A2(G45), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n675), .A2(new_n283), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(new_n680), .C2(G45), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n675), .A2(new_n278), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(G355), .B1(new_n517), .B2(new_n675), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n727), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n718), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n216), .A2(new_n312), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G190), .A3(new_n368), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n283), .B1(new_n736), .B2(new_n202), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n216), .A2(G179), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n304), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n209), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n735), .A2(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n304), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n740), .B1(G50), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n377), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n304), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n216), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n743), .B1(KEYINPUT32), .B2(new_n747), .C1(new_n208), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n735), .A2(new_n744), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n737), .B(new_n750), .C1(new_n223), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n741), .A2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n738), .A2(G190), .A3(G200), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n203), .B1(new_n756), .B2(new_n572), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(KEYINPUT32), .B2(new_n747), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  INV_X1    g0559(.A(G329), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n739), .A2(new_n759), .B1(new_n745), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT92), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n755), .A2(new_n763), .B1(new_n764), .B2(new_n749), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n742), .A2(G326), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n513), .B2(new_n756), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n278), .B1(new_n751), .B2(new_n768), .C1(new_n769), .C2(new_n736), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n765), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n753), .A2(new_n758), .B1(new_n762), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n725), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n734), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n653), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n733), .B(new_n774), .C1(new_n775), .C2(new_n724), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n721), .A2(new_n776), .ZN(G396));
  NOR2_X1   g0577(.A1(new_n725), .A2(new_n722), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n734), .B1(G77), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n754), .A2(G283), .B1(new_n752), .B2(G116), .ZN(new_n781));
  INV_X1    g0581(.A(new_n742), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n513), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n739), .A2(new_n572), .B1(new_n745), .B2(new_n768), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT94), .Z(new_n786));
  OAI221_X1 g0586(.A(new_n278), .B1(new_n736), .B2(new_n764), .C1(new_n208), .C2(new_n749), .ZN(new_n787));
  INV_X1    g0587(.A(new_n756), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n787), .B1(G107), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n784), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n736), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G143), .B1(new_n752), .B2(G159), .ZN(new_n792));
  INV_X1    g0592(.A(G137), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n792), .B1(new_n782), .B2(new_n793), .C1(new_n251), .C2(new_n755), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT34), .Z(new_n795));
  OAI22_X1  g0595(.A1(new_n322), .A2(new_n756), .B1(new_n739), .B2(new_n203), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  INV_X1    g0597(.A(new_n745), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n278), .B1(new_n798), .B2(G132), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n799), .C1(new_n202), .C2(new_n749), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n790), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n780), .B1(new_n801), .B2(new_n725), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n371), .A2(new_n372), .A3(new_n649), .ZN(new_n803));
  INV_X1    g0603(.A(new_n356), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n369), .B1(new_n804), .B2(new_n663), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(new_n805), .B2(new_n374), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n802), .B1(new_n806), .B2(new_n723), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n631), .A2(new_n663), .A3(new_n806), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT97), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n687), .A2(KEYINPUT97), .A3(new_n806), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n806), .B(KEYINPUT96), .ZN(new_n813));
  INV_X1    g0613(.A(new_n687), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n708), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n718), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(new_n708), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n807), .B1(new_n818), .B2(new_n819), .ZN(G384));
  NAND3_X1  g0620(.A1(new_n213), .A2(new_n223), .A3(new_n379), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n322), .A2(G68), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n215), .B(G13), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n262), .A2(new_n216), .A3(new_n517), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n545), .A2(new_n547), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT35), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n344), .A2(new_n350), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(new_n329), .A3(new_n649), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n329), .A2(new_n649), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n344), .A2(new_n350), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(new_n707), .A3(new_n806), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n434), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n647), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n408), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n443), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n404), .B1(new_n405), .B2(new_n317), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n393), .A2(new_n263), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n387), .A2(KEYINPUT73), .A3(new_n388), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(G68), .A3(new_n391), .ZN(new_n846));
  INV_X1    g0646(.A(new_n397), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT16), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n843), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT99), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n843), .B(KEYINPUT99), .C1(new_n844), .C2(new_n848), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n633), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n839), .A3(new_n852), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n854), .A3(new_n443), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n842), .B1(new_n855), .B2(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n325), .B1(new_n846), .B2(new_n381), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(new_n398), .B1(new_n403), .B2(new_n406), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n444), .B1(new_n859), .B2(new_n442), .ZN(new_n860));
  AND4_X1   g0660(.A1(new_n442), .A2(new_n399), .A3(new_n407), .A4(new_n448), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT78), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n862), .A2(new_n863), .B1(new_n436), .B2(new_n437), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT100), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n864), .A2(new_n865), .A3(new_n854), .ZN(new_n866));
  INV_X1    g0666(.A(new_n854), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT100), .B1(new_n452), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n857), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n634), .A2(new_n840), .A3(new_n443), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n842), .B1(KEYINPUT37), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n446), .A2(new_n449), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n840), .B1(new_n635), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n836), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n836), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n865), .B1(new_n864), .B2(new_n854), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n452), .A2(KEYINPUT100), .A3(new_n867), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n882), .B2(new_n857), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n870), .B(new_n856), .C1(new_n880), .C2(new_n881), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT101), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT101), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n857), .B1(new_n866), .B2(new_n868), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n870), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(new_n869), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n879), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n878), .B1(new_n890), .B2(new_n877), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n453), .A2(new_n707), .ZN(new_n893));
  OAI21_X1  g0693(.A(G330), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n635), .A2(new_n839), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT98), .ZN(new_n897));
  INV_X1    g0697(.A(new_n803), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n812), .B2(new_n898), .ZN(new_n899));
  AOI211_X1 g0699(.A(KEYINPUT98), .B(new_n803), .C1(new_n810), .C2(new_n811), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n835), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n885), .A2(new_n889), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n636), .A2(new_n329), .A3(new_n663), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n888), .B2(new_n869), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT102), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n906), .A2(new_n907), .B1(new_n905), .B2(new_n876), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT39), .B1(new_n883), .B2(new_n884), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT102), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n904), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n453), .A2(new_n688), .A3(new_n691), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n640), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n895), .A2(new_n915), .B1(new_n215), .B2(new_n713), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n895), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n830), .B1(new_n916), .B2(new_n917), .ZN(G367));
  OAI211_X1 g0718(.A(new_n569), .B(new_n609), .C1(new_n551), .C2(new_n663), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n621), .A2(new_n649), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT104), .B1(new_n665), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n596), .A2(new_n649), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n599), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n617), .B2(new_n925), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n667), .A2(new_n922), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n621), .B1(new_n500), .B2(new_n569), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n649), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT103), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(KEYINPUT103), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n928), .A2(new_n929), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n930), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n929), .B(new_n928), .C1(new_n941), .C2(new_n934), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n924), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n942), .A2(new_n940), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT104), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n656), .A2(new_n945), .A3(new_n664), .A4(new_n921), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n923), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n943), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n676), .B(KEYINPUT41), .Z(new_n949));
  NAND3_X1  g0749(.A1(new_n670), .A2(new_n672), .A3(new_n922), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT44), .Z(new_n951));
  AOI21_X1  g0751(.A(new_n922), .B1(new_n670), .B2(new_n672), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n665), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n665), .A3(new_n953), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n667), .B1(new_n664), .B2(new_n666), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n656), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n656), .A2(new_n958), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n709), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n956), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n949), .B1(new_n962), .B2(new_n710), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n948), .B1(new_n963), .B2(new_n715), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n928), .A2(new_n724), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n729), .A2(new_n241), .ZN(new_n966));
  INV_X1    g0766(.A(new_n351), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n727), .B1(new_n675), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n718), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n791), .A2(G150), .B1(new_n798), .B2(G137), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n970), .B(new_n283), .C1(new_n322), .C2(new_n751), .ZN(new_n971));
  INV_X1    g0771(.A(new_n749), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n972), .A2(G68), .B1(new_n788), .B2(G58), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n377), .B2(new_n755), .ZN(new_n974));
  INV_X1    g0774(.A(G143), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n782), .A2(new_n975), .B1(new_n222), .B2(new_n739), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT106), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n756), .A2(new_n517), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(KEYINPUT46), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT105), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n278), .B1(new_n751), .B2(new_n759), .ZN(new_n982));
  INV_X1    g0782(.A(G317), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n736), .A2(new_n513), .B1(new_n745), .B2(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(KEYINPUT46), .C2(new_n979), .ZN(new_n985));
  INV_X1    g0785(.A(new_n739), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n754), .A2(G294), .B1(new_n986), .B2(G97), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G107), .A2(new_n972), .B1(new_n742), .B2(G311), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n981), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n978), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT47), .Z(new_n991));
  OAI211_X1 g0791(.A(new_n965), .B(new_n969), .C1(new_n991), .C2(new_n773), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n964), .A2(new_n992), .ZN(G387));
  INV_X1    g0793(.A(new_n678), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n731), .A2(new_n994), .B1(new_n209), .B2(new_n675), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n678), .A2(KEYINPUT107), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n678), .A2(KEYINPUT107), .ZN(new_n997));
  AOI21_X1  g0797(.A(G45), .B1(G68), .B2(G77), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT108), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n254), .A2(G50), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT50), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n729), .B1(new_n238), .B2(new_n289), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n995), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n718), .B1(new_n1005), .B2(new_n726), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n283), .B1(new_n798), .B2(G326), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n749), .A2(new_n759), .B1(new_n756), .B2(new_n764), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n791), .A2(G317), .B1(new_n752), .B2(G303), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n782), .B2(new_n769), .C1(new_n768), .C2(new_n755), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1007), .B1(new_n517), .B2(new_n739), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n278), .B1(new_n798), .B2(G150), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n208), .B2(new_n739), .C1(new_n222), .C2(new_n756), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT109), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n749), .A2(new_n351), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n791), .A2(G50), .B1(new_n752), .B2(G68), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n377), .B2(new_n782), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(new_n405), .C2(new_n754), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1016), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1006), .B1(new_n1024), .B2(new_n773), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n664), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(new_n724), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n959), .A2(new_n960), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(new_n715), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n961), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n676), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1028), .A2(new_n710), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G393));
  INV_X1    g0833(.A(new_n957), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n665), .B1(new_n951), .B2(new_n953), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(new_n962), .A3(new_n676), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n922), .A2(new_n724), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n726), .B1(new_n208), .B2(new_n219), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n729), .B2(new_n245), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT110), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G150), .A2(new_n742), .B1(new_n791), .B2(G159), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT51), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n755), .A2(new_n322), .B1(new_n321), .B2(new_n749), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n283), .B1(new_n745), .B2(new_n975), .C1(new_n254), .C2(new_n751), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n203), .A2(new_n756), .B1(new_n739), .B2(new_n572), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n283), .B(new_n740), .C1(G294), .C2(new_n752), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n756), .A2(new_n759), .B1(new_n745), .B2(new_n769), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT111), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(KEYINPUT111), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G116), .A2(new_n972), .B1(new_n754), .B2(G303), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G317), .A2(new_n742), .B1(new_n791), .B2(G311), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT52), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1044), .A2(new_n1048), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n718), .B(new_n1042), .C1(new_n1057), .C2(new_n725), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT112), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1038), .A2(new_n715), .B1(new_n1039), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1037), .A2(new_n1060), .ZN(G390));
  INV_X1    g0861(.A(new_n835), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n707), .A2(G330), .A3(new_n806), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n805), .A2(new_n374), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n690), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n835), .B1(new_n1066), .B2(new_n803), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n869), .A2(new_n875), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n904), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n901), .A2(new_n904), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n907), .B(KEYINPUT39), .C1(new_n883), .C2(new_n884), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n869), .A2(new_n905), .A3(new_n875), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n888), .A2(new_n869), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n907), .B1(new_n1075), .B2(KEYINPUT39), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1064), .B(new_n1070), .C1(new_n1071), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1064), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT97), .B1(new_n687), .B2(new_n806), .ZN(new_n1080));
  AND4_X1   g0880(.A1(KEYINPUT97), .A2(new_n631), .A3(new_n663), .A4(new_n806), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n898), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT98), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n812), .A2(new_n897), .A3(new_n898), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1062), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n904), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n910), .B(new_n908), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1079), .B1(new_n1087), .B2(new_n1069), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1078), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n453), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n913), .B(new_n640), .C1(new_n1090), .C2(new_n708), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1064), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1066), .A2(new_n803), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1062), .B1(new_n708), .B2(new_n813), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1079), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1091), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n677), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1086), .B1(new_n1092), .B2(new_n835), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n910), .A2(new_n1073), .A3(new_n1072), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1069), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1064), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1087), .A2(new_n1079), .A3(new_n1069), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1091), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT113), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT113), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1110), .B(new_n1098), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1099), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n718), .B1(new_n258), .B2(new_n778), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n755), .A2(new_n793), .B1(new_n751), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G159), .B2(new_n972), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT114), .Z(new_n1117));
  AOI21_X1  g0917(.A(new_n278), .B1(new_n798), .B2(G125), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n322), .B2(new_n739), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT115), .Z(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n788), .B2(G150), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n788), .A2(new_n1121), .A3(G150), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n791), .A2(G132), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1124), .C1(new_n782), .C2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1120), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n782), .A2(new_n759), .B1(new_n321), .B2(new_n749), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n278), .B1(new_n745), .B2(new_n764), .C1(new_n736), .C2(new_n517), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n203), .A2(new_n739), .B1(new_n756), .B2(new_n572), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n754), .A2(G107), .B1(new_n752), .B2(G97), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT117), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1117), .A2(new_n1127), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1113), .B1(new_n773), .B2(new_n1134), .C1(new_n1101), .C2(new_n723), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1105), .B2(new_n714), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1112), .A2(new_n1137), .ZN(G378));
  OAI21_X1  g0938(.A(KEYINPUT120), .B1(new_n903), .B2(new_n911), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n272), .A2(new_n647), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n316), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1140), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n309), .B2(new_n315), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OR3_X1    g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n891), .B2(G330), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n879), .A2(KEYINPUT40), .A3(new_n1068), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT101), .B1(new_n883), .B2(new_n884), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n888), .A2(new_n886), .A3(new_n869), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n836), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(G330), .B(new_n1150), .C1(new_n1153), .C2(KEYINPUT40), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1139), .B1(new_n1149), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n891), .A2(G330), .A3(new_n1148), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1086), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1085), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1162), .A3(new_n896), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1158), .A2(KEYINPUT120), .A3(new_n1159), .A4(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1157), .A2(new_n715), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n734), .B1(G50), .B2(new_n779), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n755), .A2(new_n208), .B1(new_n739), .B2(new_n202), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G116), .B2(new_n742), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n278), .A2(new_n288), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G283), .B2(new_n798), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n791), .A2(G107), .B1(new_n752), .B2(new_n967), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n972), .A2(G68), .B1(new_n223), .B2(new_n788), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1169), .B(new_n322), .C1(G33), .C2(G41), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n754), .A2(G132), .B1(new_n752), .B2(G137), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT118), .Z(new_n1179));
  OAI22_X1  g0979(.A1(new_n736), .A2(new_n1125), .B1(new_n756), .B2(new_n1114), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT119), .Z(new_n1181));
  AOI22_X1  g0981(.A1(G150), .A2(new_n972), .B1(new_n742), .B2(G125), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n986), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1177), .B1(new_n1174), .B2(new_n1173), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1166), .B1(new_n1189), .B2(new_n725), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1148), .B2(new_n723), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT121), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT121), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1165), .A2(new_n1194), .A3(new_n1191), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1091), .B1(new_n1089), .B2(new_n1106), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1157), .A2(new_n1164), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1163), .B1(new_n1149), .B2(new_n1156), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n912), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1103), .A2(new_n1104), .A3(new_n1098), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1107), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n677), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1200), .A2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1196), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(G375));
  NAND2_X1  g1009(.A1(new_n1062), .A2(new_n722), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n734), .B1(G68), .B2(new_n779), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n755), .A2(new_n517), .B1(new_n782), .B2(new_n764), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G97), .B2(new_n788), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n736), .A2(new_n759), .B1(new_n751), .B2(new_n209), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n283), .B(new_n1214), .C1(G303), .C2(new_n798), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1020), .B1(G77), .B2(new_n986), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT123), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n736), .A2(new_n793), .B1(new_n745), .B2(new_n1125), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n278), .B(new_n1220), .C1(G150), .C2(new_n752), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n742), .A2(G132), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1114), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G50), .A2(new_n972), .B1(new_n754), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n788), .A2(G159), .B1(new_n986), .B2(G58), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1219), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1211), .B1(new_n1228), .B2(new_n725), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT124), .Z(new_n1230));
  AOI22_X1  g1030(.A1(new_n1106), .A2(new_n715), .B1(new_n1210), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1091), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT122), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1232), .B(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1098), .A2(new_n949), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1231), .B1(new_n1234), .B2(new_n1235), .ZN(G381));
  OR3_X1    g1036(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(G387), .A2(new_n1237), .A3(G390), .A4(G381), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT125), .ZN(new_n1239));
  INV_X1    g1039(.A(G378), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1208), .ZN(G407));
  INV_X1    g1041(.A(G213), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(G343), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1208), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G407), .A2(G213), .A3(new_n1244), .ZN(G409));
  NAND3_X1  g1045(.A1(new_n1196), .A2(new_n1207), .A3(G378), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1198), .A2(new_n949), .A3(new_n1199), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1191), .B1(new_n1248), .B2(new_n714), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1112), .B(new_n1137), .C1(new_n1247), .C2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1243), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1232), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n677), .B1(new_n1254), .B2(KEYINPUT60), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1234), .B2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(KEYINPUT126), .B(new_n807), .C1(new_n818), .C2(new_n819), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1257), .A2(new_n1231), .A3(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(G384), .B(KEYINPUT126), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1257), .B2(new_n1231), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1243), .A2(G2897), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G2897), .B(new_n1243), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n964), .A2(new_n992), .A3(G390), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(G396), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G390), .B1(new_n964), .B2(new_n992), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1269), .A2(new_n1274), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1243), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1262), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1279), .B2(new_n1262), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1267), .B(new_n1278), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1279), .A2(new_n1284), .A3(new_n1262), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1286), .B1(new_n1279), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1284), .B1(new_n1279), .B2(new_n1262), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1285), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1283), .B1(new_n1290), .B2(new_n1278), .ZN(G405));
  INV_X1    g1091(.A(new_n1262), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1276), .A2(new_n1277), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1292), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1208), .B(G378), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1208), .B(new_n1240), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1278), .A2(new_n1262), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(new_n1293), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1297), .A2(new_n1300), .ZN(G402));
endmodule


