

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n610), .A2(n515), .ZN(n611) );
  AND2_X1 U550 ( .A1(n684), .A2(n683), .ZN(n514) );
  AND2_X1 U551 ( .A1(n609), .A2(n608), .ZN(n515) );
  AND2_X1 U552 ( .A1(n614), .A2(G1996), .ZN(n595) );
  INV_X1 U553 ( .A(n954), .ZN(n688) );
  NOR2_X1 U554 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U555 ( .A1(G2105), .A2(n522), .ZN(n869) );
  NOR2_X1 U556 ( .A1(G651), .A2(n577), .ZN(n775) );
  NOR2_X1 U557 ( .A1(n527), .A2(n526), .ZN(n594) );
  BUF_X1 U558 ( .A(n594), .Z(G160) );
  NAND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  XOR2_X2 U560 ( .A(KEYINPUT66), .B(n516), .Z(n866) );
  NAND2_X1 U561 ( .A1(n866), .A2(G113), .ZN(n517) );
  XOR2_X1 U562 ( .A(KEYINPUT67), .B(n517), .Z(n520) );
  INV_X1 U563 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U564 ( .A1(G101), .A2(n869), .ZN(n518) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U566 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X1 U568 ( .A(KEYINPUT17), .B(n521), .Z(n871) );
  NAND2_X1 U569 ( .A1(G137), .A2(n871), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n522), .A2(G2105), .ZN(n523) );
  XNOR2_X1 U571 ( .A(n523), .B(KEYINPUT65), .ZN(n865) );
  NAND2_X1 U572 ( .A1(G125), .A2(n865), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n869), .A2(G102), .ZN(n530) );
  NAND2_X1 U575 ( .A1(G114), .A2(n866), .ZN(n528) );
  XOR2_X1 U576 ( .A(n528), .B(KEYINPUT87), .Z(n529) );
  NAND2_X1 U577 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U578 ( .A1(G138), .A2(n871), .ZN(n532) );
  NAND2_X1 U579 ( .A1(G126), .A2(n865), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n534), .A2(n533), .ZN(G164) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  INV_X1 U583 ( .A(G651), .ZN(n541) );
  NOR2_X1 U584 ( .A1(n577), .A2(n541), .ZN(n779) );
  NAND2_X1 U585 ( .A1(n779), .A2(G77), .ZN(n535) );
  XNOR2_X1 U586 ( .A(KEYINPUT69), .B(n535), .ZN(n538) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n778) );
  NAND2_X1 U588 ( .A1(n778), .A2(G90), .ZN(n536) );
  XOR2_X1 U589 ( .A(n536), .B(KEYINPUT68), .Z(n537) );
  NOR2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  XNOR2_X1 U592 ( .A(KEYINPUT70), .B(n540), .ZN(n546) );
  NOR2_X1 U593 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n542), .Z(n774) );
  NAND2_X1 U595 ( .A1(G64), .A2(n774), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G52), .A2(n775), .ZN(n543) );
  AND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(G301) );
  NAND2_X1 U599 ( .A1(n778), .A2(G89), .ZN(n547) );
  XNOR2_X1 U600 ( .A(n547), .B(KEYINPUT4), .ZN(n549) );
  NAND2_X1 U601 ( .A1(G76), .A2(n779), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n550), .B(KEYINPUT5), .ZN(n555) );
  NAND2_X1 U604 ( .A1(G63), .A2(n774), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G51), .A2(n775), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U609 ( .A(n556), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(G50), .A2(n775), .ZN(n563) );
  NAND2_X1 U612 ( .A1(G88), .A2(n778), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G62), .A2(n774), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n779), .A2(G75), .ZN(n559) );
  XOR2_X1 U616 ( .A(KEYINPUT82), .B(n559), .Z(n560) );
  NOR2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U619 ( .A(n564), .B(KEYINPUT83), .ZN(G166) );
  INV_X1 U620 ( .A(G166), .ZN(G303) );
  NAND2_X1 U621 ( .A1(G86), .A2(n778), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G61), .A2(n774), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n779), .A2(G73), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT2), .B(n567), .Z(n568) );
  NOR2_X1 U626 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U627 ( .A1(n775), .A2(G48), .ZN(n570) );
  NAND2_X1 U628 ( .A1(n571), .A2(n570), .ZN(G305) );
  NAND2_X1 U629 ( .A1(G651), .A2(G74), .ZN(n572) );
  XNOR2_X1 U630 ( .A(n572), .B(KEYINPUT80), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G49), .A2(n775), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U633 ( .A(KEYINPUT81), .B(n575), .Z(n576) );
  NOR2_X1 U634 ( .A1(n774), .A2(n576), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n577), .A2(G87), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U637 ( .A1(G85), .A2(n778), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G72), .A2(n779), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U640 ( .A1(G60), .A2(n774), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G47), .A2(n775), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n584) );
  OR2_X1 U643 ( .A1(n585), .A2(n584), .ZN(G290) );
  NAND2_X1 U644 ( .A1(G66), .A2(n774), .ZN(n592) );
  NAND2_X1 U645 ( .A1(G92), .A2(n778), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G79), .A2(n779), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U648 ( .A1(n775), .A2(G54), .ZN(n588) );
  XOR2_X1 U649 ( .A(KEYINPUT78), .B(n588), .Z(n589) );
  NOR2_X1 U650 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U651 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U652 ( .A(n593), .B(KEYINPUT15), .ZN(n970) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n698) );
  AND2_X1 U654 ( .A1(n594), .A2(G40), .ZN(n696) );
  AND2_X1 U655 ( .A1(n698), .A2(n696), .ZN(n614) );
  XOR2_X1 U656 ( .A(n595), .B(KEYINPUT26), .Z(n610) );
  XNOR2_X1 U657 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n601) );
  NAND2_X1 U658 ( .A1(n778), .A2(G81), .ZN(n596) );
  XNOR2_X1 U659 ( .A(n596), .B(KEYINPUT12), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G68), .A2(n779), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U662 ( .A(n599), .B(KEYINPUT13), .ZN(n600) );
  XNOR2_X1 U663 ( .A(n601), .B(n600), .ZN(n605) );
  NAND2_X1 U664 ( .A1(G56), .A2(n774), .ZN(n602) );
  XNOR2_X1 U665 ( .A(n602), .B(KEYINPUT14), .ZN(n603) );
  XNOR2_X1 U666 ( .A(KEYINPUT75), .B(n603), .ZN(n604) );
  NOR2_X1 U667 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U668 ( .A1(n775), .A2(G43), .ZN(n606) );
  NAND2_X2 U669 ( .A1(n607), .A2(n606), .ZN(n958) );
  INV_X1 U670 ( .A(n958), .ZN(n609) );
  NAND2_X1 U671 ( .A1(n698), .A2(n696), .ZN(n654) );
  NAND2_X1 U672 ( .A1(n654), .A2(G1341), .ZN(n608) );
  XNOR2_X1 U673 ( .A(n611), .B(KEYINPUT64), .ZN(n613) );
  NOR2_X1 U674 ( .A1(n970), .A2(n613), .ZN(n612) );
  XNOR2_X1 U675 ( .A(n612), .B(KEYINPUT93), .ZN(n620) );
  NAND2_X1 U676 ( .A1(n970), .A2(n613), .ZN(n618) );
  INV_X1 U677 ( .A(n654), .ZN(n638) );
  NOR2_X1 U678 ( .A1(n638), .A2(G1348), .ZN(n616) );
  NOR2_X1 U679 ( .A1(G2067), .A2(n654), .ZN(n615) );
  NOR2_X1 U680 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U681 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U682 ( .A1(n620), .A2(n619), .ZN(n631) );
  NAND2_X1 U683 ( .A1(G65), .A2(n774), .ZN(n622) );
  NAND2_X1 U684 ( .A1(G53), .A2(n775), .ZN(n621) );
  NAND2_X1 U685 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U686 ( .A1(G91), .A2(n778), .ZN(n624) );
  NAND2_X1 U687 ( .A1(G78), .A2(n779), .ZN(n623) );
  NAND2_X1 U688 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U689 ( .A1(n626), .A2(n625), .ZN(n959) );
  NAND2_X1 U690 ( .A1(n638), .A2(G2072), .ZN(n627) );
  XNOR2_X1 U691 ( .A(n627), .B(KEYINPUT27), .ZN(n629) );
  INV_X1 U692 ( .A(G1956), .ZN(n988) );
  NOR2_X1 U693 ( .A1(n988), .A2(n638), .ZN(n628) );
  NOR2_X1 U694 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U695 ( .A1(n959), .A2(n632), .ZN(n630) );
  NAND2_X1 U696 ( .A1(n631), .A2(n630), .ZN(n635) );
  NOR2_X1 U697 ( .A1(n959), .A2(n632), .ZN(n633) );
  XOR2_X1 U698 ( .A(n633), .B(KEYINPUT28), .Z(n634) );
  NAND2_X1 U699 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U700 ( .A(n636), .B(KEYINPUT29), .ZN(n642) );
  XOR2_X1 U701 ( .A(G2078), .B(KEYINPUT25), .Z(n637) );
  XNOR2_X1 U702 ( .A(KEYINPUT92), .B(n637), .ZN(n943) );
  NOR2_X1 U703 ( .A1(n654), .A2(n943), .ZN(n640) );
  NOR2_X1 U704 ( .A1(n638), .A2(G1961), .ZN(n639) );
  NOR2_X1 U705 ( .A1(n640), .A2(n639), .ZN(n643) );
  NOR2_X1 U706 ( .A1(G301), .A2(n643), .ZN(n641) );
  NOR2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n652) );
  AND2_X1 U708 ( .A1(G301), .A2(n643), .ZN(n648) );
  NAND2_X1 U709 ( .A1(G8), .A2(n654), .ZN(n686) );
  NOR2_X1 U710 ( .A1(G1966), .A2(n686), .ZN(n663) );
  NOR2_X1 U711 ( .A1(G2084), .A2(n654), .ZN(n664) );
  NOR2_X1 U712 ( .A1(n663), .A2(n664), .ZN(n644) );
  NAND2_X1 U713 ( .A1(G8), .A2(n644), .ZN(n645) );
  XNOR2_X1 U714 ( .A(KEYINPUT30), .B(n645), .ZN(n646) );
  NOR2_X1 U715 ( .A1(G168), .A2(n646), .ZN(n647) );
  NOR2_X1 U716 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U717 ( .A(KEYINPUT31), .B(n649), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT94), .B(n650), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n652), .A2(n651), .ZN(n662) );
  INV_X1 U720 ( .A(n662), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n653), .A2(G286), .ZN(n659) );
  NOR2_X1 U722 ( .A1(G1971), .A2(n686), .ZN(n656) );
  NOR2_X1 U723 ( .A1(G2090), .A2(n654), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n657), .A2(G303), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n660), .A2(G8), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n661), .B(KEYINPUT32), .ZN(n669) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U730 ( .A1(G8), .A2(n664), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT95), .B(n667), .Z(n668) );
  NAND2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n680) );
  NOR2_X1 U734 ( .A1(G2090), .A2(G303), .ZN(n670) );
  NAND2_X1 U735 ( .A1(G8), .A2(n670), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n680), .A2(n671), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT96), .ZN(n673) );
  AND2_X1 U738 ( .A1(n673), .A2(n686), .ZN(n694) );
  NOR2_X1 U739 ( .A1(G1981), .A2(G305), .ZN(n674) );
  XOR2_X1 U740 ( .A(n674), .B(KEYINPUT24), .Z(n675) );
  NOR2_X1 U741 ( .A1(n686), .A2(n675), .ZN(n676) );
  XNOR2_X1 U742 ( .A(KEYINPUT91), .B(n676), .ZN(n692) );
  NOR2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U744 ( .A1(G1971), .A2(G303), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n685), .A2(n677), .ZN(n963) );
  INV_X1 U746 ( .A(KEYINPUT33), .ZN(n678) );
  AND2_X1 U747 ( .A1(n963), .A2(n678), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n684) );
  INV_X1 U749 ( .A(n686), .ZN(n681) );
  NAND2_X1 U750 ( .A1(G1976), .A2(G288), .ZN(n962) );
  AND2_X1 U751 ( .A1(n681), .A2(n962), .ZN(n682) );
  OR2_X1 U752 ( .A1(KEYINPUT33), .A2(n682), .ZN(n683) );
  NAND2_X1 U753 ( .A1(n685), .A2(KEYINPUT33), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n689) );
  XOR2_X1 U755 ( .A(G1981), .B(G305), .Z(n954) );
  NAND2_X1 U756 ( .A1(n514), .A2(n690), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U759 ( .A(n695), .B(KEYINPUT97), .ZN(n731) );
  XNOR2_X1 U760 ( .A(G1986), .B(G290), .ZN(n968) );
  INV_X1 U761 ( .A(n696), .ZN(n697) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n744) );
  NAND2_X1 U763 ( .A1(n968), .A2(n744), .ZN(n729) );
  NAND2_X1 U764 ( .A1(G95), .A2(n869), .ZN(n700) );
  NAND2_X1 U765 ( .A1(G131), .A2(n871), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U767 ( .A1(n865), .A2(G119), .ZN(n702) );
  NAND2_X1 U768 ( .A1(G107), .A2(n866), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n877) );
  NAND2_X1 U771 ( .A1(G1991), .A2(n877), .ZN(n705) );
  XNOR2_X1 U772 ( .A(n705), .B(KEYINPUT89), .ZN(n714) );
  NAND2_X1 U773 ( .A1(G141), .A2(n871), .ZN(n707) );
  NAND2_X1 U774 ( .A1(G129), .A2(n865), .ZN(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U776 ( .A1(n869), .A2(G105), .ZN(n708) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n708), .Z(n709) );
  NOR2_X1 U778 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U779 ( .A1(G117), .A2(n866), .ZN(n711) );
  NAND2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n882) );
  AND2_X1 U781 ( .A1(G1996), .A2(n882), .ZN(n713) );
  NOR2_X1 U782 ( .A1(n714), .A2(n713), .ZN(n909) );
  INV_X1 U783 ( .A(n744), .ZN(n715) );
  NOR2_X1 U784 ( .A1(n909), .A2(n715), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n735), .B(KEYINPUT90), .ZN(n727) );
  NAND2_X1 U786 ( .A1(G104), .A2(n869), .ZN(n717) );
  NAND2_X1 U787 ( .A1(G140), .A2(n871), .ZN(n716) );
  NAND2_X1 U788 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U789 ( .A(KEYINPUT34), .B(n718), .ZN(n723) );
  NAND2_X1 U790 ( .A1(n865), .A2(G128), .ZN(n720) );
  NAND2_X1 U791 ( .A1(G116), .A2(n866), .ZN(n719) );
  NAND2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U793 ( .A(KEYINPUT35), .B(n721), .Z(n722) );
  NOR2_X1 U794 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U795 ( .A(KEYINPUT36), .B(n724), .ZN(n864) );
  XNOR2_X1 U796 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  NOR2_X1 U797 ( .A1(n864), .A2(n742), .ZN(n925) );
  NAND2_X1 U798 ( .A1(n925), .A2(n744), .ZN(n725) );
  XNOR2_X1 U799 ( .A(n725), .B(KEYINPUT88), .ZN(n740) );
  INV_X1 U800 ( .A(n740), .ZN(n726) );
  NOR2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n728) );
  AND2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n747) );
  XOR2_X1 U804 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n732) );
  XNOR2_X1 U805 ( .A(KEYINPUT39), .B(n732), .ZN(n739) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n882), .ZN(n916) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n733) );
  NOR2_X1 U808 ( .A1(G1991), .A2(n877), .ZN(n907) );
  NOR2_X1 U809 ( .A1(n733), .A2(n907), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U811 ( .A(n736), .B(KEYINPUT98), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n916), .A2(n737), .ZN(n738) );
  XNOR2_X1 U813 ( .A(n739), .B(n738), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n864), .A2(n742), .ZN(n922) );
  NAND2_X1 U816 ( .A1(n743), .A2(n922), .ZN(n745) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U819 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U820 ( .A1(G99), .A2(n869), .ZN(n750) );
  NAND2_X1 U821 ( .A1(G135), .A2(n871), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n753) );
  NAND2_X1 U823 ( .A1(n865), .A2(G123), .ZN(n751) );
  XOR2_X1 U824 ( .A(KEYINPUT18), .B(n751), .Z(n752) );
  NOR2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U826 ( .A1(G111), .A2(n866), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n904) );
  XNOR2_X1 U828 ( .A(G2096), .B(n904), .ZN(n756) );
  OR2_X1 U829 ( .A1(G2100), .A2(n756), .ZN(G156) );
  INV_X1 U830 ( .A(G57), .ZN(G237) );
  INV_X1 U831 ( .A(G132), .ZN(G219) );
  NAND2_X1 U832 ( .A1(G94), .A2(G452), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n757), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n758) );
  XNOR2_X1 U835 ( .A(n758), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U836 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n760) );
  XNOR2_X1 U837 ( .A(G223), .B(KEYINPUT73), .ZN(n819) );
  NAND2_X1 U838 ( .A1(G567), .A2(n819), .ZN(n759) );
  XNOR2_X1 U839 ( .A(n760), .B(n759), .ZN(G234) );
  INV_X1 U840 ( .A(G860), .ZN(n773) );
  OR2_X1 U841 ( .A1(n958), .A2(n773), .ZN(G153) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n762) );
  OR2_X1 U843 ( .A1(n970), .A2(G868), .ZN(n761) );
  NAND2_X1 U844 ( .A1(n762), .A2(n761), .ZN(G284) );
  INV_X1 U845 ( .A(n959), .ZN(G299) );
  INV_X1 U846 ( .A(G868), .ZN(n763) );
  NOR2_X1 U847 ( .A1(G286), .A2(n763), .ZN(n765) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n764) );
  NOR2_X1 U849 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n773), .A2(G559), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n766), .A2(n970), .ZN(n767) );
  XNOR2_X1 U852 ( .A(n767), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U853 ( .A1(G868), .A2(n958), .ZN(n768) );
  XOR2_X1 U854 ( .A(KEYINPUT79), .B(n768), .Z(n771) );
  NAND2_X1 U855 ( .A1(G868), .A2(n970), .ZN(n769) );
  NOR2_X1 U856 ( .A1(G559), .A2(n769), .ZN(n770) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(G282) );
  NAND2_X1 U858 ( .A1(G559), .A2(n970), .ZN(n772) );
  XOR2_X1 U859 ( .A(n958), .B(n772), .Z(n790) );
  NAND2_X1 U860 ( .A1(n773), .A2(n790), .ZN(n784) );
  NAND2_X1 U861 ( .A1(G67), .A2(n774), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G55), .A2(n775), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n783) );
  NAND2_X1 U864 ( .A1(G93), .A2(n778), .ZN(n781) );
  NAND2_X1 U865 ( .A1(G80), .A2(n779), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n792) );
  XOR2_X1 U868 ( .A(n784), .B(n792), .Z(G145) );
  XNOR2_X1 U869 ( .A(KEYINPUT19), .B(G290), .ZN(n785) );
  XNOR2_X1 U870 ( .A(n785), .B(G305), .ZN(n786) );
  XOR2_X1 U871 ( .A(n786), .B(n792), .Z(n788) );
  XNOR2_X1 U872 ( .A(G166), .B(n959), .ZN(n787) );
  XNOR2_X1 U873 ( .A(n788), .B(n787), .ZN(n789) );
  XNOR2_X1 U874 ( .A(n789), .B(G288), .ZN(n893) );
  XNOR2_X1 U875 ( .A(n790), .B(n893), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n791), .A2(G868), .ZN(n794) );
  OR2_X1 U877 ( .A1(G868), .A2(n792), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(G295) );
  NAND2_X1 U879 ( .A1(G2084), .A2(G2078), .ZN(n795) );
  XOR2_X1 U880 ( .A(KEYINPUT20), .B(n795), .Z(n796) );
  NAND2_X1 U881 ( .A1(G2090), .A2(n796), .ZN(n797) );
  XNOR2_X1 U882 ( .A(KEYINPUT21), .B(n797), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n798), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U884 ( .A(KEYINPUT84), .B(G44), .ZN(n799) );
  XNOR2_X1 U885 ( .A(n799), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U886 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NAND2_X1 U887 ( .A1(G483), .A2(G661), .ZN(n808) );
  NOR2_X1 U888 ( .A1(G220), .A2(G219), .ZN(n801) );
  XNOR2_X1 U889 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n800) );
  XNOR2_X1 U890 ( .A(n801), .B(n800), .ZN(n802) );
  NOR2_X1 U891 ( .A1(G218), .A2(n802), .ZN(n803) );
  NAND2_X1 U892 ( .A1(G96), .A2(n803), .ZN(n823) );
  NAND2_X1 U893 ( .A1(n823), .A2(G2106), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G69), .A2(G120), .ZN(n804) );
  NOR2_X1 U895 ( .A1(G237), .A2(n804), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G108), .A2(n805), .ZN(n824) );
  NAND2_X1 U897 ( .A1(n824), .A2(G567), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n825) );
  NOR2_X1 U899 ( .A1(n808), .A2(n825), .ZN(n809) );
  XNOR2_X1 U900 ( .A(n809), .B(KEYINPUT86), .ZN(n822) );
  NAND2_X1 U901 ( .A1(G36), .A2(n822), .ZN(G176) );
  XNOR2_X1 U902 ( .A(G1341), .B(G2454), .ZN(n810) );
  XNOR2_X1 U903 ( .A(n810), .B(G2430), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n811), .B(G1348), .ZN(n817) );
  XOR2_X1 U905 ( .A(G2443), .B(G2427), .Z(n813) );
  XNOR2_X1 U906 ( .A(G2438), .B(G2446), .ZN(n812) );
  XNOR2_X1 U907 ( .A(n813), .B(n812), .ZN(n815) );
  XOR2_X1 U908 ( .A(G2451), .B(G2435), .Z(n814) );
  XNOR2_X1 U909 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n817), .B(n816), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n818), .A2(G14), .ZN(n897) );
  XNOR2_X1 U912 ( .A(KEYINPUT101), .B(n897), .ZN(G401) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U915 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(G188) );
  NOR2_X1 U918 ( .A1(n824), .A2(n823), .ZN(G325) );
  XOR2_X1 U919 ( .A(KEYINPUT102), .B(G325), .Z(G261) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  INV_X1 U924 ( .A(n825), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2096), .B(G2090), .Z(n827) );
  XNOR2_X1 U926 ( .A(G2067), .B(G2072), .ZN(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n837) );
  XOR2_X1 U928 ( .A(KEYINPUT42), .B(KEYINPUT103), .Z(n829) );
  XNOR2_X1 U929 ( .A(KEYINPUT104), .B(KEYINPUT106), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U931 ( .A(G2100), .B(KEYINPUT43), .Z(n831) );
  XNOR2_X1 U932 ( .A(G2678), .B(KEYINPUT105), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U934 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U935 ( .A(G2084), .B(G2078), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U937 ( .A(n837), .B(n836), .Z(G227) );
  XOR2_X1 U938 ( .A(G1961), .B(G1966), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1981), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U941 ( .A(G1956), .B(G1971), .Z(n841) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1976), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U944 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2474), .B(KEYINPUT41), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U947 ( .A(G1991), .B(KEYINPUT107), .Z(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U949 ( .A1(G100), .A2(n869), .ZN(n849) );
  NAND2_X1 U950 ( .A1(G136), .A2(n871), .ZN(n848) );
  NAND2_X1 U951 ( .A1(n849), .A2(n848), .ZN(n855) );
  NAND2_X1 U952 ( .A1(G124), .A2(n865), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n850), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U954 ( .A1(n866), .A2(G112), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n851), .B(KEYINPUT108), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U957 ( .A1(n855), .A2(n854), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G103), .A2(n869), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G139), .A2(n871), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n865), .A2(G127), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G115), .A2(n866), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U964 ( .A(KEYINPUT47), .B(n860), .Z(n861) );
  NOR2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(KEYINPUT111), .B(n863), .Z(n910) );
  XNOR2_X1 U967 ( .A(n910), .B(n864), .ZN(n881) );
  NAND2_X1 U968 ( .A1(n865), .A2(G130), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G118), .A2(n866), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n876) );
  NAND2_X1 U971 ( .A1(n869), .A2(G106), .ZN(n870) );
  XOR2_X1 U972 ( .A(KEYINPUT109), .B(n870), .Z(n873) );
  NAND2_X1 U973 ( .A1(n871), .A2(G142), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U978 ( .A(G164), .B(n879), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(n889) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  XOR2_X1 U981 ( .A(n882), .B(KEYINPUT110), .Z(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n887) );
  XOR2_X1 U983 ( .A(G160), .B(G162), .Z(n885) );
  XNOR2_X1 U984 ( .A(n904), .B(n885), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U987 ( .A1(G37), .A2(n890), .ZN(G395) );
  INV_X1 U988 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U989 ( .A(n958), .B(KEYINPUT112), .ZN(n892) );
  XNOR2_X1 U990 ( .A(G171), .B(n970), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n895) );
  XNOR2_X1 U992 ( .A(G286), .B(n893), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U994 ( .A1(G37), .A2(n896), .ZN(G397) );
  NAND2_X1 U995 ( .A1(G319), .A2(n897), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n898) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(n898), .Z(n899) );
  XNOR2_X1 U998 ( .A(n899), .B(KEYINPUT49), .ZN(n900) );
  NOR2_X1 U999 ( .A1(n901), .A2(n900), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1004 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n927) );
  XNOR2_X1 U1005 ( .A(G160), .B(G2084), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U1007 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n921) );
  XOR2_X1 U1009 ( .A(G2072), .B(n910), .Z(n912) );
  XOR2_X1 U1010 ( .A(G164), .B(G2078), .Z(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(KEYINPUT114), .B(n913), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(KEYINPUT50), .ZN(n919) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1016 ( .A(KEYINPUT51), .B(n917), .Z(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1022 ( .A1(KEYINPUT55), .A2(n928), .ZN(n929) );
  XOR2_X1 U1023 ( .A(KEYINPUT116), .B(n929), .Z(n930) );
  NAND2_X1 U1024 ( .A1(G29), .A2(n930), .ZN(n1014) );
  XOR2_X1 U1025 ( .A(G2090), .B(G35), .Z(n934) );
  XNOR2_X1 U1026 ( .A(KEYINPUT54), .B(G34), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(KEYINPUT119), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(G2084), .B(n932), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n949) );
  XNOR2_X1 U1030 ( .A(G1996), .B(G32), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(G1991), .B(G25), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1033 ( .A(G2072), .B(G33), .Z(n937) );
  NAND2_X1 U1034 ( .A1(n937), .A2(G28), .ZN(n940) );
  XOR2_X1 U1035 ( .A(KEYINPUT117), .B(G2067), .Z(n938) );
  XNOR2_X1 U1036 ( .A(G26), .B(n938), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(G27), .B(n943), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT118), .B(n944), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT53), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT55), .B(n950), .ZN(n952) );
  INV_X1 U1045 ( .A(G29), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(G11), .ZN(n1012) );
  XNOR2_X1 U1048 ( .A(G16), .B(KEYINPUT56), .ZN(n981) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G168), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT120), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT57), .B(n957), .ZN(n979) );
  XNOR2_X1 U1053 ( .A(n958), .B(G1341), .ZN(n977) );
  XNOR2_X1 U1054 ( .A(G1956), .B(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(G1971), .A2(G303), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n966), .B(KEYINPUT121), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(KEYINPUT122), .B(n969), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G1348), .B(n970), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G301), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT123), .B(n975), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n1010) );
  INV_X1 U1070 ( .A(G16), .ZN(n1008) );
  XNOR2_X1 U1071 ( .A(KEYINPUT125), .B(G1981), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n982), .B(G6), .ZN(n987) );
  XOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .Z(n983) );
  XNOR2_X1 U1074 ( .A(G4), .B(n983), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(G19), .B(G1341), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G20), .B(n988), .Z(n989) );
  XNOR2_X1 U1079 ( .A(KEYINPUT124), .B(n989), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(KEYINPUT126), .B(n992), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n993), .B(KEYINPUT60), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G21), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G1961), .B(G5), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1005) );
  XOR2_X1 U1087 ( .A(G1986), .B(G24), .Z(n1001) );
  XNOR2_X1 U1088 ( .A(G1976), .B(G23), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(KEYINPUT127), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1015), .Z(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

