

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(KEYINPUT17), .B(n523), .Z(n892) );
  NOR2_X1 U552 ( .A1(n972), .A2(n698), .ZN(n699) );
  OR2_X1 U553 ( .A1(n767), .A2(n776), .ZN(n518) );
  INV_X1 U554 ( .A(n724), .ZN(n703) );
  NOR2_X1 U555 ( .A1(G299), .A2(n718), .ZN(n714) );
  XNOR2_X1 U556 ( .A(n702), .B(KEYINPUT94), .ZN(n724) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U558 ( .A(n723), .B(n722), .ZN(n729) );
  NAND2_X1 U559 ( .A1(n518), .A2(n963), .ZN(n768) );
  NAND2_X1 U560 ( .A1(G160), .A2(G40), .ZN(n796) );
  INV_X1 U561 ( .A(KEYINPUT13), .ZN(n579) );
  XNOR2_X1 U562 ( .A(KEYINPUT65), .B(n528), .ZN(n651) );
  NOR2_X1 U563 ( .A1(G651), .A2(n533), .ZN(n656) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n532), .Z(n660) );
  NAND2_X1 U565 ( .A1(n586), .A2(n585), .ZN(n972) );
  AND2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U567 ( .A1(n888), .A2(G113), .ZN(n522) );
  INV_X1 U568 ( .A(G2105), .ZN(n519) );
  AND2_X1 U569 ( .A1(n519), .A2(G2104), .ZN(n891) );
  NAND2_X1 U570 ( .A1(G101), .A2(n891), .ZN(n520) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n520), .Z(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NAND2_X1 U574 ( .A1(G137), .A2(n892), .ZN(n525) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n519), .ZN(n887) );
  NAND2_X1 U576 ( .A1(G125), .A2(n887), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n527), .A2(n526), .ZN(G160) );
  INV_X1 U579 ( .A(G651), .ZN(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n533) );
  OR2_X1 U581 ( .A1(n531), .A2(n533), .ZN(n528) );
  NAND2_X1 U582 ( .A1(G78), .A2(n651), .ZN(n530) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U584 ( .A1(G91), .A2(n652), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n530), .A2(n529), .ZN(n537) );
  NOR2_X1 U586 ( .A1(G543), .A2(n531), .ZN(n532) );
  NAND2_X1 U587 ( .A1(G65), .A2(n660), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G53), .A2(n656), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U590 ( .A1(n537), .A2(n536), .ZN(G299) );
  NAND2_X1 U591 ( .A1(n892), .A2(G138), .ZN(n544) );
  NAND2_X1 U592 ( .A1(G126), .A2(n887), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G114), .A2(n888), .ZN(n538) );
  AND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n891), .A2(G102), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n540), .B(KEYINPUT92), .ZN(n541) );
  AND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  AND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(G164) );
  XOR2_X1 U599 ( .A(G2443), .B(G2446), .Z(n546) );
  XNOR2_X1 U600 ( .A(G2427), .B(G2451), .ZN(n545) );
  XNOR2_X1 U601 ( .A(n546), .B(n545), .ZN(n552) );
  XOR2_X1 U602 ( .A(G2430), .B(G2454), .Z(n548) );
  XNOR2_X1 U603 ( .A(G1348), .B(G1341), .ZN(n547) );
  XNOR2_X1 U604 ( .A(n548), .B(n547), .ZN(n550) );
  XOR2_X1 U605 ( .A(G2435), .B(G2438), .Z(n549) );
  XNOR2_X1 U606 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U607 ( .A(n552), .B(n551), .Z(n553) );
  AND2_X1 U608 ( .A1(G14), .A2(n553), .ZN(G401) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  INV_X1 U611 ( .A(G120), .ZN(G236) );
  INV_X1 U612 ( .A(G69), .ZN(G235) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  NAND2_X1 U614 ( .A1(G64), .A2(n660), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G52), .A2(n656), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G77), .A2(n651), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G90), .A2(n652), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  XNOR2_X1 U621 ( .A(KEYINPUT68), .B(n559), .ZN(n560) );
  NOR2_X1 U622 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U623 ( .A1(G63), .A2(n660), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G51), .A2(n656), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(n564), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n652), .A2(G89), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G76), .A2(n651), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U631 ( .A(n568), .B(KEYINPUT5), .Z(n569) );
  NOR2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT7), .B(n571), .Z(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT75), .B(n572), .Z(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U638 ( .A(G223), .B(KEYINPUT70), .Z(n828) );
  NAND2_X1 U639 ( .A1(n828), .A2(G567), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U641 ( .A1(G68), .A2(n651), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G81), .A2(n652), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n575), .B(KEYINPUT72), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G56), .A2(n660), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT71), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n582), .B(KEYINPUT14), .ZN(n583) );
  NOR2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n656), .A2(G43), .ZN(n585) );
  XNOR2_X1 U652 ( .A(G860), .B(KEYINPUT73), .ZN(n599) );
  OR2_X1 U653 ( .A1(n972), .A2(n599), .ZN(G153) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U656 ( .A1(G54), .A2(n656), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G79), .A2(n651), .ZN(n588) );
  NAND2_X1 U658 ( .A1(G66), .A2(n660), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n652), .A2(G92), .ZN(n589) );
  XOR2_X1 U661 ( .A(KEYINPUT74), .B(n589), .Z(n590) );
  NOR2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(KEYINPUT15), .ZN(n976) );
  INV_X1 U665 ( .A(n976), .ZN(n602) );
  INV_X1 U666 ( .A(G868), .ZN(n672) );
  NAND2_X1 U667 ( .A1(n602), .A2(n672), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(G284) );
  NOR2_X1 U669 ( .A1(G286), .A2(n672), .ZN(n598) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U672 ( .A1(G559), .A2(n599), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT76), .B(n600), .Z(n601) );
  NOR2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT77), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U677 ( .A1(n976), .A2(G868), .ZN(n605) );
  XNOR2_X1 U678 ( .A(KEYINPUT78), .B(n605), .ZN(n606) );
  NOR2_X1 U679 ( .A1(G559), .A2(n606), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT79), .B(n607), .Z(n609) );
  NOR2_X1 U681 ( .A1(G868), .A2(n972), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G99), .A2(n891), .ZN(n611) );
  NAND2_X1 U684 ( .A1(G111), .A2(n888), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n617) );
  NAND2_X1 U686 ( .A1(G123), .A2(n887), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n612), .B(KEYINPUT18), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G135), .A2(n892), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n613), .B(KEYINPUT80), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n909) );
  XNOR2_X1 U692 ( .A(G2096), .B(n909), .ZN(n619) );
  INV_X1 U693 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G55), .A2(n656), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT82), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n651), .A2(G80), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U699 ( .A1(G93), .A2(n652), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G67), .A2(n660), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n671) );
  NAND2_X1 U703 ( .A1(G559), .A2(n976), .ZN(n627) );
  XOR2_X1 U704 ( .A(n972), .B(n627), .Z(n668) );
  XNOR2_X1 U705 ( .A(KEYINPUT81), .B(n668), .ZN(n628) );
  NOR2_X1 U706 ( .A1(G860), .A2(n628), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n671), .B(n629), .ZN(G145) );
  NAND2_X1 U708 ( .A1(G75), .A2(n651), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G88), .A2(n652), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G50), .A2(n656), .ZN(n632) );
  XNOR2_X1 U712 ( .A(KEYINPUT85), .B(n632), .ZN(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n660), .A2(G62), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(G303) );
  INV_X1 U716 ( .A(G303), .ZN(G166) );
  XOR2_X1 U717 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n638) );
  NAND2_X1 U718 ( .A1(G73), .A2(n651), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n638), .B(n637), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G86), .A2(n652), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G48), .A2(n656), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n660), .A2(G61), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G49), .A2(n656), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U729 ( .A(KEYINPUT83), .B(n647), .Z(n648) );
  NOR2_X1 U730 ( .A1(n660), .A2(n648), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n533), .A2(G87), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U733 ( .A1(G72), .A2(n651), .ZN(n654) );
  NAND2_X1 U734 ( .A1(G85), .A2(n652), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U736 ( .A(KEYINPUT66), .B(n655), .ZN(n659) );
  NAND2_X1 U737 ( .A1(G47), .A2(n656), .ZN(n657) );
  XNOR2_X1 U738 ( .A(KEYINPUT67), .B(n657), .ZN(n658) );
  NOR2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n660), .A2(G60), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n662), .A2(n661), .ZN(G290) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(G299), .ZN(n667) );
  XNOR2_X1 U743 ( .A(G166), .B(n671), .ZN(n665) );
  XNOR2_X1 U744 ( .A(G305), .B(G288), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n663), .B(G290), .ZN(n664) );
  XNOR2_X1 U746 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n667), .B(n666), .ZN(n837) );
  XNOR2_X1 U748 ( .A(n668), .B(n837), .ZN(n669) );
  XNOR2_X1 U749 ( .A(KEYINPUT86), .B(n669), .ZN(n670) );
  NOR2_X1 U750 ( .A1(n672), .A2(n670), .ZN(n674) );
  AND2_X1 U751 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U752 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U757 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G235), .A2(G236), .ZN(n679) );
  XNOR2_X1 U761 ( .A(n679), .B(KEYINPUT89), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G237), .A2(n680), .ZN(n681) );
  XNOR2_X1 U763 ( .A(KEYINPUT90), .B(n681), .ZN(n682) );
  NAND2_X1 U764 ( .A1(n682), .A2(G108), .ZN(n834) );
  AND2_X1 U765 ( .A1(G567), .A2(n834), .ZN(n689) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n684) );
  XNOR2_X1 U767 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n683) );
  XNOR2_X1 U768 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X1 U769 ( .A1(n685), .A2(G218), .ZN(n686) );
  NAND2_X1 U770 ( .A1(G96), .A2(n686), .ZN(n833) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n833), .ZN(n687) );
  XOR2_X1 U772 ( .A(KEYINPUT88), .B(n687), .Z(n688) );
  NOR2_X1 U773 ( .A1(n689), .A2(n688), .ZN(G319) );
  INV_X1 U774 ( .A(G319), .ZN(n902) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U776 ( .A1(n902), .A2(n690), .ZN(n832) );
  NAND2_X1 U777 ( .A1(G36), .A2(n832), .ZN(n691) );
  XOR2_X1 U778 ( .A(KEYINPUT91), .B(n691), .Z(G176) );
  XNOR2_X1 U779 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n827) );
  INV_X1 U780 ( .A(n796), .ZN(n692) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n795) );
  NAND2_X1 U782 ( .A1(n692), .A2(n795), .ZN(n702) );
  INV_X1 U783 ( .A(n702), .ZN(n725) );
  INV_X1 U784 ( .A(n725), .ZN(n740) );
  NAND2_X1 U785 ( .A1(G8), .A2(n740), .ZN(n776) );
  INV_X1 U786 ( .A(G1996), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n702), .A2(n693), .ZN(n695) );
  XOR2_X1 U788 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n694) );
  XNOR2_X1 U789 ( .A(n695), .B(n694), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n740), .A2(G1341), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U792 ( .A(n699), .B(KEYINPUT64), .ZN(n701) );
  NOR2_X1 U793 ( .A1(n976), .A2(n701), .ZN(n700) );
  XNOR2_X1 U794 ( .A(n700), .B(KEYINPUT97), .ZN(n709) );
  NAND2_X1 U795 ( .A1(n976), .A2(n701), .ZN(n707) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n740), .ZN(n705) );
  NAND2_X1 U797 ( .A1(G2067), .A2(n703), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n717) );
  INV_X1 U801 ( .A(KEYINPUT98), .ZN(n715) );
  INV_X1 U802 ( .A(G2072), .ZN(n920) );
  NOR2_X1 U803 ( .A1(n724), .A2(n920), .ZN(n711) );
  XOR2_X1 U804 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n710) );
  XNOR2_X1 U805 ( .A(n711), .B(n710), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n724), .A2(G1956), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n718) );
  XNOR2_X1 U808 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U810 ( .A1(G299), .A2(n718), .ZN(n719) );
  XNOR2_X1 U811 ( .A(n719), .B(KEYINPUT28), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .Z(n943) );
  NOR2_X1 U814 ( .A1(n943), .A2(n724), .ZN(n727) );
  NOR2_X1 U815 ( .A1(n725), .A2(G1961), .ZN(n726) );
  NOR2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n730) );
  OR2_X1 U817 ( .A1(n730), .A2(G301), .ZN(n728) );
  NAND2_X1 U818 ( .A1(n729), .A2(n728), .ZN(n739) );
  NAND2_X1 U819 ( .A1(n730), .A2(G301), .ZN(n731) );
  XNOR2_X1 U820 ( .A(n731), .B(KEYINPUT99), .ZN(n736) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n776), .ZN(n754) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n740), .ZN(n751) );
  NOR2_X1 U823 ( .A1(n754), .A2(n751), .ZN(n732) );
  NAND2_X1 U824 ( .A1(G8), .A2(n732), .ZN(n733) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n734), .A2(G168), .ZN(n735) );
  NOR2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U828 ( .A(KEYINPUT31), .B(n737), .Z(n738) );
  NAND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n752) );
  NAND2_X1 U830 ( .A1(n752), .A2(G286), .ZN(n749) );
  INV_X1 U831 ( .A(G8), .ZN(n747) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n776), .ZN(n742) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U835 ( .A(KEYINPUT100), .B(n743), .Z(n744) );
  NOR2_X1 U836 ( .A1(G166), .A2(n744), .ZN(n745) );
  XNOR2_X1 U837 ( .A(n745), .B(KEYINPUT101), .ZN(n746) );
  OR2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U840 ( .A(n750), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U841 ( .A1(G8), .A2(n751), .ZN(n756) );
  INV_X1 U842 ( .A(n752), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n772) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n766), .A2(n759), .ZN(n971) );
  XNOR2_X1 U849 ( .A(KEYINPUT102), .B(n971), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n772), .A2(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G288), .A2(G1976), .ZN(n761) );
  XOR2_X1 U852 ( .A(KEYINPUT103), .B(n761), .Z(n977) );
  NAND2_X1 U853 ( .A1(n762), .A2(n977), .ZN(n763) );
  XNOR2_X1 U854 ( .A(n763), .B(KEYINPUT104), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n776), .A2(n764), .ZN(n765) );
  NOR2_X1 U856 ( .A1(KEYINPUT33), .A2(n765), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n963) );
  NOR2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n781) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U861 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n773), .A2(n776), .ZN(n779) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XOR2_X1 U865 ( .A(n774), .B(KEYINPUT24), .Z(n775) );
  NOR2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U867 ( .A(KEYINPUT93), .B(n777), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n808) );
  NAND2_X1 U870 ( .A1(G141), .A2(n892), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G117), .A2(n888), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n891), .A2(G105), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n887), .A2(G129), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n873) );
  AND2_X1 U878 ( .A1(n873), .A2(G1996), .ZN(n910) );
  NAND2_X1 U879 ( .A1(G95), .A2(n891), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G131), .A2(n892), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G119), .A2(n887), .ZN(n792) );
  NAND2_X1 U883 ( .A1(G107), .A2(n888), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n868) );
  INV_X1 U886 ( .A(G1991), .ZN(n940) );
  NOR2_X1 U887 ( .A1(n868), .A2(n940), .ZN(n912) );
  OR2_X1 U888 ( .A1(n910), .A2(n912), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n822) );
  NAND2_X1 U890 ( .A1(n797), .A2(n822), .ZN(n811) );
  XNOR2_X1 U891 ( .A(KEYINPUT37), .B(G2067), .ZN(n819) );
  NAND2_X1 U892 ( .A1(G104), .A2(n891), .ZN(n799) );
  NAND2_X1 U893 ( .A1(G140), .A2(n892), .ZN(n798) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U895 ( .A(KEYINPUT34), .B(n800), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G128), .A2(n887), .ZN(n802) );
  NAND2_X1 U897 ( .A1(G116), .A2(n888), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U899 ( .A(KEYINPUT35), .B(n803), .Z(n804) );
  NOR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U901 ( .A(KEYINPUT36), .B(n806), .ZN(n872) );
  NOR2_X1 U902 ( .A1(n819), .A2(n872), .ZN(n916) );
  NAND2_X1 U903 ( .A1(n822), .A2(n916), .ZN(n817) );
  NAND2_X1 U904 ( .A1(n811), .A2(n817), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n810) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n980) );
  NAND2_X1 U907 ( .A1(n980), .A2(n822), .ZN(n809) );
  NAND2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n825) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n873), .ZN(n925) );
  INV_X1 U910 ( .A(n811), .ZN(n814) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n812) );
  AND2_X1 U912 ( .A1(n940), .A2(n868), .ZN(n911) );
  NOR2_X1 U913 ( .A1(n812), .A2(n911), .ZN(n813) );
  NOR2_X1 U914 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U915 ( .A1(n925), .A2(n815), .ZN(n816) );
  XNOR2_X1 U916 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U917 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n819), .A2(n872), .ZN(n932) );
  NAND2_X1 U919 ( .A1(n820), .A2(n932), .ZN(n821) );
  NAND2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U921 ( .A(KEYINPUT105), .B(n823), .Z(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n827), .B(n826), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n830) );
  XOR2_X1 U928 ( .A(KEYINPUT107), .B(n830), .Z(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(n972), .B(G286), .ZN(n836) );
  XNOR2_X1 U936 ( .A(G171), .B(n976), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  NOR2_X1 U939 ( .A1(G37), .A2(n839), .ZN(G397) );
  XOR2_X1 U940 ( .A(G2096), .B(G2678), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2090), .B(KEYINPUT43), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n842), .B(KEYINPUT42), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U946 ( .A(KEYINPUT108), .B(G2100), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1986), .B(G1966), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1981), .B(G1976), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(n851), .B(G2474), .Z(n853) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U956 ( .A(KEYINPUT41), .B(G1971), .Z(n855) );
  XNOR2_X1 U957 ( .A(G1961), .B(G1956), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G112), .A2(n888), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G100), .A2(n891), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G136), .A2(n892), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n864) );
  XOR2_X1 U964 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n861) );
  NAND2_X1 U965 ( .A1(G124), .A2(n887), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U967 ( .A(KEYINPUT109), .B(n862), .Z(n863) );
  NOR2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT111), .ZN(G162) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U972 ( .A(n868), .B(KEYINPUT112), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n875) );
  XOR2_X1 U975 ( .A(G164), .B(n873), .Z(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n876), .B(n909), .Z(n878) );
  XNOR2_X1 U978 ( .A(G160), .B(G162), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n900) );
  NAND2_X1 U980 ( .A1(G103), .A2(n891), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G139), .A2(n892), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n888), .A2(G115), .ZN(n881) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n881), .Z(n883) );
  NAND2_X1 U985 ( .A1(n887), .A2(G127), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n919) );
  NAND2_X1 U989 ( .A1(G130), .A2(n887), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G118), .A2(n888), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U992 ( .A1(G106), .A2(n891), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G142), .A2(n892), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(KEYINPUT45), .B(n895), .Z(n896) );
  NOR2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n919), .B(n898), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U999 ( .A1(G37), .A2(n901), .ZN(G395) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n902), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G397), .A2(n904), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n907), .A2(G395), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(KEYINPUT114), .ZN(G308) );
  INV_X1 U1007 ( .A(G308), .ZN(G225) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n918) );
  XNOR2_X1 U1009 ( .A(G160), .B(G2084), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n930) );
  XOR2_X1 U1014 ( .A(G164), .B(G2078), .Z(n922) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(KEYINPUT50), .B(n923), .ZN(n928) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n926), .Z(n927) );
  NAND2_X1 U1021 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(n933), .B(KEYINPUT52), .ZN(n934) );
  XNOR2_X1 U1025 ( .A(KEYINPUT115), .B(n934), .ZN(n935) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n958) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n958), .ZN(n936) );
  NAND2_X1 U1028 ( .A1(n936), .A2(G29), .ZN(n1020) );
  XOR2_X1 U1029 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n957) );
  XNOR2_X1 U1030 ( .A(G2090), .B(G35), .ZN(n952) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(G2072), .B(G33), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n939), .B(KEYINPUT116), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(n940), .B(G25), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n949) );
  XNOR2_X1 U1037 ( .A(G1996), .B(G32), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(n943), .B(G27), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1040 ( .A(KEYINPUT117), .B(n946), .Z(n947) );
  NAND2_X1 U1041 ( .A1(n947), .A2(G28), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT53), .B(n950), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G2084), .B(G34), .Z(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(n953), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n957), .B(n956), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(n959), .B(n958), .ZN(n961) );
  INV_X1 U1050 ( .A(G29), .ZN(n960) );
  NAND2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n962), .ZN(n1018) );
  XNOR2_X1 U1053 ( .A(G16), .B(KEYINPUT56), .ZN(n987) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n964) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(KEYINPUT57), .B(n965), .ZN(n985) );
  XNOR2_X1 U1057 ( .A(G171), .B(G1961), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(G1971), .A2(G303), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(G1956), .B(G299), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(G1341), .B(n972), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT120), .B(n973), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n982) );
  XNOR2_X1 U1066 ( .A(n976), .B(G1348), .ZN(n978) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1070 ( .A(KEYINPUT121), .B(n983), .ZN(n984) );
  NAND2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1072 ( .A1(n987), .A2(n986), .ZN(n1016) );
  INV_X1 U1073 ( .A(G16), .ZN(n1014) );
  XOR2_X1 U1074 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n994) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G1986), .B(G24), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G1976), .B(KEYINPUT125), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(n990), .B(G23), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n994), .B(n993), .ZN(n1009) );
  XNOR2_X1 U1082 ( .A(KEYINPUT123), .B(G1981), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n995), .B(G6), .ZN(n1002) );
  XOR2_X1 U1084 ( .A(KEYINPUT124), .B(G4), .Z(n997) );
  XNOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n997), .B(n996), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT122), .B(G1956), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(G20), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G19), .B(G1341), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G21), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G5), .B(G1961), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(n1021), .B(KEYINPUT127), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1022), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

