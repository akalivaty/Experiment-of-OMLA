

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  INV_X1 U324 ( .A(n564), .ZN(n388) );
  XNOR2_X1 U325 ( .A(n397), .B(G50GAT), .ZN(n398) );
  XNOR2_X1 U326 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U327 ( .A(n402), .B(n292), .ZN(n403) );
  XNOR2_X1 U328 ( .A(n450), .B(n293), .ZN(n451) );
  XNOR2_X1 U329 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U330 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n292) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U332 ( .A(KEYINPUT18), .B(KEYINPUT88), .Z(n294) );
  XOR2_X1 U333 ( .A(KEYINPUT54), .B(n559), .Z(n295) );
  INV_X1 U334 ( .A(KEYINPUT46), .ZN(n511) );
  XNOR2_X1 U335 ( .A(n511), .B(KEYINPUT114), .ZN(n512) );
  XNOR2_X1 U336 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U337 ( .A(n520), .B(n519), .ZN(n523) );
  XOR2_X1 U338 ( .A(G36GAT), .B(n374), .Z(n375) );
  XNOR2_X1 U339 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U340 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n526) );
  XOR2_X1 U341 ( .A(G190GAT), .B(G218GAT), .Z(n444) );
  XNOR2_X1 U342 ( .A(n331), .B(n330), .ZN(n334) );
  XNOR2_X1 U343 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U344 ( .A(G169GAT), .B(G8GAT), .Z(n383) );
  XNOR2_X1 U345 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U346 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U347 ( .A(KEYINPUT19), .B(n311), .ZN(n374) );
  XNOR2_X1 U348 ( .A(n465), .B(G106GAT), .ZN(n466) );
  XNOR2_X1 U349 ( .A(KEYINPUT40), .B(G43GAT), .ZN(n460) );
  XNOR2_X1 U350 ( .A(n467), .B(n466), .ZN(G1339GAT) );
  XNOR2_X1 U351 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT87), .B(G176GAT), .Z(n297) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n309) );
  XOR2_X1 U355 ( .A(G120GAT), .B(G71GAT), .Z(n338) );
  XOR2_X1 U356 ( .A(KEYINPUT86), .B(G99GAT), .Z(n299) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U359 ( .A(n338), .B(n300), .Z(n302) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U362 ( .A(n303), .B(KEYINPUT89), .Z(n307) );
  XOR2_X1 U363 ( .A(G127GAT), .B(KEYINPUT0), .Z(n305) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(G134GAT), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n352) );
  XNOR2_X1 U366 ( .A(n352), .B(KEYINPUT20), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n312) );
  XNOR2_X1 U369 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n294), .B(n310), .ZN(n311) );
  XNOR2_X2 U371 ( .A(n312), .B(n374), .ZN(n564) );
  XOR2_X1 U372 ( .A(G43GAT), .B(G29GAT), .Z(n314) );
  XNOR2_X1 U373 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U375 ( .A(n315), .B(KEYINPUT69), .Z(n317) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n443) );
  XOR2_X1 U378 ( .A(G113GAT), .B(G197GAT), .Z(n319) );
  XOR2_X1 U379 ( .A(G141GAT), .B(G22GAT), .Z(n392) );
  XNOR2_X1 U380 ( .A(n392), .B(n383), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n324) );
  INV_X1 U382 ( .A(n324), .ZN(n323) );
  XOR2_X1 U383 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n321) );
  XNOR2_X1 U384 ( .A(KEYINPUT71), .B(KEYINPUT67), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n325) );
  INV_X1 U386 ( .A(n325), .ZN(n322) );
  NAND2_X1 U387 ( .A1(n323), .A2(n322), .ZN(n327) );
  NAND2_X1 U388 ( .A1(n325), .A2(n324), .ZN(n326) );
  NAND2_X1 U389 ( .A1(n327), .A2(n326), .ZN(n331) );
  AND2_X1 U390 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  INV_X1 U391 ( .A(KEYINPUT68), .ZN(n328) );
  XNOR2_X1 U392 ( .A(G15GAT), .B(G1GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n332), .B(KEYINPUT70), .ZN(n434) );
  XNOR2_X1 U394 ( .A(n434), .B(KEYINPUT30), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n443), .B(n335), .ZN(n510) );
  XOR2_X1 U397 ( .A(n510), .B(KEYINPUT72), .Z(n566) );
  XOR2_X1 U398 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n337) );
  XNOR2_X1 U399 ( .A(G204GAT), .B(KEYINPUT76), .ZN(n336) );
  XOR2_X1 U400 ( .A(n337), .B(n336), .Z(n351) );
  XNOR2_X1 U401 ( .A(G176GAT), .B(G64GAT), .ZN(n386) );
  XOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT13), .Z(n433) );
  XNOR2_X1 U403 ( .A(n386), .B(n433), .ZN(n340) );
  XOR2_X1 U404 ( .A(G148GAT), .B(G78GAT), .Z(n391) );
  XNOR2_X1 U405 ( .A(n338), .B(n391), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U407 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n342) );
  NAND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U410 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U411 ( .A(KEYINPUT75), .B(G92GAT), .Z(n346) );
  XNOR2_X1 U412 ( .A(G99GAT), .B(G85GAT), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U414 ( .A(G106GAT), .B(n347), .Z(n442) );
  XNOR2_X1 U415 ( .A(n442), .B(KEYINPUT33), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n521) );
  INV_X1 U418 ( .A(n521), .ZN(n586) );
  NOR2_X1 U419 ( .A1(n566), .A2(n586), .ZN(n473) );
  XOR2_X1 U420 ( .A(G85GAT), .B(n352), .Z(n354) );
  NAND2_X1 U421 ( .A1(G225GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U423 ( .A(G29GAT), .B(n355), .ZN(n371) );
  XOR2_X1 U424 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n357) );
  XNOR2_X1 U425 ( .A(G57GAT), .B(KEYINPUT97), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U427 ( .A(G148GAT), .B(G162GAT), .Z(n359) );
  XNOR2_X1 U428 ( .A(G141GAT), .B(G120GAT), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n369) );
  XOR2_X1 U431 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n367) );
  XNOR2_X1 U432 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n362), .B(KEYINPUT2), .ZN(n402) );
  XOR2_X1 U434 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n364) );
  XNOR2_X1 U435 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n402), .B(n365), .ZN(n366) );
  XNOR2_X1 U438 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n560) );
  XOR2_X1 U441 ( .A(G204GAT), .B(G211GAT), .Z(n373) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n373), .B(n372), .ZN(n396) );
  XOR2_X1 U444 ( .A(G92GAT), .B(n396), .Z(n376) );
  XNOR2_X1 U445 ( .A(n376), .B(n375), .ZN(n378) );
  INV_X1 U446 ( .A(n378), .ZN(n377) );
  NAND2_X1 U447 ( .A1(n444), .A2(n377), .ZN(n381) );
  INV_X1 U448 ( .A(n444), .ZN(n379) );
  NAND2_X1 U449 ( .A1(n379), .A2(n378), .ZN(n380) );
  NAND2_X1 U450 ( .A1(n381), .A2(n380), .ZN(n385) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n557) );
  OR2_X1 U453 ( .A1(n388), .A2(n557), .ZN(n407) );
  XOR2_X1 U454 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n390) );
  XNOR2_X1 U455 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n406) );
  XOR2_X1 U457 ( .A(G106GAT), .B(G218GAT), .Z(n394) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U460 ( .A(n395), .B(KEYINPUT92), .Z(n401) );
  XOR2_X1 U461 ( .A(KEYINPUT77), .B(G162GAT), .Z(n445) );
  XOR2_X1 U462 ( .A(n445), .B(n396), .Z(n399) );
  NAND2_X1 U463 ( .A1(G228GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n404) );
  XOR2_X1 U465 ( .A(n406), .B(n405), .Z(n562) );
  NAND2_X1 U466 ( .A1(n407), .A2(n562), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT25), .ZN(n410) );
  INV_X1 U468 ( .A(KEYINPUT98), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n413) );
  NOR2_X1 U470 ( .A1(n564), .A2(n562), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n411), .B(KEYINPUT26), .ZN(n580) );
  INV_X1 U472 ( .A(n557), .ZN(n506) );
  XNOR2_X1 U473 ( .A(KEYINPUT27), .B(n506), .ZN(n416) );
  NAND2_X1 U474 ( .A1(n580), .A2(n416), .ZN(n412) );
  NAND2_X1 U475 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U476 ( .A(KEYINPUT99), .B(n414), .ZN(n415) );
  NOR2_X1 U477 ( .A1(n560), .A2(n415), .ZN(n419) );
  NAND2_X1 U478 ( .A1(n416), .A2(n560), .ZN(n528) );
  XNOR2_X1 U479 ( .A(n562), .B(KEYINPUT28), .ZN(n501) );
  INV_X1 U480 ( .A(n501), .ZN(n530) );
  OR2_X1 U481 ( .A1(n528), .A2(n530), .ZN(n417) );
  NOR2_X1 U482 ( .A1(n564), .A2(n417), .ZN(n418) );
  NOR2_X1 U483 ( .A1(n419), .A2(n418), .ZN(n471) );
  XOR2_X1 U484 ( .A(G211GAT), .B(G71GAT), .Z(n421) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(G183GAT), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U487 ( .A(KEYINPUT84), .B(G64GAT), .Z(n423) );
  XNOR2_X1 U488 ( .A(G8GAT), .B(G127GAT), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U490 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U491 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n427) );
  NAND2_X1 U492 ( .A1(G231GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U494 ( .A(KEYINPUT12), .B(n428), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n440) );
  XOR2_X1 U496 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n432) );
  XNOR2_X1 U497 ( .A(KEYINPUT15), .B(KEYINPUT85), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n432), .B(n431), .ZN(n438) );
  XOR2_X1 U499 ( .A(n433), .B(G78GAT), .Z(n436) );
  XNOR2_X1 U500 ( .A(n434), .B(G155GAT), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U502 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n589) );
  NOR2_X1 U504 ( .A1(n471), .A2(n589), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n441), .B(KEYINPUT104), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT11), .B(n444), .Z(n447) );
  XNOR2_X1 U508 ( .A(G134GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT79), .B(KEYINPUT9), .Z(n449) );
  XNOR2_X1 U511 ( .A(KEYINPUT10), .B(KEYINPUT78), .ZN(n448) );
  XNOR2_X1 U512 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n454), .B(n453), .ZN(n515) );
  INV_X1 U514 ( .A(n515), .ZN(n554) );
  XOR2_X1 U515 ( .A(KEYINPUT80), .B(n554), .Z(n576) );
  INV_X1 U516 ( .A(n576), .ZN(n468) );
  XNOR2_X1 U517 ( .A(KEYINPUT36), .B(n468), .ZN(n592) );
  NAND2_X1 U518 ( .A1(n455), .A2(n592), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n456), .B(KEYINPUT105), .ZN(n457) );
  XOR2_X1 U520 ( .A(KEYINPUT37), .B(n457), .Z(n463) );
  NAND2_X1 U521 ( .A1(n473), .A2(n463), .ZN(n459) );
  XOR2_X1 U522 ( .A(KEYINPUT106), .B(KEYINPUT38), .Z(n458) );
  XNOR2_X2 U523 ( .A(n459), .B(n458), .ZN(n488) );
  NAND2_X1 U524 ( .A1(n564), .A2(n488), .ZN(n461) );
  INV_X1 U525 ( .A(KEYINPUT41), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n462), .B(n521), .ZN(n571) );
  NOR2_X1 U527 ( .A1(n571), .A2(n510), .ZN(n493) );
  NAND2_X1 U528 ( .A1(n493), .A2(n463), .ZN(n464) );
  XNOR2_X2 U529 ( .A(n464), .B(KEYINPUT111), .ZN(n508) );
  NAND2_X1 U530 ( .A1(n508), .A2(n530), .ZN(n467) );
  XOR2_X1 U531 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n465) );
  INV_X1 U532 ( .A(n560), .ZN(n494) );
  INV_X1 U533 ( .A(n589), .ZN(n574) );
  NOR2_X1 U534 ( .A1(n574), .A2(n468), .ZN(n469) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  NOR2_X1 U536 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U537 ( .A(KEYINPUT100), .B(n472), .ZN(n492) );
  NAND2_X1 U538 ( .A1(n473), .A2(n492), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n494), .A2(n480), .ZN(n475) );
  XNOR2_X1 U540 ( .A(KEYINPUT101), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U541 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n557), .A2(n480), .ZN(n477) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n388), .A2(n480), .ZN(n479) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U547 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n501), .A2(n480), .ZN(n481) );
  XOR2_X1 U549 ( .A(KEYINPUT102), .B(n481), .Z(n482) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  NAND2_X1 U551 ( .A1(n488), .A2(n560), .ZN(n485) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n483) );
  XNOR2_X1 U553 ( .A(n483), .B(KEYINPUT39), .ZN(n484) );
  XNOR2_X1 U554 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  XOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT107), .Z(n487) );
  NAND2_X1 U556 ( .A1(n506), .A2(n488), .ZN(n486) );
  XNOR2_X1 U557 ( .A(n487), .B(n486), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n530), .A2(n488), .ZN(n489) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n489), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n491) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n490) );
  XNOR2_X1 U562 ( .A(n491), .B(n490), .ZN(n496) );
  NAND2_X1 U563 ( .A1(n493), .A2(n492), .ZN(n500) );
  NOR2_X1 U564 ( .A1(n494), .A2(n500), .ZN(n495) );
  XOR2_X1 U565 ( .A(n496), .B(n495), .Z(G1332GAT) );
  NOR2_X1 U566 ( .A1(n557), .A2(n500), .ZN(n497) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n497), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n388), .A2(n500), .ZN(n498) );
  XOR2_X1 U569 ( .A(KEYINPUT110), .B(n498), .Z(n499) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n499), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n501), .A2(n500), .ZN(n503) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n502) );
  XNOR2_X1 U573 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n505) );
  NAND2_X1 U575 ( .A1(n560), .A2(n508), .ZN(n504) );
  XNOR2_X1 U576 ( .A(n505), .B(n504), .ZN(G1336GAT) );
  NAND2_X1 U577 ( .A1(n508), .A2(n506), .ZN(n507) );
  XNOR2_X1 U578 ( .A(n507), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U579 ( .A1(n564), .A2(n508), .ZN(n509) );
  XNOR2_X1 U580 ( .A(n509), .B(G99GAT), .ZN(G1338GAT) );
  INV_X1 U581 ( .A(n571), .ZN(n548) );
  NAND2_X1 U582 ( .A1(n510), .A2(n548), .ZN(n513) );
  NOR2_X1 U583 ( .A1(n589), .A2(n514), .ZN(n516) );
  NAND2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n518) );
  XOR2_X1 U585 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n525) );
  NAND2_X1 U587 ( .A1(n592), .A2(n589), .ZN(n520) );
  XOR2_X1 U588 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n519) );
  NAND2_X1 U589 ( .A1(n566), .A2(n521), .ZN(n522) );
  NOR2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n558) );
  NOR2_X1 U593 ( .A1(n558), .A2(n528), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n545), .A2(n564), .ZN(n529) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(KEYINPUT117), .B(n531), .ZN(n540) );
  NOR2_X1 U597 ( .A1(n566), .A2(n540), .ZN(n532) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n532), .Z(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT118), .B(n533), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n571), .A2(n540), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT119), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  NOR2_X1 U604 ( .A1(n574), .A2(n540), .ZN(n538) );
  XNOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U608 ( .A1(n540), .A2(n576), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n542) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT121), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n580), .A2(n545), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n546), .B(KEYINPUT123), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n553), .A2(n510), .ZN(n547) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U618 ( .A1(n553), .A2(n548), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n589), .A2(n553), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT124), .ZN(n556) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U627 ( .A1(n560), .A2(n295), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT64), .ZN(n581) );
  NAND2_X1 U629 ( .A1(n581), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT55), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U632 ( .A1(n566), .A2(n577), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT125), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT126), .Z(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n577), .A2(n571), .ZN(n572) );
  XOR2_X1 U639 ( .A(n573), .B(n572), .Z(G1349GAT) );
  NOR2_X1 U640 ( .A1(n574), .A2(n577), .ZN(n575) );
  XOR2_X1 U641 ( .A(G183GAT), .B(n575), .Z(G1350GAT) );
  OR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT58), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n584) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(KEYINPUT127), .B(n582), .ZN(n591) );
  NAND2_X1 U648 ( .A1(n591), .A2(n510), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G197GAT), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U652 ( .A1(n591), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n589), .A2(n591), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

