

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598;

  XOR2_X1 U323 ( .A(n331), .B(n314), .Z(n540) );
  INV_X1 U324 ( .A(KEYINPUT25), .ZN(n468) );
  XNOR2_X1 U325 ( .A(n468), .B(KEYINPUT96), .ZN(n469) );
  XNOR2_X1 U326 ( .A(G204GAT), .B(KEYINPUT93), .ZN(n334) );
  XNOR2_X1 U327 ( .A(n470), .B(n469), .ZN(n479) );
  XNOR2_X1 U328 ( .A(n335), .B(n334), .ZN(n338) );
  XNOR2_X1 U329 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U330 ( .A(n414), .B(n413), .ZN(n418) );
  INV_X1 U331 ( .A(KEYINPUT41), .ZN(n419) );
  INV_X1 U332 ( .A(G190GAT), .ZN(n461) );
  NOR2_X1 U333 ( .A1(n475), .A2(n460), .ZN(n576) );
  XOR2_X1 U334 ( .A(n345), .B(n344), .Z(n528) );
  XOR2_X1 U335 ( .A(KEYINPUT28), .B(n474), .Z(n542) );
  XNOR2_X1 U336 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U337 ( .A(n489), .B(G43GAT), .ZN(n490) );
  XNOR2_X1 U338 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n491), .B(n490), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT81), .B(G134GAT), .Z(n292) );
  XNOR2_X1 U341 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U343 ( .A(G113GAT), .B(n293), .Z(n331) );
  XOR2_X1 U344 ( .A(KEYINPUT85), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U347 ( .A(G183GAT), .B(KEYINPUT86), .Z(n297) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U350 ( .A(n299), .B(n298), .Z(n313) );
  XOR2_X1 U351 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n301) );
  XNOR2_X1 U352 ( .A(KEYINPUT20), .B(KEYINPUT84), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n311) );
  XOR2_X1 U354 ( .A(G120GAT), .B(G71GAT), .Z(n416) );
  INV_X1 U355 ( .A(KEYINPUT19), .ZN(n302) );
  NAND2_X1 U356 ( .A1(KEYINPUT18), .A2(n302), .ZN(n305) );
  INV_X1 U357 ( .A(KEYINPUT18), .ZN(n303) );
  NAND2_X1 U358 ( .A1(n303), .A2(KEYINPUT19), .ZN(n304) );
  NAND2_X1 U359 ( .A1(n305), .A2(n304), .ZN(n307) );
  XNOR2_X1 U360 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n335) );
  XOR2_X1 U362 ( .A(n416), .B(n335), .Z(n309) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  INV_X1 U367 ( .A(n540), .ZN(n475) );
  XOR2_X1 U368 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n316) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(G148GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U371 ( .A(KEYINPUT4), .B(G57GAT), .Z(n318) );
  XNOR2_X1 U372 ( .A(KEYINPUT5), .B(KEYINPUT90), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U374 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U375 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n322) );
  NAND2_X1 U376 ( .A1(G225GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U378 ( .A(G1GAT), .B(n323), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n330) );
  XNOR2_X1 U380 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n326), .B(KEYINPUT2), .ZN(n451) );
  XOR2_X1 U382 ( .A(G85GAT), .B(n451), .Z(n328) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(G162GAT), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U385 ( .A(n330), .B(n329), .Z(n333) );
  XNOR2_X1 U386 ( .A(G29GAT), .B(n331), .ZN(n332) );
  XOR2_X1 U387 ( .A(n333), .B(n332), .Z(n481) );
  XOR2_X1 U388 ( .A(G169GAT), .B(G8GAT), .Z(n395) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(G218GAT), .ZN(n336) );
  XOR2_X1 U390 ( .A(G183GAT), .B(KEYINPUT75), .Z(n361) );
  XNOR2_X1 U391 ( .A(n336), .B(n361), .ZN(n337) );
  XOR2_X1 U392 ( .A(n338), .B(n337), .Z(n342) );
  XNOR2_X1 U393 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n339), .B(G211GAT), .ZN(n447) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n340), .B(G64GAT), .ZN(n399) );
  XNOR2_X1 U397 ( .A(n447), .B(n399), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U399 ( .A(n395), .B(n343), .Z(n345) );
  NAND2_X1 U400 ( .A1(G226GAT), .A2(G233GAT), .ZN(n344) );
  INV_X1 U401 ( .A(n528), .ZN(n435) );
  XOR2_X1 U402 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n434) );
  XOR2_X1 U403 ( .A(G155GAT), .B(G211GAT), .Z(n347) );
  XNOR2_X1 U404 ( .A(G127GAT), .B(G71GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U406 ( .A(n348), .B(G78GAT), .Z(n351) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G1GAT), .Z(n396) );
  INV_X1 U408 ( .A(n396), .ZN(n349) );
  XOR2_X1 U409 ( .A(n349), .B(G22GAT), .Z(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n365) );
  XOR2_X1 U411 ( .A(G57GAT), .B(KEYINPUT13), .Z(n415) );
  XOR2_X1 U412 ( .A(n415), .B(KEYINPUT14), .Z(n353) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT76), .Z(n355) );
  XNOR2_X1 U416 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U418 ( .A(n357), .B(n356), .Z(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n359) );
  XNOR2_X1 U420 ( .A(G8GAT), .B(G64GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n591) );
  INV_X1 U425 ( .A(n591), .ZN(n575) );
  XOR2_X1 U426 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n367) );
  XNOR2_X1 U427 ( .A(KEYINPUT11), .B(KEYINPUT74), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U429 ( .A(G92GAT), .B(G106GAT), .Z(n369) );
  XNOR2_X1 U430 ( .A(G134GAT), .B(G190GAT), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U432 ( .A(n371), .B(n370), .Z(n373) );
  XOR2_X1 U433 ( .A(G218GAT), .B(G162GAT), .Z(n453) );
  XOR2_X1 U434 ( .A(G99GAT), .B(G85GAT), .Z(n398) );
  XNOR2_X1 U435 ( .A(n453), .B(n398), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U437 ( .A(KEYINPUT73), .B(KEYINPUT65), .Z(n375) );
  NAND2_X1 U438 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n384) );
  XOR2_X1 U441 ( .A(G43GAT), .B(G29GAT), .Z(n379) );
  XNOR2_X1 U442 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U444 ( .A(n380), .B(KEYINPUT68), .Z(n382) );
  XNOR2_X1 U445 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n391), .B(KEYINPUT64), .ZN(n383) );
  XOR2_X1 U448 ( .A(n384), .B(n383), .Z(n550) );
  INV_X1 U449 ( .A(n550), .ZN(n565) );
  XOR2_X1 U450 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n423) );
  XOR2_X1 U451 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n386) );
  NAND2_X1 U452 ( .A1(G229GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U454 ( .A(G141GAT), .B(G22GAT), .Z(n454) );
  XOR2_X1 U455 ( .A(n387), .B(n454), .Z(n393) );
  XOR2_X1 U456 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n389) );
  XNOR2_X1 U457 ( .A(G113GAT), .B(G197GAT), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U462 ( .A(n397), .B(n396), .Z(n582) );
  INV_X1 U463 ( .A(n582), .ZN(n421) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n403) );
  INV_X1 U465 ( .A(n403), .ZN(n401) );
  AND2_X1 U466 ( .A1(G230GAT), .A2(G233GAT), .ZN(n402) );
  INV_X1 U467 ( .A(n402), .ZN(n400) );
  NAND2_X1 U468 ( .A1(n401), .A2(n400), .ZN(n405) );
  NAND2_X1 U469 ( .A1(n403), .A2(n402), .ZN(n404) );
  NAND2_X1 U470 ( .A1(n405), .A2(n404), .ZN(n406) );
  XOR2_X1 U471 ( .A(n406), .B(KEYINPUT72), .Z(n414) );
  XOR2_X1 U472 ( .A(G78GAT), .B(G148GAT), .Z(n408) );
  XNOR2_X1 U473 ( .A(G106GAT), .B(G204GAT), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n448) );
  XNOR2_X1 U475 ( .A(n448), .B(KEYINPUT71), .ZN(n412) );
  XOR2_X1 U476 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n410) );
  XNOR2_X1 U477 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n409) );
  XOR2_X1 U478 ( .A(n410), .B(n409), .Z(n411) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n588) );
  XNOR2_X1 U481 ( .A(n588), .B(n419), .ZN(n558) );
  INV_X1 U482 ( .A(n558), .ZN(n420) );
  NAND2_X1 U483 ( .A1(n421), .A2(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  NAND2_X1 U485 ( .A1(n565), .A2(n424), .ZN(n425) );
  NOR2_X1 U486 ( .A1(n575), .A2(n425), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n426), .B(KEYINPUT47), .ZN(n432) );
  XOR2_X1 U488 ( .A(KEYINPUT36), .B(n550), .Z(n596) );
  NOR2_X1 U489 ( .A1(n596), .A2(n591), .ZN(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT45), .B(n427), .ZN(n428) );
  NAND2_X1 U491 ( .A1(n428), .A2(n588), .ZN(n429) );
  XOR2_X1 U492 ( .A(KEYINPUT110), .B(n429), .Z(n430) );
  XOR2_X1 U493 ( .A(KEYINPUT69), .B(n582), .Z(n465) );
  NAND2_X1 U494 ( .A1(n430), .A2(n465), .ZN(n431) );
  AND2_X1 U495 ( .A1(n432), .A2(n431), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n537) );
  NOR2_X1 U497 ( .A1(n435), .A2(n537), .ZN(n438) );
  INV_X1 U498 ( .A(n438), .ZN(n437) );
  INV_X1 U499 ( .A(KEYINPUT54), .ZN(n436) );
  NAND2_X1 U500 ( .A1(n437), .A2(n436), .ZN(n440) );
  NAND2_X1 U501 ( .A1(KEYINPUT54), .A2(n438), .ZN(n439) );
  NAND2_X1 U502 ( .A1(n440), .A2(n439), .ZN(n441) );
  AND2_X1 U503 ( .A1(n481), .A2(n441), .ZN(n580) );
  XOR2_X1 U504 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n443) );
  XNOR2_X1 U505 ( .A(G50GAT), .B(KEYINPUT89), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n458) );
  XOR2_X1 U507 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n445) );
  NAND2_X1 U508 ( .A1(G228GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U510 ( .A(n446), .B(KEYINPUT23), .Z(n450) );
  XNOR2_X1 U511 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U513 ( .A(n452), .B(n451), .Z(n456) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n474) );
  NAND2_X1 U517 ( .A1(n580), .A2(n474), .ZN(n459) );
  XOR2_X1 U518 ( .A(n459), .B(KEYINPUT55), .Z(n460) );
  NAND2_X1 U519 ( .A1(n576), .A2(n550), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n462) );
  INV_X1 U521 ( .A(n465), .ZN(n568) );
  NAND2_X1 U522 ( .A1(n568), .A2(n588), .ZN(n496) );
  AND2_X1 U523 ( .A1(n528), .A2(n540), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT95), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n467), .A2(n474), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n528), .B(KEYINPUT27), .ZN(n473) );
  NOR2_X1 U527 ( .A1(n540), .A2(n474), .ZN(n472) );
  XNOR2_X1 U528 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n579) );
  NAND2_X1 U530 ( .A1(n473), .A2(n579), .ZN(n477) );
  INV_X1 U531 ( .A(n481), .ZN(n524) );
  NAND2_X1 U532 ( .A1(n524), .A2(n473), .ZN(n538) );
  NOR2_X1 U533 ( .A1(n538), .A2(n542), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n476), .A2(n475), .ZN(n480) );
  AND2_X1 U535 ( .A1(n477), .A2(n480), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n484) );
  INV_X1 U537 ( .A(n480), .ZN(n482) );
  OR2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n483) );
  AND2_X1 U539 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U540 ( .A(KEYINPUT97), .B(n485), .Z(n494) );
  NAND2_X1 U541 ( .A1(n591), .A2(n494), .ZN(n486) );
  NOR2_X1 U542 ( .A1(n486), .A2(n596), .ZN(n487) );
  XNOR2_X1 U543 ( .A(n487), .B(KEYINPUT37), .ZN(n523) );
  NOR2_X1 U544 ( .A1(n496), .A2(n523), .ZN(n488) );
  XNOR2_X1 U545 ( .A(n488), .B(KEYINPUT38), .ZN(n510) );
  NAND2_X1 U546 ( .A1(n540), .A2(n510), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n489) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n498) );
  XOR2_X1 U549 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n493) );
  NAND2_X1 U550 ( .A1(n575), .A2(n565), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n495) );
  NAND2_X1 U552 ( .A1(n495), .A2(n494), .ZN(n512) );
  NOR2_X1 U553 ( .A1(n496), .A2(n512), .ZN(n504) );
  NAND2_X1 U554 ( .A1(n524), .A2(n504), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n498), .B(n497), .ZN(G1324GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n500) );
  NAND2_X1 U557 ( .A1(n504), .A2(n528), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U559 ( .A(G8GAT), .B(n501), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n503) );
  NAND2_X1 U561 ( .A1(n504), .A2(n540), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n542), .A2(n504), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n505), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U565 ( .A1(n524), .A2(n510), .ZN(n507) );
  XOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .Z(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NAND2_X1 U568 ( .A1(n510), .A2(n528), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n508), .B(KEYINPUT100), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n509), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n510), .A2(n542), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n511), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n515) );
  NAND2_X1 U574 ( .A1(n582), .A2(n420), .ZN(n522) );
  NOR2_X1 U575 ( .A1(n512), .A2(n522), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(KEYINPUT102), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n524), .A2(n519), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n519), .A2(n528), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT103), .Z(n518) );
  NAND2_X1 U582 ( .A1(n540), .A2(n519), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U585 ( .A1(n519), .A2(n542), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n526) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n533), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n533), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n531) );
  NAND2_X1 U595 ( .A1(n533), .A2(n540), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n532), .ZN(G1338GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U599 ( .A1(n533), .A2(n542), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U601 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  NOR2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT112), .ZN(n555) );
  NAND2_X1 U604 ( .A1(n540), .A2(n555), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n568), .A2(n551), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U609 ( .A1(n551), .A2(n420), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n549) );
  XOR2_X1 U612 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n547) );
  NAND2_X1 U613 ( .A1(n551), .A2(n575), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U619 ( .A(G134GAT), .B(n554), .Z(G1343GAT) );
  NAND2_X1 U620 ( .A1(n579), .A2(n555), .ZN(n564) );
  NOR2_X1 U621 ( .A1(n582), .A2(n564), .ZN(n556) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n556), .Z(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT116), .B(n557), .ZN(G1344GAT) );
  NOR2_X1 U624 ( .A1(n564), .A2(n558), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n591), .A2(n564), .ZN(n563) );
  XOR2_X1 U630 ( .A(G155GAT), .B(n563), .Z(G1346GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT118), .B(n566), .Z(n567) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n576), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n571) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT56), .B(n572), .Z(n574) );
  NAND2_X1 U640 ( .A1(n576), .A2(n420), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  XOR2_X1 U642 ( .A(G183GAT), .B(KEYINPUT121), .Z(n578) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1350GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT123), .B(n581), .Z(n595) );
  NOR2_X1 U647 ( .A1(n582), .A2(n595), .ZN(n587) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(KEYINPUT124), .B(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1352GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n595), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  NOR2_X1 U656 ( .A1(n591), .A2(n595), .ZN(n592) );
  XOR2_X1 U657 ( .A(G211GAT), .B(n592), .Z(G1354GAT) );
  XOR2_X1 U658 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n594) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n594), .B(n593), .ZN(n598) );
  NOR2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U662 ( .A(n598), .B(n597), .Z(G1355GAT) );
endmodule

