//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  OR3_X1    g0012(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT65), .ZN(new_n213));
  OAI21_X1  g0013(.A(KEYINPUT65), .B1(new_n211), .B2(new_n212), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G97), .A2(G257), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT66), .Z(new_n224));
  AOI211_X1 g0024(.A(new_n222), .B(new_n224), .C1(G87), .C2(G250), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(new_n214), .B2(new_n213), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n212), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n206), .A2(new_n207), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n218), .B(new_n228), .C1(new_n230), .C2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  INV_X1    g0035(.A(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  INV_X1    g0038(.A(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n245), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(new_n208), .A2(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT8), .A2(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT69), .B(G58), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(KEYINPUT8), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n251), .A2(KEYINPUT70), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G150), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n257), .B(new_n259), .C1(KEYINPUT70), .C2(new_n251), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n229), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n207), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n261), .B(new_n229), .C1(G1), .C2(new_n212), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(new_n207), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT68), .A2(G223), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT68), .A2(G223), .ZN(new_n273));
  OAI21_X1  g0073(.A(G1698), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n229), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n280), .B(new_n282), .C1(G77), .C2(new_n277), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n284), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n283), .B(new_n287), .C1(new_n236), .C2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n269), .A2(new_n270), .B1(G200), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT72), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n271), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n271), .A2(new_n292), .A3(KEYINPUT10), .A4(new_n295), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n291), .A2(G179), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n300), .B(KEYINPUT71), .Z(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n269), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n298), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n277), .A2(G232), .A3(new_n278), .ZN(new_n306));
  INV_X1    g0106(.A(G107), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n277), .A2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(G238), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n306), .B1(new_n307), .B2(new_n277), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n286), .B1(new_n310), .B2(new_n282), .ZN(new_n311));
  INV_X1    g0111(.A(new_n290), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G244), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n302), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT15), .B(G87), .Z(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(new_n258), .B1(new_n318), .B2(new_n256), .ZN(new_n319));
  INV_X1    g0119(.A(G77), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n212), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n262), .B1(new_n320), .B2(new_n265), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n320), .B2(new_n267), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n311), .A2(new_n324), .A3(new_n313), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n315), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n314), .A2(G200), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n293), .B2(new_n314), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n328), .B2(new_n323), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n277), .B1(G232), .B2(new_n278), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G226), .A2(G1698), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n282), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n312), .A2(G238), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n287), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n336), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G179), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n334), .A2(KEYINPUT13), .A3(new_n287), .A4(new_n335), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(G169), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n342), .A2(new_n346), .A3(G169), .A4(new_n343), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n340), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n256), .A2(G77), .B1(new_n258), .B2(G50), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n212), .B2(G68), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(KEYINPUT11), .A3(new_n262), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n203), .B2(new_n267), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n264), .A2(G68), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT11), .B1(new_n350), .B2(new_n262), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n339), .A2(G190), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n342), .A2(G200), .A3(new_n343), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n277), .A2(G223), .A3(new_n278), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n308), .B2(new_n236), .ZN(new_n364));
  INV_X1    g0164(.A(G87), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n255), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n282), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n312), .A2(G232), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n287), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n302), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n367), .A2(new_n324), .A3(new_n287), .A4(new_n368), .ZN(new_n371));
  INV_X1    g0171(.A(new_n262), .ZN(new_n372));
  AND2_X1   g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  NOR2_X1   g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n375), .B2(new_n212), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NOR4_X1   g0177(.A1(new_n373), .A2(new_n374), .A3(new_n377), .A4(G20), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n258), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT69), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G58), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(G68), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(new_n204), .A3(new_n205), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n380), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT16), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n275), .A2(new_n212), .A3(new_n276), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n377), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n276), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(G68), .B1(G20), .B2(new_n385), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n380), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n372), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n254), .A2(new_n267), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n254), .B2(new_n265), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n397), .B(KEYINPUT74), .C1(new_n254), .C2(new_n265), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n370), .B(new_n371), .C1(new_n396), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n394), .B1(new_n393), .B2(new_n380), .ZN(new_n407));
  AND4_X1   g0207(.A1(new_n394), .A2(new_n379), .A3(new_n380), .A4(new_n386), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n262), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n402), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .A3(new_n370), .A4(new_n371), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT75), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n396), .A2(new_n403), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n369), .A2(G200), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n367), .A2(G190), .A3(new_n287), .A4(new_n368), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n409), .A2(new_n416), .A3(new_n417), .A4(new_n402), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n404), .A2(KEYINPUT75), .A3(new_n405), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n413), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NOR4_X1   g0223(.A1(new_n305), .A2(new_n329), .A3(new_n362), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n211), .A2(G45), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(new_n285), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(G250), .C1(new_n281), .C2(new_n229), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT77), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n289), .A2(new_n429), .A3(G250), .A4(new_n425), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(G244), .B(G1698), .C1(new_n373), .C2(new_n374), .ZN(new_n432));
  OAI211_X1 g0232(.A(G238), .B(new_n278), .C1(new_n373), .C2(new_n374), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G116), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n282), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(new_n436), .A3(G190), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT78), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n436), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT78), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n431), .A2(new_n436), .A3(new_n441), .A4(G190), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT19), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n212), .B1(new_n330), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G97), .A2(G107), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n365), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n212), .B(G68), .C1(new_n373), .C2(new_n374), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n444), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n262), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n318), .A2(new_n264), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n211), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n264), .A2(new_n456), .A3(new_n229), .A4(new_n261), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n365), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n443), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n439), .A2(new_n302), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n454), .B1(new_n452), .B2(new_n262), .ZN(new_n463));
  INV_X1    g0263(.A(new_n318), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n431), .A2(new_n436), .A3(new_n324), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT25), .ZN(new_n470));
  AOI211_X1 g0270(.A(G107), .B(new_n264), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n469), .A2(new_n470), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n473), .A2(new_n474), .B1(new_n307), .B2(new_n457), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n212), .B(G87), .C1(new_n373), .C2(new_n374), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT22), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n277), .A2(new_n478), .A3(new_n212), .A4(G87), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n434), .A2(G20), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n212), .A2(G107), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT23), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT80), .B(KEYINPUT24), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n481), .B1(new_n477), .B2(new_n479), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n486), .A3(new_n484), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n475), .B1(new_n491), .B2(new_n262), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n277), .A2(G257), .A3(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G294), .ZN(new_n494));
  OAI211_X1 g0294(.A(G250), .B(new_n278), .C1(new_n373), .C2(new_n374), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n282), .ZN(new_n497));
  INV_X1    g0297(.A(new_n425), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n282), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G264), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(G274), .A3(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G169), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n496), .A2(new_n282), .B1(G264), .B2(new_n500), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G179), .A3(new_n502), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(KEYINPUT82), .A3(new_n506), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n492), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n468), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n265), .A2(new_n248), .ZN(new_n513));
  INV_X1    g0313(.A(new_n457), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G116), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n212), .B1(new_n516), .B2(G33), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT76), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT76), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(G33), .A3(G283), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n262), .B1(new_n212), .B2(G116), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT20), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n520), .B1(G33), .B2(G283), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n518), .A2(KEYINPUT76), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n261), .A2(new_n229), .B1(G20), .B2(new_n248), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT20), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n513), .B(new_n515), .C1(new_n525), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n278), .A2(G257), .ZN(new_n533));
  OAI221_X1 g0333(.A(new_n533), .B1(new_n239), .B2(new_n278), .C1(new_n373), .C2(new_n374), .ZN(new_n534));
  INV_X1    g0334(.A(G303), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n275), .A2(new_n535), .A3(new_n276), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n282), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n499), .A2(new_n498), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(G270), .A3(new_n289), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n539), .A3(new_n502), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n532), .A2(G169), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n537), .A2(new_n502), .A3(new_n539), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n532), .A2(G179), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(G190), .ZN(new_n546));
  INV_X1    g0346(.A(new_n513), .ZN(new_n547));
  INV_X1    g0347(.A(new_n531), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n540), .A2(G200), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n546), .A2(new_n550), .A3(new_n515), .A4(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n532), .A2(KEYINPUT21), .A3(G169), .A4(new_n540), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n543), .A2(new_n545), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT79), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n392), .A2(G107), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n258), .A2(G77), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n307), .A2(KEYINPUT6), .A3(G97), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n516), .A2(new_n307), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n446), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n561), .B2(KEYINPUT6), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G20), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n262), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n265), .A2(new_n516), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n514), .A2(G97), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n538), .A2(G257), .A3(new_n289), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(new_n278), .C1(new_n373), .C2(new_n374), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .A4(new_n278), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n519), .A2(new_n521), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n569), .B1(new_n576), .B2(new_n282), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n302), .B1(new_n577), .B2(new_n502), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n282), .ZN(new_n579));
  INV_X1    g0379(.A(new_n569), .ZN(new_n580));
  AND4_X1   g0380(.A1(G179), .A2(new_n579), .A3(new_n502), .A4(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n568), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n502), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n564), .A2(new_n262), .B1(new_n516), .B2(new_n265), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n577), .A2(G190), .A3(new_n502), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n567), .A4(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n489), .A2(new_n486), .A3(new_n484), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n486), .B1(new_n489), .B2(new_n484), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n262), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n475), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n503), .A2(G200), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n505), .A2(G190), .A3(new_n502), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n582), .A2(new_n587), .A3(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n424), .A2(new_n512), .A3(new_n556), .A4(new_n595), .ZN(G372));
  NAND2_X1  g0396(.A1(new_n406), .A2(new_n411), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n326), .A2(KEYINPUT89), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n326), .A2(KEYINPUT89), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n361), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n358), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n598), .B1(new_n603), .B2(new_n421), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n298), .A2(new_n299), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n304), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT88), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT83), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n460), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n463), .A2(KEYINPUT83), .A3(new_n459), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n467), .B1(new_n443), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT84), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(KEYINPUT84), .B(new_n467), .C1(new_n443), .C2(new_n612), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n568), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT87), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n581), .B2(new_n578), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n579), .A2(G179), .A3(new_n502), .A4(new_n580), .ZN(new_n621));
  INV_X1    g0421(.A(new_n502), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n622), .B(new_n569), .C1(new_n576), .C2(new_n282), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(KEYINPUT87), .C1(new_n623), .C2(new_n302), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n618), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n608), .B(KEYINPUT26), .C1(new_n617), .C2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n445), .A2(new_n447), .B1(new_n444), .B2(new_n450), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n372), .B1(new_n627), .B2(new_n449), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n628), .A2(new_n609), .A3(new_n454), .A4(new_n458), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT83), .B1(new_n463), .B2(new_n459), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n440), .A3(new_n438), .A4(new_n442), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT84), .B1(new_n632), .B2(new_n467), .ZN(new_n633));
  INV_X1    g0433(.A(new_n616), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n625), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT88), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n468), .A2(new_n636), .A3(new_n582), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n626), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n582), .A2(new_n594), .A3(new_n587), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n615), .B2(new_n616), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n505), .A2(G179), .A3(new_n502), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n302), .B1(new_n505), .B2(new_n502), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT85), .B1(new_n492), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n543), .A2(new_n545), .A3(new_n553), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n590), .A2(new_n591), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT85), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n507), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n640), .B1(new_n642), .B2(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n640), .A2(new_n651), .A3(new_n617), .A4(new_n595), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n467), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n424), .B1(new_n639), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n607), .A2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(new_n556), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT91), .ZN(new_n658));
  INV_X1    g0458(.A(G13), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G20), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n211), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT90), .Z(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(G213), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n532), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n657), .A2(KEYINPUT91), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n658), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n647), .B2(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n511), .ZN(new_n673));
  INV_X1    g0473(.A(new_n667), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n673), .B(new_n594), .C1(new_n492), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n511), .A2(new_n667), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n647), .A2(new_n667), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n667), .B1(new_n646), .B2(new_n650), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n216), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n447), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n231), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n635), .A2(new_n636), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n608), .ZN(new_n696));
  INV_X1    g0496(.A(new_n638), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n635), .A2(KEYINPUT88), .A3(new_n636), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n467), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n651), .A2(new_n617), .A3(new_n595), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT86), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n642), .A2(new_n640), .A3(new_n651), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n667), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT93), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n674), .B1(new_n639), .B2(new_n654), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT93), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n582), .A2(new_n587), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT95), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n673), .A2(new_n647), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n594), .A3(new_n617), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n635), .A2(KEYINPUT26), .ZN(new_n717));
  OR3_X1    g0517(.A1(new_n468), .A2(KEYINPUT26), .A3(new_n582), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n467), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n717), .A2(new_n721), .A3(new_n718), .A4(new_n467), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n716), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .A3(new_n674), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n577), .A2(new_n505), .A3(new_n502), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n544), .A2(G179), .A3(new_n436), .A4(new_n431), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT92), .ZN(new_n729));
  OR3_X1    g0529(.A1(new_n726), .A2(new_n727), .A3(new_n725), .ZN(new_n730));
  AOI21_X1  g0530(.A(G179), .B1(new_n431), .B2(new_n436), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n583), .A2(new_n503), .A3(new_n540), .A4(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT92), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n733), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n729), .A2(new_n730), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n735), .A2(new_n667), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n556), .A2(new_n512), .A3(new_n595), .A4(new_n674), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(KEYINPUT31), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n730), .A2(new_n732), .A3(new_n728), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n711), .A2(new_n724), .B1(G330), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n694), .B1(new_n742), .B2(G1), .ZN(G364));
  AOI21_X1  g0543(.A(new_n211), .B1(new_n660), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n688), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n671), .B2(G330), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n671), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n212), .A2(new_n324), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G190), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n375), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(G20), .A3(new_n324), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n753), .B1(G329), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G294), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n212), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n324), .A2(G200), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n756), .B1(new_n757), .B2(new_n759), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT97), .ZN(new_n767));
  INV_X1    g0567(.A(new_n749), .ZN(new_n768));
  INV_X1    g0568(.A(G200), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n749), .A2(KEYINPUT97), .A3(G200), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n293), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n766), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n749), .A2(G190), .A3(new_n769), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G322), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n762), .A2(new_n293), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G303), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(G190), .A3(new_n771), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G326), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n775), .A2(new_n778), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n783), .A2(G87), .ZN(new_n789));
  INV_X1    g0589(.A(new_n785), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G50), .A2(new_n790), .B1(new_n773), .B2(G68), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n764), .A2(new_n307), .ZN(new_n792));
  INV_X1    g0592(.A(new_n253), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n277), .B1(new_n793), .B2(new_n776), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n759), .A2(new_n516), .B1(new_n751), .B2(new_n320), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n789), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n755), .A2(G159), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT32), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n788), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT101), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n229), .B1(G20), .B2(new_n302), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n245), .A2(G45), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n687), .A2(new_n277), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(G45), .C2(new_n692), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n216), .A2(G355), .A3(new_n277), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(G116), .C2(new_n216), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT96), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n811), .B(new_n802), .C1(new_n807), .C2(KEYINPUT96), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n801), .A2(new_n802), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n811), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n746), .B(new_n813), .C1(new_n671), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n748), .A2(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n667), .A2(new_n323), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n599), .A2(new_n600), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n329), .A2(new_n817), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n822), .A2(G330), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n741), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n822), .B1(new_n741), .B2(G330), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n826), .A2(new_n705), .ZN(new_n827));
  INV_X1    g0627(.A(new_n746), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n705), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n764), .A2(new_n203), .B1(new_n793), .B2(new_n759), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n375), .B1(new_n755), .B2(G132), .ZN(new_n832));
  INV_X1    g0632(.A(new_n751), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n790), .A2(G137), .B1(G159), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n776), .C1(new_n836), .C2(new_n772), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT34), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n832), .B1(new_n207), .B2(new_n782), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n831), .B(new_n839), .C1(new_n838), .C2(new_n837), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n375), .B1(new_n757), .B2(new_n776), .C1(new_n782), .C2(new_n307), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n763), .A2(G87), .B1(G311), .B2(new_n755), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT103), .Z(new_n843));
  OAI22_X1  g0643(.A1(new_n772), .A2(new_n765), .B1(new_n248), .B2(new_n751), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT102), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n785), .A2(new_n535), .B1(new_n516), .B2(new_n759), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n841), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n802), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n822), .B2(new_n810), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n802), .A2(new_n809), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n320), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n830), .B1(new_n828), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT104), .ZN(G384));
  INV_X1    g0653(.A(KEYINPUT40), .ZN(new_n854));
  INV_X1    g0654(.A(new_n665), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n396), .B2(new_n403), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n423), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n856), .B2(KEYINPUT105), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n404), .A2(new_n419), .A3(new_n856), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n858), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n358), .B(new_n361), .C1(new_n356), .C2(new_n674), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n357), .B(new_n667), .C1(new_n602), .C2(new_n348), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n821), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT108), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n869), .B1(new_n738), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n854), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n738), .A2(new_n872), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n861), .B(new_n859), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n856), .B1(new_n597), .B2(new_n421), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n863), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n875), .A2(KEYINPUT40), .A3(new_n880), .A4(new_n869), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n875), .A2(new_n424), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(G330), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n711), .A2(new_n886), .A3(new_n424), .A4(new_n724), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n706), .A2(new_n710), .A3(new_n424), .A4(new_n724), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT107), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n607), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n885), .B(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n858), .A2(new_n862), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n876), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n895), .B2(new_n863), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n863), .A2(new_n893), .A3(new_n879), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT106), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n864), .B2(new_n865), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n863), .A2(new_n879), .A3(new_n893), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n358), .A2(new_n667), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n898), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n598), .A2(new_n665), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n867), .A2(new_n868), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n674), .B(new_n822), .C1(new_n639), .C2(new_n654), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n326), .A2(new_n667), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n907), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n895), .A2(new_n863), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n904), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n892), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n211), .B2(new_n660), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n248), .B1(new_n562), .B2(KEYINPUT35), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n230), .C1(KEYINPUT35), .C2(new_n562), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n231), .A2(G77), .A3(new_n384), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(G50), .B2(new_n203), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n659), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n920), .A3(new_n923), .ZN(G367));
  INV_X1    g0724(.A(KEYINPUT46), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n782), .B2(new_n248), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT112), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n782), .A2(new_n925), .A3(new_n248), .ZN(new_n928));
  INV_X1    g0728(.A(new_n786), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n752), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n772), .A2(new_n757), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n763), .A2(G97), .ZN(new_n932));
  INV_X1    g0732(.A(new_n759), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G107), .ZN(new_n934));
  XNOR2_X1  g0734(.A(KEYINPUT113), .B(G317), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n277), .B1(new_n755), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n777), .A2(G303), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n932), .A2(new_n934), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  NOR4_X1   g0738(.A1(new_n928), .A2(new_n930), .A3(new_n931), .A4(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n927), .B(new_n939), .C1(new_n765), .C2(new_n751), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT114), .Z(new_n941));
  NAND2_X1  g0741(.A1(new_n783), .A2(new_n253), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n759), .A2(new_n203), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n277), .B1(new_n751), .B2(new_n207), .C1(new_n836), .C2(new_n776), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(G137), .C2(new_n755), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n786), .A2(G143), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n764), .A2(new_n320), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G159), .B2(new_n773), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n942), .A2(new_n945), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT47), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n828), .B1(new_n951), .B2(new_n802), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n811), .A2(new_n802), .ZN(new_n953));
  INV_X1    g0753(.A(new_n804), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n953), .B1(new_n216), .B2(new_n464), .C1(new_n954), .C2(new_n241), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n667), .A2(new_n612), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n467), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n617), .B2(new_n956), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n952), .B(new_n955), .C1(new_n814), .C2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n674), .A2(new_n618), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n713), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n625), .A2(new_n667), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n683), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT42), .Z(new_n966));
  NOR2_X1   g0766(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n967));
  INV_X1    g0767(.A(new_n964), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n582), .B1(new_n968), .B2(new_n673), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n674), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT109), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n967), .B1(new_n966), .B2(new_n970), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n958), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n680), .B2(new_n968), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n973), .A2(new_n679), .A3(new_n964), .A4(new_n976), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n964), .A2(new_n685), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT44), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n964), .A2(new_n685), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n964), .B2(new_n685), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n679), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT111), .ZN(new_n990));
  INV_X1    g0790(.A(new_n683), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n677), .B2(new_n681), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n672), .B(new_n992), .Z(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n742), .A3(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n983), .A2(new_n987), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n680), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT111), .B1(new_n996), .B2(new_n989), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n742), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n688), .B(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n745), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n960), .B1(new_n980), .B2(new_n1002), .ZN(G387));
  OR2_X1    g0803(.A1(new_n742), .A2(new_n993), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n742), .A2(new_n993), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n688), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n802), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n773), .A2(G311), .B1(new_n777), .B2(new_n935), .ZN(new_n1008));
  INV_X1    g0808(.A(G322), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(new_n535), .B2(new_n751), .C1(new_n929), .C2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n765), .B2(new_n759), .C1(new_n757), .C2(new_n782), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT49), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n755), .A2(G326), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n277), .B1(new_n763), .B2(G116), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n464), .A2(new_n759), .ZN(new_n1019));
  INV_X1    g0819(.A(G159), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n254), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1020), .A2(new_n785), .B1(new_n772), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1019), .B(new_n1022), .C1(G97), .C2(new_n763), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n277), .B1(new_n754), .B2(new_n836), .C1(new_n776), .C2(new_n207), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G68), .B2(new_n833), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n320), .C2(new_n782), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1007), .B1(new_n1018), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n677), .A2(new_n814), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n690), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n216), .A2(new_n277), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G45), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n237), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n316), .A2(G50), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT115), .ZN(new_n1035));
  AOI21_X1  g0835(.A(G45), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(new_n1035), .C2(new_n1029), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n203), .A2(new_n320), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n804), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1030), .B1(G107), .B2(new_n216), .C1(new_n1032), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(new_n953), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1027), .A2(new_n828), .A3(new_n1028), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n993), .B2(new_n745), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1006), .A2(new_n1043), .ZN(G393));
  NAND3_X1  g0844(.A1(new_n989), .A2(new_n745), .A3(new_n996), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n953), .B1(new_n516), .B2(new_n216), .C1(new_n954), .C2(new_n249), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n783), .A2(G68), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G87), .A2(new_n763), .B1(new_n773), .B2(G50), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n277), .B1(new_n754), .B2(new_n835), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n759), .A2(new_n320), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n317), .C2(new_n833), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n785), .A2(new_n836), .B1(new_n1020), .B2(new_n776), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n375), .B1(new_n1009), .B2(new_n754), .C1(new_n759), .C2(new_n248), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1055), .B(new_n792), .C1(G303), .C2(new_n773), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n790), .A2(G317), .B1(G311), .B2(new_n777), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(new_n765), .C2(new_n782), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n751), .A2(new_n757), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1054), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n828), .B1(new_n1061), .B2(new_n802), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1046), .B(new_n1062), .C1(new_n964), .C2(new_n814), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n688), .B1(new_n994), .B2(new_n997), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n993), .A2(new_n742), .B1(new_n989), .B2(new_n996), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1045), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(G390));
  OAI21_X1  g0866(.A(KEYINPUT116), .B1(new_n911), .B2(new_n903), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n898), .A2(new_n902), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT116), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n903), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n909), .B1(new_n705), .B2(new_n822), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1070), .C1(new_n1071), .C2(new_n907), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n723), .A2(new_n674), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n909), .B1(new_n1074), .B2(new_n822), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1070), .B(new_n880), .C1(new_n1075), .C2(new_n907), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n824), .A2(new_n906), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1073), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n875), .A2(new_n823), .A3(new_n906), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1079), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n745), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1068), .A2(new_n809), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n790), .A2(G128), .ZN(new_n1086));
  INV_X1    g0886(.A(G132), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n277), .B1(new_n776), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G159), .B2(new_n933), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1086), .B(new_n1089), .C1(new_n764), .C2(new_n207), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n783), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT53), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n782), .B2(new_n836), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1090), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  AOI22_X1  g0895(.A1(new_n773), .A2(G137), .B1(new_n833), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT117), .ZN(new_n1097));
  INV_X1    g0897(.A(G125), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1094), .B(new_n1097), .C1(new_n1098), .C2(new_n754), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n375), .B1(new_n754), .B2(new_n757), .C1(new_n776), .C2(new_n248), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G97), .B2(new_n833), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n764), .B2(new_n203), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G107), .A2(new_n773), .B1(new_n790), .B2(G283), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n789), .B(new_n1103), .C1(new_n320), .C2(new_n759), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1099), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1105), .A2(new_n802), .B1(new_n1021), .B2(new_n850), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1085), .A2(new_n746), .A3(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1073), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1082), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n875), .A2(new_n823), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1075), .B(new_n1077), .C1(new_n906), .C2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1081), .B1(new_n824), .B2(new_n906), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1071), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n883), .A2(G330), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n890), .A2(new_n1116), .A3(new_n607), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n688), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n888), .A2(KEYINPUT107), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n888), .A2(KEYINPUT107), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n607), .B(new_n1117), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1083), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1084), .B(new_n1107), .C1(new_n1119), .C2(new_n1125), .ZN(G378));
  NAND2_X1  g0926(.A1(new_n783), .A2(new_n1095), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT118), .Z(new_n1128));
  NAND2_X1  g0928(.A1(new_n833), .A2(G137), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n785), .A2(new_n1098), .B1(new_n836), .B2(new_n759), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT119), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n773), .A2(G132), .B1(G128), .B2(new_n777), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1136));
  AOI21_X1  g0936(.A(G33), .B1(new_n755), .B2(G124), .ZN(new_n1137));
  AOI21_X1  g0937(.A(G41), .B1(new_n763), .B2(G159), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n207), .B1(new_n373), .B2(G41), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n763), .A2(new_n253), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n776), .A2(new_n307), .B1(new_n765), .B2(new_n754), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n318), .B2(new_n833), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n943), .A2(G41), .A3(new_n277), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G97), .B2(new_n773), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n320), .B2(new_n782), .C1(new_n248), .C2(new_n785), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT58), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1139), .A2(new_n1140), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n828), .B1(new_n1149), .B2(new_n802), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n305), .A2(KEYINPUT121), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT121), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n298), .A2(new_n1152), .A3(new_n299), .A4(new_n304), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n269), .A2(new_n855), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1155), .B(new_n1156), .Z(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1154), .B(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n809), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n850), .A2(new_n207), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1150), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n873), .B1(new_n895), .B2(new_n863), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G330), .B(new_n881), .C1(new_n1164), .C2(KEYINPUT40), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n874), .A2(new_n1159), .A3(G330), .A4(new_n881), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n915), .A2(new_n1169), .A3(KEYINPUT122), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n914), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(KEYINPUT122), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1163), .B1(new_n1172), .B2(new_n745), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1117), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n606), .B(new_n1174), .C1(new_n887), .C2(new_n889), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n1116), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1122), .A2(KEYINPUT123), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT123), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n890), .A2(new_n1178), .A3(new_n607), .A4(new_n1117), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT57), .B1(new_n1181), .B2(new_n1172), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1083), .A2(new_n1124), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n915), .A2(new_n1169), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n914), .B1(new_n1168), .B2(new_n1167), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n688), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1173), .B1(new_n1182), .B2(new_n1187), .ZN(G375));
  NAND2_X1  g0988(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n1118), .A3(new_n1001), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT124), .Z(new_n1191));
  NAND2_X1  g0991(.A1(new_n907), .A2(new_n809), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n375), .B1(new_n754), .B2(new_n535), .C1(new_n751), .C2(new_n307), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1193), .B(new_n947), .C1(G283), .C2(new_n777), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n248), .A2(new_n772), .B1(new_n785), .B2(new_n757), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n1019), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(new_n516), .C2(new_n782), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1141), .A2(new_n277), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT125), .Z(new_n1199));
  AOI22_X1  g0999(.A1(new_n777), .A2(G137), .B1(G128), .B2(new_n755), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n207), .B2(new_n759), .C1(new_n785), .C2(new_n1087), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n773), .B2(new_n1095), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1199), .B(new_n1202), .C1(new_n1020), .C2(new_n782), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n751), .A2(new_n836), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1197), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1205), .A2(new_n802), .B1(new_n203), .B2(new_n850), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1192), .A2(new_n746), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1116), .B2(new_n745), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1191), .A2(new_n1208), .ZN(G381));
  NOR3_X1   g1009(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1210));
  INV_X1    g1010(.A(G378), .ZN(new_n1211));
  INV_X1    g1011(.A(G375), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(G407));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n666), .A3(new_n1211), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(G407), .A2(G213), .A3(new_n1215), .ZN(G409));
  NAND3_X1  g1016(.A1(new_n1181), .A2(new_n1001), .A3(new_n1172), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n745), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1162), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1211), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G378), .B(new_n1173), .C1(new_n1182), .C2(new_n1187), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n666), .A2(G213), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n689), .B1(new_n1189), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1122), .A2(KEYINPUT60), .A3(new_n1123), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1118), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1208), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(G384), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT104), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n852), .B(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1227), .A3(new_n1208), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1222), .A2(new_n1223), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n666), .A2(G213), .A3(G2897), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1232), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1231), .B1(new_n1208), .B2(new_n1227), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1229), .A2(new_n1232), .A3(new_n1237), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1236), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT61), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1222), .A2(new_n1246), .A3(new_n1233), .A4(new_n1223), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1235), .A2(new_n1244), .A3(new_n1245), .A4(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G387), .A2(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(G393), .B(G396), .Z(new_n1251));
  OAI211_X1 g1051(.A(new_n960), .B(G390), .C1(new_n980), .C2(new_n1002), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1248), .A2(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1222), .A2(new_n1223), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT63), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1234), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1222), .A2(KEYINPUT63), .A3(new_n1233), .A4(new_n1223), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1255), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1262), .A3(new_n1245), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(G405));
  NOR2_X1   g1064(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT127), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT127), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1233), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G375), .A2(new_n1211), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1221), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1221), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(KEYINPUT127), .C1(new_n1266), .C2(new_n1265), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1271), .A2(new_n1255), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1255), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G402));
endmodule


