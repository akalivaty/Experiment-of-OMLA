

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744;

  NAND2_X1 U375 ( .A1(n510), .A2(n683), .ZN(n680) );
  XNOR2_X1 U376 ( .A(n432), .B(KEYINPUT4), .ZN(n477) );
  AND2_X2 U377 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U378 ( .A(G119), .B(G116), .ZN(n435) );
  INV_X1 U379 ( .A(G953), .ZN(n728) );
  AND2_X2 U380 ( .A1(n714), .A2(n362), .ZN(n371) );
  XNOR2_X2 U381 ( .A(n517), .B(KEYINPUT1), .ZN(n556) );
  XNOR2_X1 U382 ( .A(n479), .B(G134), .ZN(n454) );
  XNOR2_X1 U383 ( .A(n401), .B(G110), .ZN(n478) );
  XNOR2_X2 U384 ( .A(n398), .B(n557), .ZN(n582) );
  NOR2_X2 U385 ( .A1(n556), .A2(n680), .ZN(n398) );
  XNOR2_X2 U386 ( .A(n366), .B(n367), .ZN(n597) );
  NOR2_X2 U387 ( .A1(n589), .A2(n571), .ZN(n366) );
  NOR2_X1 U388 ( .A1(n492), .A2(n395), .ZN(n394) );
  INV_X1 U389 ( .A(G146), .ZN(n401) );
  INV_X1 U390 ( .A(KEYINPUT73), .ZN(n557) );
  NAND2_X1 U391 ( .A1(n606), .A2(KEYINPUT44), .ZN(n385) );
  INV_X1 U392 ( .A(KEYINPUT83), .ZN(n569) );
  AND2_X1 U393 ( .A1(n545), .A2(n546), .ZN(n384) );
  INV_X1 U394 ( .A(KEYINPUT66), .ZN(n432) );
  INV_X1 U395 ( .A(G128), .ZN(n430) );
  NOR2_X1 U396 ( .A1(n531), .A2(n509), .ZN(n388) );
  NAND2_X2 U397 ( .A1(n376), .A2(n374), .ZN(n517) );
  OR2_X1 U398 ( .A1(n368), .A2(n375), .ZN(n374) );
  NAND2_X1 U399 ( .A1(n379), .A2(G902), .ZN(n377) );
  XNOR2_X1 U400 ( .A(n726), .B(n442), .ZN(n633) );
  XNOR2_X1 U401 ( .A(n725), .B(n409), .ZN(n412) );
  XNOR2_X1 U402 ( .A(G119), .B(G137), .ZN(n402) );
  XNOR2_X1 U403 ( .A(G146), .B(KEYINPUT67), .ZN(n433) );
  NOR2_X1 U404 ( .A1(n548), .A2(n553), .ZN(n497) );
  BUF_X1 U405 ( .A(n556), .Z(n681) );
  XNOR2_X1 U406 ( .A(n392), .B(n537), .ZN(n544) );
  AND2_X1 U407 ( .A1(n445), .A2(n596), .ZN(n446) );
  NAND2_X1 U408 ( .A1(n503), .A2(n475), .ZN(n375) );
  AND2_X1 U409 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U410 ( .A1(n383), .A2(n381), .ZN(n727) );
  XNOR2_X1 U411 ( .A(n384), .B(KEYINPUT48), .ZN(n383) );
  INV_X1 U412 ( .A(n669), .ZN(n382) );
  INV_X1 U413 ( .A(G122), .ZN(n449) );
  XOR2_X1 U414 ( .A(G143), .B(G122), .Z(n464) );
  NAND2_X1 U415 ( .A1(n371), .A2(n372), .ZN(n370) );
  XNOR2_X1 U416 ( .A(n727), .B(n373), .ZN(n372) );
  INV_X1 U417 ( .A(KEYINPUT74), .ZN(n373) );
  XNOR2_X1 U418 ( .A(G107), .B(G101), .ZN(n498) );
  XOR2_X1 U419 ( .A(G110), .B(G104), .Z(n499) );
  XNOR2_X1 U420 ( .A(n454), .B(n477), .ZN(n380) );
  INV_X1 U421 ( .A(KEYINPUT33), .ZN(n396) );
  NOR2_X1 U422 ( .A1(n389), .A2(n387), .ZN(n530) );
  XNOR2_X1 U423 ( .A(n414), .B(n413), .ZN(n644) );
  XNOR2_X1 U424 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U425 ( .A(n393), .B(KEYINPUT40), .ZN(n743) );
  OR2_X1 U426 ( .A1(n547), .A2(n663), .ZN(n393) );
  XNOR2_X1 U427 ( .A(n505), .B(KEYINPUT111), .ZN(n742) );
  XNOR2_X1 U428 ( .A(n586), .B(n585), .ZN(n667) );
  INV_X1 U429 ( .A(KEYINPUT92), .ZN(n583) );
  XOR2_X1 U430 ( .A(n502), .B(n501), .Z(n356) );
  OR2_X1 U431 ( .A1(n522), .A2(n655), .ZN(n357) );
  XOR2_X1 U432 ( .A(n520), .B(n519), .Z(n358) );
  NOR2_X1 U433 ( .A1(n596), .A2(n595), .ZN(n359) );
  AND2_X1 U434 ( .A1(n390), .A2(n391), .ZN(n360) );
  XNOR2_X1 U435 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n361) );
  NOR2_X1 U436 ( .A1(n492), .A2(KEYINPUT2), .ZN(n362) );
  XOR2_X1 U437 ( .A(n709), .B(n708), .Z(n363) );
  INV_X1 U438 ( .A(KEYINPUT2), .ZN(n395) );
  NAND2_X1 U439 ( .A1(n370), .A2(n369), .ZN(n364) );
  NAND2_X1 U440 ( .A1(n370), .A2(n369), .ZN(n365) );
  NAND2_X1 U441 ( .A1(n670), .A2(n394), .ZN(n369) );
  NAND2_X1 U442 ( .A1(n370), .A2(n369), .ZN(n707) );
  XOR2_X1 U443 ( .A(KEYINPUT71), .B(KEYINPUT22), .Z(n367) );
  OR2_X2 U444 ( .A1(n623), .A2(n625), .ZN(n607) );
  OR2_X1 U445 ( .A1(n627), .A2(n615), .ZN(n495) );
  NAND2_X1 U446 ( .A1(n368), .A2(n379), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n368), .B(n363), .ZN(n710) );
  XNOR2_X2 U448 ( .A(n726), .B(n356), .ZN(n368) );
  NAND2_X1 U449 ( .A1(n714), .A2(n614), .ZN(n670) );
  XNOR2_X2 U450 ( .A(n613), .B(KEYINPUT45), .ZN(n714) );
  INV_X1 U451 ( .A(n503), .ZN(n379) );
  AND2_X2 U452 ( .A1(n575), .A2(n574), .ZN(n623) );
  NAND2_X1 U453 ( .A1(n567), .A2(n566), .ZN(n386) );
  NOR2_X2 U454 ( .A1(n700), .A2(n589), .ZN(n564) );
  XNOR2_X2 U455 ( .A(n563), .B(KEYINPUT0), .ZN(n589) );
  XNOR2_X2 U456 ( .A(n380), .B(n434), .ZN(n726) );
  XNOR2_X2 U457 ( .A(n431), .B(n430), .ZN(n479) );
  AND2_X1 U458 ( .A1(n737), .A2(n382), .ZN(n381) );
  XNOR2_X1 U459 ( .A(n385), .B(n569), .ZN(n603) );
  XNOR2_X2 U460 ( .A(n386), .B(n568), .ZN(n606) );
  XNOR2_X1 U461 ( .A(n508), .B(n361), .ZN(n390) );
  NAND2_X1 U462 ( .A1(n360), .A2(n588), .ZN(n528) );
  NAND2_X1 U463 ( .A1(n390), .A2(n388), .ZN(n387) );
  INV_X1 U464 ( .A(n588), .ZN(n389) );
  INV_X1 U465 ( .A(n509), .ZN(n391) );
  NAND2_X1 U466 ( .A1(n743), .A2(n744), .ZN(n392) );
  XNOR2_X2 U467 ( .A(n397), .B(n396), .ZN(n700) );
  NAND2_X1 U468 ( .A1(n582), .A2(n596), .ZN(n397) );
  OR2_X1 U469 ( .A1(n659), .A2(n526), .ZN(n399) );
  OR2_X1 U470 ( .A1(n562), .A2(n561), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U472 ( .A(n489), .B(n440), .ZN(n441) );
  XNOR2_X1 U473 ( .A(n478), .B(n402), .ZN(n406) );
  XNOR2_X1 U474 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n551) );
  XNOR2_X1 U475 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U476 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U477 ( .A(n555), .B(KEYINPUT108), .ZN(n737) );
  INV_X1 U478 ( .A(KEYINPUT123), .ZN(n621) );
  XOR2_X1 U479 ( .A(KEYINPUT23), .B(KEYINPUT79), .Z(n404) );
  XNOR2_X1 U480 ( .A(G128), .B(KEYINPUT24), .ZN(n403) );
  XNOR2_X1 U481 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U482 ( .A(n406), .B(n405), .Z(n414) );
  XOR2_X1 U483 ( .A(G125), .B(G140), .Z(n407) );
  XNOR2_X2 U484 ( .A(KEYINPUT10), .B(n407), .ZN(n725) );
  INV_X1 U485 ( .A(KEYINPUT86), .ZN(n408) );
  XNOR2_X1 U486 ( .A(n408), .B(KEYINPUT87), .ZN(n409) );
  NAND2_X1 U487 ( .A1(G234), .A2(n728), .ZN(n410) );
  XOR2_X1 U488 ( .A(KEYINPUT8), .B(n410), .Z(n455) );
  NAND2_X1 U489 ( .A1(G221), .A2(n455), .ZN(n411) );
  INV_X1 U490 ( .A(G902), .ZN(n475) );
  NAND2_X1 U491 ( .A1(n644), .A2(n475), .ZN(n421) );
  XOR2_X1 U492 ( .A(KEYINPUT25), .B(KEYINPUT89), .Z(n417) );
  XNOR2_X1 U493 ( .A(KEYINPUT15), .B(G902), .ZN(n492) );
  NAND2_X1 U494 ( .A1(G234), .A2(n492), .ZN(n415) );
  XNOR2_X1 U495 ( .A(KEYINPUT20), .B(n415), .ZN(n427) );
  NAND2_X1 U496 ( .A1(n427), .A2(G217), .ZN(n416) );
  XNOR2_X1 U497 ( .A(n417), .B(n416), .ZN(n419) );
  INV_X1 U498 ( .A(KEYINPUT88), .ZN(n418) );
  XNOR2_X1 U499 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X2 U500 ( .A(n421), .B(n420), .ZN(n510) );
  NAND2_X1 U501 ( .A1(G237), .A2(G234), .ZN(n422) );
  XNOR2_X1 U502 ( .A(n422), .B(KEYINPUT14), .ZN(n423) );
  NAND2_X1 U503 ( .A1(G952), .A2(n423), .ZN(n697) );
  NOR2_X1 U504 ( .A1(n697), .A2(G953), .ZN(n562) );
  NAND2_X1 U505 ( .A1(G902), .A2(n423), .ZN(n558) );
  NOR2_X1 U506 ( .A1(G900), .A2(n558), .ZN(n424) );
  NAND2_X1 U507 ( .A1(G953), .A2(n424), .ZN(n425) );
  XNOR2_X1 U508 ( .A(KEYINPUT103), .B(n425), .ZN(n426) );
  NOR2_X1 U509 ( .A1(n562), .A2(n426), .ZN(n509) );
  NOR2_X1 U510 ( .A1(n510), .A2(n509), .ZN(n429) );
  AND2_X1 U511 ( .A1(n427), .A2(G221), .ZN(n428) );
  XNOR2_X1 U512 ( .A(n428), .B(KEYINPUT21), .ZN(n683) );
  NAND2_X1 U513 ( .A1(n429), .A2(n683), .ZN(n515) );
  INV_X1 U514 ( .A(n515), .ZN(n445) );
  XNOR2_X2 U515 ( .A(G143), .B(KEYINPUT64), .ZN(n431) );
  XNOR2_X1 U516 ( .A(n433), .B(G131), .ZN(n466) );
  XOR2_X1 U517 ( .A(n466), .B(G137), .Z(n434) );
  XNOR2_X1 U518 ( .A(n435), .B(KEYINPUT3), .ZN(n437) );
  XNOR2_X1 U519 ( .A(G101), .B(KEYINPUT69), .ZN(n436) );
  XNOR2_X1 U520 ( .A(n437), .B(n436), .ZN(n489) );
  XOR2_X1 U521 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n439) );
  NOR2_X1 U522 ( .A1(G953), .A2(G237), .ZN(n460) );
  NAND2_X1 U523 ( .A1(G210), .A2(n460), .ZN(n438) );
  XNOR2_X1 U524 ( .A(n441), .B(G113), .ZN(n442) );
  NAND2_X1 U525 ( .A1(n633), .A2(n475), .ZN(n444) );
  INV_X1 U526 ( .A(G472), .ZN(n443) );
  XNOR2_X2 U527 ( .A(n444), .B(n443), .ZN(n507) );
  XNOR2_X2 U528 ( .A(n507), .B(KEYINPUT6), .ZN(n596) );
  XNOR2_X1 U529 ( .A(n446), .B(KEYINPUT104), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT96), .B(KEYINPUT7), .Z(n448) );
  XNOR2_X1 U531 ( .A(G116), .B(KEYINPUT97), .ZN(n447) );
  XNOR2_X1 U532 ( .A(n448), .B(n447), .ZN(n453) );
  XOR2_X1 U533 ( .A(KEYINPUT98), .B(KEYINPUT95), .Z(n451) );
  XNOR2_X1 U534 ( .A(n449), .B(G107), .ZN(n487) );
  XNOR2_X1 U535 ( .A(n487), .B(KEYINPUT9), .ZN(n450) );
  XNOR2_X1 U536 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U537 ( .A(n453), .B(n452), .Z(n458) );
  NAND2_X1 U538 ( .A1(G217), .A2(n455), .ZN(n456) );
  XNOR2_X1 U539 ( .A(n454), .B(n456), .ZN(n457) );
  XNOR2_X1 U540 ( .A(n458), .B(n457), .ZN(n616) );
  NAND2_X1 U541 ( .A1(n616), .A2(n475), .ZN(n459) );
  XNOR2_X1 U542 ( .A(n459), .B(G478), .ZN(n533) );
  XOR2_X1 U543 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n462) );
  NAND2_X1 U544 ( .A1(n460), .A2(G214), .ZN(n461) );
  XNOR2_X1 U545 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U546 ( .A(n463), .B(n725), .ZN(n468) );
  XNOR2_X2 U547 ( .A(G113), .B(G104), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(n464), .ZN(n465) );
  XNOR2_X1 U549 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U550 ( .A(n468), .B(n467), .ZN(n639) );
  NAND2_X1 U551 ( .A1(n639), .A2(n475), .ZN(n470) );
  XNOR2_X1 U552 ( .A(KEYINPUT13), .B(G475), .ZN(n469) );
  XNOR2_X1 U553 ( .A(n470), .B(n469), .ZN(n521) );
  OR2_X1 U554 ( .A1(n533), .A2(n521), .ZN(n471) );
  XNOR2_X1 U555 ( .A(n471), .B(KEYINPUT99), .ZN(n522) );
  INV_X1 U556 ( .A(n522), .ZN(n663) );
  NAND2_X1 U557 ( .A1(n472), .A2(n522), .ZN(n473) );
  XNOR2_X1 U558 ( .A(n473), .B(KEYINPUT105), .ZN(n476) );
  INV_X1 U559 ( .A(G237), .ZN(n474) );
  NAND2_X1 U560 ( .A1(n475), .A2(n474), .ZN(n493) );
  NAND2_X1 U561 ( .A1(n493), .A2(G214), .ZN(n671) );
  NAND2_X1 U562 ( .A1(n476), .A2(n671), .ZN(n548) );
  XNOR2_X1 U563 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X1 U564 ( .A(n480), .B(n479), .ZN(n485) );
  XOR2_X1 U565 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n483) );
  NAND2_X1 U566 ( .A1(G224), .A2(n728), .ZN(n481) );
  XNOR2_X1 U567 ( .A(n481), .B(G125), .ZN(n482) );
  XNOR2_X1 U568 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U569 ( .A(n485), .B(n484), .ZN(n491) );
  XNOR2_X1 U570 ( .A(n486), .B(KEYINPUT16), .ZN(n488) );
  XNOR2_X1 U571 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U572 ( .A(n490), .B(n489), .ZN(n720) );
  XNOR2_X1 U573 ( .A(n491), .B(n720), .ZN(n627) );
  INV_X1 U574 ( .A(n492), .ZN(n615) );
  AND2_X1 U575 ( .A1(n493), .A2(G210), .ZN(n494) );
  XNOR2_X2 U576 ( .A(n495), .B(n494), .ZN(n527) );
  INV_X1 U577 ( .A(n527), .ZN(n553) );
  XNOR2_X1 U578 ( .A(KEYINPUT36), .B(KEYINPUT84), .ZN(n496) );
  XNOR2_X1 U579 ( .A(n497), .B(n496), .ZN(n504) );
  XNOR2_X1 U580 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U581 ( .A(G140), .B(n500), .Z(n502) );
  NAND2_X1 U582 ( .A1(G227), .A2(n728), .ZN(n501) );
  XNOR2_X1 U583 ( .A(KEYINPUT68), .B(G469), .ZN(n503) );
  INV_X1 U584 ( .A(n681), .ZN(n550) );
  NAND2_X1 U585 ( .A1(n504), .A2(n550), .ZN(n505) );
  INV_X1 U586 ( .A(n521), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n506) );
  XNOR2_X1 U588 ( .A(n506), .B(KEYINPUT102), .ZN(n565) );
  INV_X1 U589 ( .A(n507), .ZN(n514) );
  NAND2_X1 U590 ( .A1(n514), .A2(n671), .ZN(n508) );
  NOR2_X1 U591 ( .A1(n680), .A2(n517), .ZN(n511) );
  XNOR2_X1 U592 ( .A(n511), .B(KEYINPUT90), .ZN(n588) );
  NOR2_X1 U593 ( .A1(n528), .A2(n553), .ZN(n512) );
  XOR2_X1 U594 ( .A(KEYINPUT110), .B(n512), .Z(n513) );
  NOR2_X1 U595 ( .A1(n565), .A2(n513), .ZN(n659) );
  INV_X1 U596 ( .A(n514), .ZN(n587) );
  NOR2_X1 U597 ( .A1(n515), .A2(n587), .ZN(n516) );
  XOR2_X1 U598 ( .A(KEYINPUT28), .B(n516), .Z(n518) );
  NOR2_X1 U599 ( .A1(n518), .A2(n517), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n527), .A2(n671), .ZN(n520) );
  XNOR2_X1 U601 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n519) );
  NAND2_X1 U602 ( .A1(n535), .A2(n358), .ZN(n539) );
  AND2_X1 U603 ( .A1(n533), .A2(n521), .ZN(n655) );
  XNOR2_X1 U604 ( .A(KEYINPUT100), .B(n357), .ZN(n593) );
  XNOR2_X1 U605 ( .A(KEYINPUT72), .B(n593), .ZN(n524) );
  INV_X1 U606 ( .A(KEYINPUT47), .ZN(n523) );
  NAND2_X1 U607 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U608 ( .A1(n539), .A2(n525), .ZN(n526) );
  NOR2_X1 U609 ( .A1(n742), .A2(n399), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n527), .B(KEYINPUT38), .ZN(n531) );
  XNOR2_X1 U611 ( .A(KEYINPUT70), .B(KEYINPUT39), .ZN(n529) );
  XNOR2_X1 U612 ( .A(n530), .B(n529), .ZN(n547) );
  INV_X1 U613 ( .A(n531), .ZN(n672) );
  NAND2_X1 U614 ( .A1(n672), .A2(n671), .ZN(n676) );
  NOR2_X1 U615 ( .A1(n533), .A2(n532), .ZN(n570) );
  INV_X1 U616 ( .A(n570), .ZN(n674) );
  NOR2_X1 U617 ( .A1(n676), .A2(n674), .ZN(n534) );
  XOR2_X1 U618 ( .A(KEYINPUT41), .B(n534), .Z(n698) );
  NAND2_X1 U619 ( .A1(n698), .A2(n535), .ZN(n536) );
  XNOR2_X1 U620 ( .A(n536), .B(KEYINPUT42), .ZN(n744) );
  XOR2_X1 U621 ( .A(KEYINPUT46), .B(KEYINPUT81), .Z(n537) );
  INV_X1 U622 ( .A(n593), .ZN(n675) );
  NAND2_X1 U623 ( .A1(n675), .A2(KEYINPUT47), .ZN(n538) );
  XNOR2_X1 U624 ( .A(n538), .B(KEYINPUT78), .ZN(n542) );
  INV_X1 U625 ( .A(n539), .ZN(n661) );
  NAND2_X1 U626 ( .A1(n661), .A2(KEYINPUT72), .ZN(n540) );
  NAND2_X1 U627 ( .A1(n540), .A2(KEYINPUT47), .ZN(n541) );
  NAND2_X1 U628 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U629 ( .A1(n544), .A2(n543), .ZN(n545) );
  INV_X1 U630 ( .A(n655), .ZN(n666) );
  NOR2_X1 U631 ( .A1(n547), .A2(n666), .ZN(n669) );
  XNOR2_X1 U632 ( .A(KEYINPUT106), .B(n548), .ZN(n549) );
  NOR2_X1 U633 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U634 ( .A1(n554), .A2(n553), .ZN(n555) );
  INV_X1 U635 ( .A(n727), .ZN(n614) );
  INV_X1 U636 ( .A(n558), .ZN(n559) );
  NOR2_X1 U637 ( .A1(G898), .A2(n728), .ZN(n721) );
  NAND2_X1 U638 ( .A1(n559), .A2(n721), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n560), .B(KEYINPUT85), .ZN(n561) );
  NAND2_X1 U640 ( .A1(n358), .A2(n400), .ZN(n563) );
  XNOR2_X1 U641 ( .A(n564), .B(KEYINPUT34), .ZN(n567) );
  INV_X1 U642 ( .A(n565), .ZN(n566) );
  XNOR2_X1 U643 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n568) );
  NAND2_X1 U644 ( .A1(n570), .A2(n683), .ZN(n571) );
  NAND2_X1 U645 ( .A1(n597), .A2(n681), .ZN(n572) );
  XNOR2_X1 U646 ( .A(n572), .B(KEYINPUT101), .ZN(n575) );
  INV_X1 U647 ( .A(n510), .ZN(n573) );
  AND2_X1 U648 ( .A1(n587), .A2(n573), .ZN(n574) );
  INV_X1 U649 ( .A(n597), .ZN(n578) );
  OR2_X1 U650 ( .A1(n681), .A2(n510), .ZN(n576) );
  OR2_X1 U651 ( .A1(n596), .A2(n576), .ZN(n577) );
  NOR2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n579) );
  XNOR2_X1 U654 ( .A(n579), .B(KEYINPUT65), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n581), .B(n580), .ZN(n625) );
  NAND2_X1 U656 ( .A1(n607), .A2(KEYINPUT44), .ZN(n601) );
  NAND2_X1 U657 ( .A1(n582), .A2(n514), .ZN(n688) );
  NOR2_X1 U658 ( .A1(n688), .A2(n589), .ZN(n586) );
  XNOR2_X1 U659 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n584) );
  AND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n591) );
  INV_X1 U661 ( .A(n589), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n652) );
  NAND2_X1 U663 ( .A1(n667), .A2(n652), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT94), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n681), .A2(n510), .ZN(n595) );
  AND2_X1 U667 ( .A1(n359), .A2(n597), .ZN(n648) );
  INV_X1 U668 ( .A(n648), .ZN(n598) );
  AND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U671 ( .A(KEYINPUT82), .ZN(n604) );
  XNOR2_X1 U672 ( .A(n605), .B(n604), .ZN(n612) );
  INV_X1 U673 ( .A(n607), .ZN(n609) );
  INV_X1 U674 ( .A(KEYINPUT44), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U676 ( .A1(n606), .A2(n610), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n364), .A2(G478), .ZN(n618) );
  INV_X1 U679 ( .A(n616), .ZN(n617) );
  XNOR2_X1 U680 ( .A(n618), .B(n617), .ZN(n620) );
  INV_X1 U681 ( .A(G952), .ZN(n619) );
  AND2_X1 U682 ( .A1(n619), .A2(G953), .ZN(n713) );
  NOR2_X2 U683 ( .A1(n620), .A2(n713), .ZN(n622) );
  XNOR2_X1 U684 ( .A(n622), .B(n621), .ZN(G63) );
  XOR2_X1 U685 ( .A(G110), .B(KEYINPUT113), .Z(n624) );
  XOR2_X1 U686 ( .A(n624), .B(n623), .Z(G12) );
  XOR2_X1 U687 ( .A(G119), .B(n625), .Z(G21) );
  NAND2_X1 U688 ( .A1(n707), .A2(G210), .ZN(n629) );
  XOR2_X1 U689 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n626) );
  XNOR2_X1 U690 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U691 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X2 U692 ( .A1(n630), .A2(n713), .ZN(n632) );
  XNOR2_X1 U693 ( .A(KEYINPUT80), .B(KEYINPUT56), .ZN(n631) );
  XNOR2_X1 U694 ( .A(n632), .B(n631), .ZN(G51) );
  NAND2_X1 U695 ( .A1(n707), .A2(G472), .ZN(n635) );
  XOR2_X1 U696 ( .A(KEYINPUT62), .B(n633), .Z(n634) );
  XNOR2_X1 U697 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X2 U698 ( .A1(n636), .A2(n713), .ZN(n638) );
  INV_X1 U699 ( .A(KEYINPUT63), .ZN(n637) );
  XNOR2_X1 U700 ( .A(n638), .B(n637), .ZN(G57) );
  NAND2_X1 U701 ( .A1(n365), .A2(G475), .ZN(n641) );
  XNOR2_X1 U702 ( .A(n639), .B(KEYINPUT59), .ZN(n640) );
  XNOR2_X1 U703 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X2 U704 ( .A1(n642), .A2(n713), .ZN(n643) );
  XNOR2_X1 U705 ( .A(n643), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n364), .A2(G217), .ZN(n646) );
  XOR2_X1 U707 ( .A(KEYINPUT124), .B(n644), .Z(n645) );
  XNOR2_X1 U708 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X1 U709 ( .A1(n647), .A2(n713), .ZN(G66) );
  XOR2_X1 U710 ( .A(G101), .B(n648), .Z(G3) );
  NOR2_X1 U711 ( .A1(n663), .A2(n652), .ZN(n649) );
  XOR2_X1 U712 ( .A(G104), .B(n649), .Z(G6) );
  XOR2_X1 U713 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n651) );
  XNOR2_X1 U714 ( .A(G107), .B(KEYINPUT112), .ZN(n650) );
  XNOR2_X1 U715 ( .A(n651), .B(n650), .ZN(n654) );
  NOR2_X1 U716 ( .A1(n666), .A2(n652), .ZN(n653) );
  XOR2_X1 U717 ( .A(n654), .B(n653), .Z(G9) );
  XOR2_X1 U718 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n657) );
  NAND2_X1 U719 ( .A1(n661), .A2(n655), .ZN(n656) );
  XNOR2_X1 U720 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U721 ( .A(G128), .B(n658), .ZN(G30) );
  XNOR2_X1 U722 ( .A(G143), .B(n659), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n660), .B(KEYINPUT115), .ZN(G45) );
  NAND2_X1 U724 ( .A1(n661), .A2(n522), .ZN(n662) );
  XNOR2_X1 U725 ( .A(n662), .B(G146), .ZN(G48) );
  NOR2_X1 U726 ( .A1(n667), .A2(n663), .ZN(n664) );
  XOR2_X1 U727 ( .A(KEYINPUT116), .B(n664), .Z(n665) );
  XNOR2_X1 U728 ( .A(G113), .B(n665), .ZN(G15) );
  NOR2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U730 ( .A(G116), .B(n668), .Z(G18) );
  XOR2_X1 U731 ( .A(G134), .B(n669), .Z(G36) );
  XOR2_X1 U732 ( .A(KEYINPUT2), .B(n670), .Z(n704) );
  NOR2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n678) );
  NOR2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U737 ( .A1(n679), .A2(n700), .ZN(n694) );
  NAND2_X1 U738 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n682), .B(KEYINPUT50), .ZN(n687) );
  NOR2_X1 U740 ( .A1(n683), .A2(n510), .ZN(n684) );
  XOR2_X1 U741 ( .A(KEYINPUT49), .B(n684), .Z(n685) );
  NOR2_X1 U742 ( .A1(n514), .A2(n685), .ZN(n686) );
  NAND2_X1 U743 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U744 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U745 ( .A(KEYINPUT51), .B(n690), .Z(n691) );
  NAND2_X1 U746 ( .A1(n698), .A2(n691), .ZN(n692) );
  XOR2_X1 U747 ( .A(KEYINPUT120), .B(n692), .Z(n693) );
  NOR2_X1 U748 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n695), .B(KEYINPUT52), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n697), .A2(n696), .ZN(n702) );
  INV_X1 U751 ( .A(n698), .ZN(n699) );
  NOR2_X1 U752 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U753 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U754 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U755 ( .A1(n705), .A2(G953), .ZN(n706) );
  XNOR2_X1 U756 ( .A(n706), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U757 ( .A1(n365), .A2(G469), .ZN(n711) );
  XOR2_X1 U758 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n709) );
  XNOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U761 ( .A1(n713), .A2(n712), .ZN(G54) );
  NAND2_X1 U762 ( .A1(n714), .A2(n728), .ZN(n715) );
  XOR2_X1 U763 ( .A(KEYINPUT125), .B(n715), .Z(n719) );
  NAND2_X1 U764 ( .A1(G953), .A2(G224), .ZN(n716) );
  XNOR2_X1 U765 ( .A(KEYINPUT61), .B(n716), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n717), .A2(G898), .ZN(n718) );
  NAND2_X1 U767 ( .A1(n719), .A2(n718), .ZN(n724) );
  XNOR2_X1 U768 ( .A(n720), .B(G110), .ZN(n722) );
  NOR2_X1 U769 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U770 ( .A(n724), .B(n723), .ZN(G69) );
  XNOR2_X1 U771 ( .A(n726), .B(n725), .ZN(n731) );
  XNOR2_X1 U772 ( .A(n731), .B(n727), .ZN(n729) );
  NAND2_X1 U773 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U774 ( .A(n730), .B(KEYINPUT126), .ZN(n735) );
  XNOR2_X1 U775 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U776 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U777 ( .A1(n733), .A2(G953), .ZN(n734) );
  NAND2_X1 U778 ( .A1(n735), .A2(n734), .ZN(G72) );
  XNOR2_X1 U779 ( .A(G122), .B(KEYINPUT127), .ZN(n736) );
  XNOR2_X1 U780 ( .A(n736), .B(n606), .ZN(G24) );
  XOR2_X1 U781 ( .A(G140), .B(n737), .Z(n738) );
  XNOR2_X1 U782 ( .A(KEYINPUT119), .B(n738), .ZN(G42) );
  XOR2_X1 U783 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n740) );
  XNOR2_X1 U784 ( .A(G125), .B(KEYINPUT118), .ZN(n739) );
  XNOR2_X1 U785 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U786 ( .A(n742), .B(n741), .ZN(G27) );
  XNOR2_X1 U787 ( .A(n743), .B(G131), .ZN(G33) );
  XNOR2_X1 U788 ( .A(G137), .B(n744), .ZN(G39) );
endmodule

