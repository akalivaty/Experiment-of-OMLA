//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n208), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(G58), .A2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  NOR3_X1   g0030(.A1(new_n221), .A2(new_n227), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G226), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  INV_X1    g0038(.A(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  NAND2_X1  g0041(.A1(G68), .A2(G77), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n203), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT66), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G107), .ZN(new_n248));
  INV_X1    g0048(.A(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT7), .B1(new_n254), .B2(new_n225), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(G68), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G159), .ZN(new_n264));
  INV_X1    g0064(.A(G58), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n201), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n266), .B2(new_n222), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n262), .A2(KEYINPUT16), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n226), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT16), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n258), .A2(new_n225), .A3(new_n259), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n201), .B1(new_n274), .B2(new_n260), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n267), .A2(new_n264), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n268), .A2(new_n270), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G87), .ZN(new_n279));
  OAI211_X1 g0079(.A(G226), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n282));
  OAI22_X1  g0082(.A1(new_n252), .A2(new_n253), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n279), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G41), .B2(G45), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n287), .A2(G232), .A3(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n290), .B(G274), .C1(G41), .C2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT8), .B(G58), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n290), .A2(G13), .A3(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n270), .B1(new_n290), .B2(G20), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n298), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT76), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n294), .B1(new_n285), .B2(new_n288), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G190), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n278), .A2(new_n297), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT17), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n289), .B2(new_n295), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n310), .B(new_n294), .C1(new_n285), .C2(new_n288), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT77), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n289), .A2(G179), .A3(new_n295), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT77), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(new_n308), .C2(new_n304), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n312), .A2(new_n315), .B1(new_n303), .B2(new_n278), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT18), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n315), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n278), .A2(new_n303), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT18), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n307), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT78), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n287), .A2(new_n291), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n293), .B1(new_n327), .B2(new_n218), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT67), .Z(new_n329));
  INV_X1    g0129(.A(KEYINPUT69), .ZN(new_n330));
  INV_X1    g0130(.A(G222), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n283), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT3), .B(G33), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT68), .B(G1698), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT69), .A4(G222), .ZN(new_n335));
  INV_X1    g0135(.A(G1698), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n258), .B2(new_n259), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G223), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n333), .A2(new_n202), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n288), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n329), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT72), .B(G200), .Z(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n329), .A2(new_n341), .A3(G190), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n223), .B2(G50), .ZN(new_n348));
  INV_X1    g0148(.A(G150), .ZN(new_n349));
  INV_X1    g0149(.A(new_n263), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n225), .A2(G33), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n348), .B1(new_n349), .B2(new_n350), .C1(new_n351), .C2(new_n298), .ZN(new_n352));
  INV_X1    g0152(.A(new_n299), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n352), .A2(new_n270), .B1(new_n217), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n301), .A2(G50), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT9), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n356), .B(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n326), .B1(new_n347), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n356), .B(KEYINPUT9), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n342), .A2(new_n343), .B1(new_n325), .B2(KEYINPUT10), .ZN(new_n361));
  INV_X1    g0161(.A(new_n326), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(new_n345), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n342), .A2(new_n308), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n356), .C1(G179), .C2(new_n342), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n337), .A2(G238), .ZN(new_n368));
  INV_X1    g0168(.A(G107), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n333), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n333), .A2(new_n334), .A3(G232), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n288), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G244), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n372), .B(new_n293), .C1(new_n373), .C2(new_n327), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(G179), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n308), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n298), .A2(new_n350), .B1(new_n225), .B2(new_n202), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n351), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n270), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n353), .A2(new_n202), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n301), .A2(G77), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n375), .A2(new_n376), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n374), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n382), .A2(KEYINPUT71), .A3(new_n383), .A4(new_n384), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n374), .A2(new_n343), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n388), .A2(new_n390), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n324), .A2(new_n367), .A3(new_n386), .A4(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(G226), .B1(new_n281), .B2(new_n282), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G232), .A2(G1698), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n254), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G97), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n288), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  INV_X1    g0201(.A(new_n327), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G238), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n400), .A2(new_n401), .A3(new_n293), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT74), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT75), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n400), .A2(new_n293), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n406), .A2(new_n407), .A3(G179), .A4(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n400), .A2(new_n403), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n411), .A2(new_n405), .A3(new_n401), .A4(new_n293), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n409), .A3(G179), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n409), .A2(new_n404), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G169), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n419), .A3(G169), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n410), .A2(new_n415), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n350), .A2(new_n217), .B1(new_n351), .B2(new_n202), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n225), .A2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n270), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n301), .A2(G68), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n299), .A2(G68), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT12), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n421), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT78), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n307), .A2(new_n322), .A3(new_n434), .A4(new_n318), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n406), .A2(G190), .A3(new_n409), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n416), .A2(G200), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n431), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT79), .B1(new_n394), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n386), .ZN(new_n441));
  INV_X1    g0241(.A(new_n393), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n441), .B(new_n442), .C1(new_n323), .C2(KEYINPUT78), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .A4(new_n367), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n270), .B1(new_n225), .B2(G116), .ZN(new_n448));
  AOI21_X1  g0248(.A(G20), .B1(new_n257), .B2(G97), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(G33), .B2(G283), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT83), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n449), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(KEYINPUT83), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(G33), .A3(G283), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT87), .A3(new_n449), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n448), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT88), .B1(new_n461), .B2(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(KEYINPUT20), .ZN(new_n463));
  INV_X1    g0263(.A(new_n448), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n459), .A2(KEYINPUT87), .A3(new_n449), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT87), .B1(new_n459), .B2(new_n449), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT88), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n462), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n290), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n299), .A2(new_n472), .A3(new_n226), .A4(new_n269), .ZN(new_n473));
  MUX2_X1   g0273(.A(new_n299), .B(new_n473), .S(G116), .Z(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT5), .B(G41), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(G274), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n226), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n476), .A2(new_n478), .B1(new_n481), .B2(new_n286), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n480), .B1(G270), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n334), .A2(G257), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G264), .A2(G1698), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n333), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G303), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n254), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n288), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n475), .A2(G179), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n490), .A2(new_n389), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(G200), .B2(new_n490), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(new_n471), .A3(new_n474), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n490), .A2(G169), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n475), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g0299(.A(KEYINPUT21), .B(new_n497), .C1(new_n471), .C2(new_n474), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n492), .B(new_n495), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n283), .B2(new_n373), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n337), .A2(G250), .B1(new_n458), .B2(new_n457), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT4), .A4(G244), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n288), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n478), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n287), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n479), .B1(new_n512), .B2(new_n212), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(G190), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT84), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n473), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n473), .A2(new_n517), .ZN(new_n519));
  OAI21_X1  g0319(.A(G97), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n353), .A2(new_n211), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT81), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n255), .B2(new_n261), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT80), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n369), .A2(KEYINPUT6), .A3(G97), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n211), .A2(new_n369), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n526), .B1(new_n529), .B2(KEYINPUT6), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n274), .A2(new_n260), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n525), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n523), .B1(new_n535), .B2(new_n270), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n508), .A2(new_n514), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G200), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n513), .B1(new_n507), .B2(new_n288), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(G190), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n516), .A2(new_n536), .A3(new_n538), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n308), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n539), .A2(new_n310), .ZN(new_n544));
  INV_X1    g0344(.A(new_n270), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n533), .B1(new_n532), .B2(G107), .ZN(new_n546));
  AOI211_X1 g0346(.A(KEYINPUT80), .B(new_n369), .C1(new_n274), .C2(new_n260), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n548), .B2(new_n531), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n543), .B(new_n544), .C1(new_n549), .C2(new_n523), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n542), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n333), .A2(new_n225), .A3(G68), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n528), .A2(new_n209), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n398), .A2(new_n225), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n398), .A2(KEYINPUT19), .A3(G20), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT86), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n553), .B(KEYINPUT86), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n270), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n473), .B(new_n517), .ZN(new_n564));
  INV_X1    g0364(.A(new_n378), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n378), .A2(new_n353), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G244), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  INV_X1    g0370(.A(G238), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n283), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n288), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n478), .A2(G274), .ZN(new_n574));
  INV_X1    g0374(.A(new_n478), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(G250), .A3(new_n287), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n573), .A2(G179), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n576), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n572), .B2(new_n288), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n308), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n568), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n343), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n564), .A2(G87), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(new_n567), .A3(new_n563), .A4(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n580), .A2(G190), .A3(new_n574), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n552), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n551), .B1(new_n542), .B2(new_n550), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n225), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT89), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n333), .A2(KEYINPUT89), .A3(new_n225), .A4(G87), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT22), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n225), .A2(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT23), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT22), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n592), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n225), .A2(G33), .A3(G116), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n596), .A2(new_n598), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT24), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n600), .A2(new_n601), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n598), .A4(new_n596), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n270), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G294), .ZN(new_n609));
  OAI211_X1 g0409(.A(G257), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n609), .B(new_n610), .C1(new_n283), .C2(new_n210), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n288), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n511), .A2(G264), .A3(new_n287), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT91), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT91), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n482), .A2(new_n615), .A3(G264), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n612), .A2(new_n479), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(G200), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n612), .A2(new_n389), .A3(new_n479), .A4(new_n613), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n564), .A2(G107), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n353), .A2(new_n369), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n623), .B(KEYINPUT25), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n608), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT90), .ZN(new_n627));
  AOI221_X4 g0427(.A(new_n480), .B1(new_n482), .B2(G264), .C1(new_n611), .C2(new_n288), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n628), .B2(new_n308), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n616), .A2(new_n614), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(G179), .A3(new_n479), .A4(new_n612), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n612), .A2(new_n479), .A3(new_n613), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(KEYINPUT90), .A3(G169), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n629), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n545), .B1(new_n603), .B2(new_n606), .ZN(new_n635));
  INV_X1    g0435(.A(new_n625), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n626), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n591), .A2(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n447), .A2(new_n502), .A3(new_n590), .A4(new_n639), .ZN(G372));
  INV_X1    g0440(.A(KEYINPUT93), .ZN(new_n641));
  INV_X1    g0441(.A(new_n574), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n642), .B(new_n579), .C1(new_n572), .C2(new_n288), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n577), .B(KEYINPUT92), .C1(new_n643), .C2(new_n308), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n583), .A2(G169), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT92), .B1(new_n646), .B2(new_n577), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n568), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n563), .A2(new_n567), .A3(new_n585), .ZN(new_n649));
  INV_X1    g0449(.A(new_n343), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n580), .B2(new_n574), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n649), .A2(new_n587), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n626), .A2(new_n542), .A3(new_n550), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n641), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n536), .A2(new_n538), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n539), .A2(new_n540), .A3(G190), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n540), .B1(new_n539), .B2(G190), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(G169), .B1(new_n508), .B2(new_n514), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n535), .A2(new_n270), .ZN(new_n662));
  INV_X1    g0462(.A(new_n523), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n657), .A2(new_n660), .B1(new_n664), .B2(new_n544), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT92), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n578), .B2(new_n581), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n644), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n652), .B1(new_n668), .B2(new_n568), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n665), .A2(new_n669), .A3(KEYINPUT93), .A4(new_n626), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n629), .A2(new_n631), .A3(new_n633), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n635), .B2(new_n636), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n672), .B(new_n492), .C1(new_n499), .C2(new_n500), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n656), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n539), .A2(new_n310), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n536), .A2(new_n676), .A3(new_n661), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n648), .A2(new_n675), .A3(new_n677), .A4(new_n653), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT26), .B1(new_n588), .B2(new_n550), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n678), .A2(new_n648), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n447), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT94), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n438), .A2(new_n307), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n433), .B2(new_n386), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n313), .B1(new_n308), .B2(new_n304), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n320), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(new_n317), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n359), .B(new_n363), .C1(new_n685), .C2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(new_n365), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n683), .A2(new_n691), .ZN(G369));
  OR2_X1    g0492(.A1(new_n499), .A2(new_n500), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n492), .ZN(new_n694));
  INV_X1    g0494(.A(G13), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G20), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n290), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n475), .A2(new_n702), .ZN(new_n703));
  MUX2_X1   g0503(.A(new_n694), .B(new_n502), .S(new_n703), .Z(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT95), .Z(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n638), .ZN(new_n707));
  INV_X1    g0507(.A(new_n702), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n637), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n672), .B2(new_n708), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n672), .A2(new_n702), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n702), .B1(new_n693), .B2(new_n492), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(G399));
  NOR2_X1   g0516(.A1(new_n555), .A2(G116), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT96), .Z(new_n718));
  INV_X1    g0518(.A(new_n228), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n718), .A2(new_n290), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n224), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n720), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  NAND4_X1  g0524(.A1(new_n502), .A2(new_n639), .A3(new_n590), .A4(new_n708), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n630), .A2(new_n612), .ZN(new_n726));
  NOR4_X1   g0526(.A1(new_n537), .A2(new_n726), .A3(new_n577), .A4(new_n490), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n491), .A2(new_n643), .A3(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n537), .A3(new_n617), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n702), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  AOI211_X1 g0537(.A(KEYINPUT29), .B(new_n702), .C1(new_n674), .C2(new_n680), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(new_n655), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n673), .A2(new_n669), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n669), .A2(new_n742), .A3(KEYINPUT26), .A4(new_n677), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n648), .A2(KEYINPUT26), .A3(new_n677), .A4(new_n653), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n675), .B1(new_n588), .B2(new_n550), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT97), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n741), .A2(new_n648), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n739), .B1(new_n747), .B2(new_n708), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n738), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n737), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n724), .B1(new_n751), .B2(G1), .ZN(G364));
  AOI21_X1  g0552(.A(new_n290), .B1(new_n696), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n720), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n246), .A2(new_n477), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(KEYINPUT99), .B1(new_n477), .B2(new_n722), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n719), .A2(new_n333), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(KEYINPUT99), .C2(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n719), .A2(new_n254), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT98), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G355), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n760), .B(new_n763), .C1(G116), .C2(new_n228), .ZN(new_n764));
  AND2_X1   g0564(.A1(KEYINPUT100), .A2(G169), .ZN(new_n765));
  NOR2_X1   g0565(.A1(KEYINPUT100), .A2(G169), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n226), .B1(new_n767), .B2(G20), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n756), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT101), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n310), .A2(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n225), .A2(G190), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n254), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n779), .B1(G329), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n225), .A2(new_n389), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n343), .A2(new_n310), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G303), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n225), .B1(new_n780), .B2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n389), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n789), .A2(G294), .B1(G326), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n790), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(G317), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n783), .A2(new_n787), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n343), .A2(new_n310), .A3(new_n776), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT102), .Z(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n784), .A2(new_n775), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n798), .B(new_n802), .C1(G322), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n800), .A2(new_n369), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n254), .B1(new_n804), .B2(G58), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G50), .A2(new_n791), .B1(new_n793), .B2(G68), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(new_n209), .C2(new_n785), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n777), .A2(new_n202), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OR3_X1    g0611(.A1(new_n781), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n789), .A2(G97), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT32), .B1(new_n781), .B2(new_n811), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n806), .A2(new_n809), .A3(new_n810), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n768), .B1(new_n805), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n771), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n774), .B(new_n817), .C1(new_n704), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n705), .A2(G330), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n756), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n705), .A2(G330), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(G396));
  INV_X1    g0623(.A(new_n800), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G87), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n778), .B2(new_n781), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT103), .Z(new_n827));
  INV_X1    g0627(.A(new_n793), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n813), .B1(new_n828), .B2(new_n801), .ZN(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n254), .B1(new_n830), .B2(new_n803), .C1(new_n785), .C2(new_n369), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(G303), .C2(new_n791), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n827), .B(new_n832), .C1(new_n249), .C2(new_n777), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n804), .A2(G143), .ZN(new_n835));
  INV_X1    g0635(.A(new_n777), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G159), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n793), .A2(G150), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n791), .A2(G137), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n835), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n824), .A2(G68), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n333), .B1(new_n265), .B2(new_n788), .C1(new_n785), .C2(new_n217), .ZN(new_n842));
  INV_X1    g0642(.A(new_n840), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(KEYINPUT34), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n841), .B(new_n844), .C1(new_n845), .C2(new_n781), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n833), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n756), .B1(new_n847), .B2(new_n768), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n768), .A2(new_n769), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n202), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n385), .A2(new_n702), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n386), .B1(new_n442), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n441), .A2(new_n708), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n848), .B(new_n850), .C1(new_n770), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n702), .B1(new_n674), .B2(new_n680), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(new_n854), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(new_n737), .Z(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n859), .B2(new_n755), .ZN(G384));
  NAND2_X1  g0660(.A1(new_n432), .A2(new_n702), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n433), .A2(new_n438), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n438), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n432), .B(new_n702), .C1(new_n863), .C2(new_n421), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n734), .A2(new_n735), .A3(new_n855), .A4(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(new_n700), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n320), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(new_n306), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n871), .B2(new_n687), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n321), .A2(new_n868), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n306), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT105), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT105), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT37), .B1(new_n319), .B2(new_n320), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n872), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n870), .B1(new_n688), .B2(new_n307), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n867), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n687), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n874), .B2(new_n882), .ZN(new_n883));
  NOR4_X1   g0683(.A1(new_n874), .A2(new_n316), .A3(KEYINPUT105), .A4(KEYINPUT37), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n876), .B1(new_n871), .B2(new_n877), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n323), .A2(new_n320), .A3(new_n869), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT38), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT40), .B1(new_n866), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI221_X4 g0691(.A(KEYINPUT18), .B1(new_n278), .B2(new_n303), .C1(new_n312), .C2(new_n315), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n870), .B1(new_n894), .B2(new_n307), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n867), .B1(new_n879), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n888), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT106), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n886), .A2(new_n887), .A3(new_n899), .A4(KEYINPUT38), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n866), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n891), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n447), .A2(new_n736), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(G330), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n681), .A2(new_n708), .A3(new_n855), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n853), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT104), .A3(new_n865), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT104), .ZN(new_n911));
  INV_X1    g0711(.A(new_n853), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n857), .B2(new_n855), .ZN(new_n913));
  INV_X1    g0713(.A(new_n865), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n897), .A2(new_n900), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n910), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n433), .A2(new_n702), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT39), .B1(new_n881), .B2(new_n888), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n918), .B(new_n920), .C1(new_n916), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n689), .A2(new_n700), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n434), .B1(new_n894), .B2(new_n307), .ZN(new_n925));
  NOR4_X1   g0725(.A1(new_n925), .A2(new_n366), .A3(new_n441), .A4(new_n442), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n445), .B1(new_n926), .B2(new_n444), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n394), .A2(KEYINPUT79), .A3(new_n439), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n927), .A2(new_n928), .B1(new_n738), .B2(new_n748), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n691), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n924), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n907), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n290), .B2(new_n696), .ZN(new_n933));
  OAI211_X1 g0733(.A(G20), .B(new_n481), .C1(new_n530), .C2(KEYINPUT35), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n249), .B(new_n934), .C1(KEYINPUT35), .C2(new_n530), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT36), .Z(new_n936));
  OAI21_X1  g0736(.A(G77), .B1(new_n265), .B2(new_n201), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n224), .A2(new_n937), .B1(G50), .B2(new_n201), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(G1), .A3(new_n695), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n936), .A3(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n649), .A2(new_n702), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n648), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n669), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n714), .A2(new_n707), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n665), .B1(new_n536), .B2(new_n708), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n550), .B1(new_n947), .B2(new_n672), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT108), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n708), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n947), .B1(new_n550), .B2(new_n708), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n711), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT107), .B(KEYINPUT110), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n962), .B1(new_n961), .B2(new_n963), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n945), .B(new_n957), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n966), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n957), .A2(new_n945), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n964), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n720), .B(KEYINPUT41), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n715), .A2(new_n958), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n715), .A2(new_n958), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n711), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n946), .B1(new_n710), .B2(new_n714), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n820), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n751), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n973), .B1(new_n985), .B2(new_n751), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n754), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT112), .B1(new_n971), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n967), .A2(new_n970), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT112), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(new_n754), .C2(new_n986), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n788), .A2(new_n201), .ZN(new_n993));
  INV_X1    g0793(.A(new_n791), .ZN(new_n994));
  INV_X1    g0794(.A(G143), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n993), .B(new_n996), .C1(G159), .C2(new_n793), .ZN(new_n997));
  INV_X1    g0797(.A(new_n799), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(G77), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n333), .B1(new_n803), .B2(new_n349), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G50), .B2(new_n836), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n786), .A2(G58), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G137), .B2(new_n782), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT113), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n803), .A2(new_n487), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n786), .A2(G116), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT46), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n828), .A2(new_n830), .B1(new_n788), .B2(new_n369), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G311), .B2(new_n791), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n254), .B1(new_n781), .B2(new_n794), .C1(new_n801), .C2(new_n777), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G97), .B2(new_n998), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1005), .B1(new_n1006), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT47), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n756), .B1(new_n1015), .B2(new_n768), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n759), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n772), .B1(new_n228), .B2(new_n378), .C1(new_n240), .C2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(new_n818), .C2(new_n944), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n992), .A2(new_n1019), .ZN(G387));
  NAND2_X1  g0820(.A1(new_n984), .A2(new_n720), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT116), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n751), .B2(new_n983), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n333), .B1(new_n781), .B2(new_n349), .C1(new_n217), .C2(new_n803), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n789), .A2(new_n565), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n994), .B2(new_n811), .C1(new_n298), .C2(new_n828), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(G77), .C2(new_n786), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n201), .B2(new_n777), .C1(new_n211), .C2(new_n800), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n804), .A2(G317), .B1(G322), .B2(new_n791), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n487), .B2(new_n777), .C1(new_n778), .C2(new_n828), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n1032));
  AOI22_X1  g0832(.A1(new_n1031), .A2(new_n1032), .B1(G283), .B2(new_n789), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n830), .B2(new_n785), .C1(new_n1032), .C2(new_n1031), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT49), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n782), .A2(G326), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n254), .C1(new_n799), .C2(new_n249), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT115), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1028), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n756), .B1(new_n1039), .B2(new_n768), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1017), .B1(new_n236), .B2(G45), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n718), .B2(new_n762), .ZN(new_n1042));
  OR3_X1    g0842(.A1(new_n298), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT50), .B1(new_n298), .B2(G50), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1043), .A2(new_n1044), .A3(new_n477), .A4(new_n242), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n718), .A2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1042), .A2(new_n1046), .B1(G107), .B2(new_n228), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n772), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1040), .B(new_n1048), .C1(new_n710), .C2(new_n818), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1023), .B(new_n1049), .C1(new_n753), .C2(new_n982), .ZN(G393));
  OR2_X1    g0850(.A1(new_n980), .A2(KEYINPUT117), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n980), .A2(KEYINPUT117), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n754), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n720), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n980), .B2(new_n984), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n985), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n806), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n782), .A2(G322), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n254), .B1(new_n777), .B2(new_n830), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n828), .A2(new_n487), .B1(new_n788), .B2(new_n249), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G283), .C2(new_n786), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n994), .A2(new_n794), .B1(new_n803), .B2(new_n778), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .A4(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT120), .Z(new_n1066));
  AOI22_X1  g0866(.A1(new_n804), .A2(G159), .B1(G150), .B2(new_n791), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n333), .B1(new_n777), .B2(new_n298), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n828), .A2(new_n217), .B1(new_n788), .B2(new_n202), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n785), .A2(new_n201), .B1(new_n995), .B2(new_n781), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT118), .Z(new_n1074));
  NAND3_X1  g0874(.A1(new_n825), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n756), .B1(new_n1076), .B2(new_n768), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n772), .B1(new_n211), .B2(new_n228), .C1(new_n250), .C2(new_n1017), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n818), .C2(new_n958), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1053), .A2(new_n1056), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(G390));
  AOI21_X1  g0881(.A(new_n921), .B1(new_n897), .B2(new_n900), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n914), .B1(new_n908), .B2(new_n853), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1082), .A2(new_n919), .B1(new_n1083), .B2(new_n918), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n747), .A2(new_n708), .A3(new_n852), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n853), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n865), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n889), .A2(new_n918), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND4_X1   g0889(.A1(new_n734), .A2(new_n735), .A3(new_n855), .A4(new_n865), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(G330), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1084), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n754), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n769), .B1(new_n1082), .B2(new_n919), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n849), .A2(new_n298), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n803), .A2(new_n249), .B1(new_n788), .B2(new_n202), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT122), .Z(new_n1099));
  AOI22_X1  g0899(.A1(G107), .A2(new_n793), .B1(new_n791), .B2(G283), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n254), .C1(new_n211), .C2(new_n777), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G87), .C2(new_n786), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n201), .B2(new_n800), .C1(new_n830), .C2(new_n781), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n777), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n785), .A2(new_n349), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n994), .A2(new_n1109), .B1(new_n788), .B2(new_n811), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G137), .B2(new_n793), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n333), .B1(new_n781), .B2(new_n1112), .C1(new_n845), .C2(new_n803), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G50), .B2(new_n998), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1108), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1103), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n756), .B1(new_n1116), .B2(new_n768), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1097), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1095), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n447), .A2(new_n736), .A3(G330), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1120), .A2(new_n929), .A3(new_n691), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n734), .A2(G330), .A3(new_n735), .A4(new_n855), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1122), .A2(new_n914), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n866), .A2(new_n906), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1086), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n914), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n913), .B1(new_n1091), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1121), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1120), .A2(new_n929), .A3(new_n691), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n909), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1086), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1091), .A2(new_n1132), .A3(new_n1126), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n897), .A2(new_n900), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n919), .B1(new_n1135), .B2(KEYINPUT39), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n918), .B1(new_n909), .B2(new_n865), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1089), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1124), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1084), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1134), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1129), .A2(new_n720), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT121), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1129), .A2(new_n1141), .A3(KEYINPUT121), .A4(new_n720), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1119), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT123), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(G378));
  NAND2_X1  g0948(.A1(new_n1141), .A2(new_n1121), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n916), .A2(new_n898), .A3(new_n1090), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n906), .B1(new_n1150), .B2(new_n890), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n924), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(G330), .B1(new_n891), .B2(new_n902), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1136), .A2(new_n918), .B1(new_n689), .B2(new_n700), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n917), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n356), .A2(new_n869), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n366), .B(new_n1156), .Z(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT55), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT56), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1152), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1149), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1149), .B(KEYINPUT57), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n720), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1159), .A2(new_n769), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n849), .A2(new_n217), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n803), .A2(new_n1109), .B1(new_n788), .B2(new_n349), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n828), .A2(new_n845), .B1(new_n994), .B2(new_n1112), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n786), .C2(new_n1104), .ZN(new_n1171));
  INV_X1    g0971(.A(G137), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n777), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT59), .Z(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n998), .B2(G159), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G33), .B1(new_n782), .B2(G124), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n217), .B1(new_n252), .B2(G41), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G107), .A2(new_n804), .B1(new_n782), .B2(G283), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n378), .B2(new_n777), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n799), .A2(new_n265), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n333), .A2(G41), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n785), .B2(new_n202), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n993), .B1(new_n791), .B2(G116), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n211), .C2(new_n828), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT58), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1177), .A2(new_n1178), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n756), .B1(new_n1188), .B2(new_n768), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1167), .A2(new_n1168), .A3(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT124), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n754), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1166), .A2(new_n1193), .ZN(G375));
  NOR2_X1   g0994(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1130), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n972), .A3(new_n1128), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n254), .B1(new_n781), .B2(new_n487), .C1(new_n801), .C2(new_n803), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1025), .B1(new_n994), .B2(new_n830), .C1(new_n249), .C2(new_n828), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(G97), .C2(new_n786), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n202), .B2(new_n800), .C1(new_n369), .C2(new_n777), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n777), .A2(new_n349), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n333), .B1(new_n803), .B2(new_n1172), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1203), .B(new_n1181), .C1(G128), .C2(new_n782), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1105), .A2(new_n828), .B1(new_n217), .B2(new_n788), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G132), .B2(new_n791), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n811), .C2(new_n785), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1201), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n756), .B1(new_n1208), .B2(new_n768), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n865), .B2(new_n770), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n201), .B2(new_n849), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1195), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n754), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1197), .A2(new_n1213), .ZN(G381));
  INV_X1    g1014(.A(G387), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(G393), .A2(G396), .A3(G390), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1119), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1142), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G375), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(G381), .A2(G384), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1215), .A2(new_n1216), .A3(new_n1219), .A4(new_n1220), .ZN(G407));
  INV_X1    g1021(.A(G213), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1219), .B2(new_n701), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G407), .A2(new_n1223), .ZN(G409));
  NAND2_X1  g1024(.A1(new_n1192), .A2(new_n754), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n1190), .C1(new_n973), .C2(new_n1162), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1218), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1166), .A2(new_n1193), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(G378), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1147), .B1(new_n1232), .B2(new_n1217), .ZN(new_n1233));
  AOI211_X1 g1033(.A(KEYINPUT123), .B(new_n1119), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1235), .A2(G375), .A3(KEYINPUT125), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1228), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1222), .A2(G343), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1054), .B1(new_n1196), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n1128), .C1(new_n1240), .C2(new_n1196), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1213), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(G384), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1237), .A2(new_n1239), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1237), .A2(KEYINPUT126), .A3(new_n1239), .A4(new_n1244), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1238), .A2(G2897), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1244), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1244), .A2(new_n1252), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT127), .B1(new_n1256), .B2(KEYINPUT61), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(G378), .A2(new_n1230), .A3(new_n1229), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT125), .B1(new_n1235), .B2(G375), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1260), .A2(new_n1261), .B1(new_n1227), .B2(new_n1226), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(new_n1238), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1258), .B(new_n1259), .C1(new_n1263), .C2(new_n1255), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1250), .A2(new_n1251), .A3(new_n1257), .A4(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(G393), .B(G396), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n992), .A2(new_n1019), .A3(G390), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G390), .B1(new_n992), .B2(new_n1019), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G387), .A2(new_n1080), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1266), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n992), .A2(new_n1019), .A3(G390), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1265), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT63), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1245), .A2(new_n1277), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1279), .A2(KEYINPUT61), .A3(new_n1256), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1278), .A2(new_n1280), .A3(new_n1273), .A4(new_n1269), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1275), .A2(new_n1281), .ZN(G405));
  OAI22_X1  g1082(.A1(new_n1231), .A2(new_n1236), .B1(new_n1230), .B2(new_n1218), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1244), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1274), .B(new_n1284), .ZN(G402));
endmodule


