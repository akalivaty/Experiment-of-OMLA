//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n474), .A2(G137), .B1(G101), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(new_n465), .B2(new_n475), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(G136), .B2(new_n474), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n463), .B2(new_n464), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n499), .B(new_n502), .C1(new_n464), .C2(new_n463), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT69), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(new_n511), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(new_n516), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT69), .B(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n514), .A2(new_n522), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n513), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n521), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n523), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n525), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT70), .Z(new_n540));
  OAI21_X1  g115(.A(new_n520), .B1(new_n525), .B2(new_n505), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n523), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n542), .A2(new_n543), .B1(new_n512), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n540), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n513), .A2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n521), .A2(G81), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n525), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n512), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n541), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n523), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT71), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n506), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n521), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G299));
  NAND3_X1  g144(.A1(new_n541), .A2(G49), .A3(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n541), .A2(G87), .A3(new_n523), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND3_X1  g148(.A1(new_n541), .A2(G86), .A3(new_n523), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n541), .A2(G48), .A3(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n515), .B2(new_n516), .ZN(new_n577));
  AND2_X1   g152(.A1(G73), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n518), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n525), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT72), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n513), .A2(G47), .B1(new_n521), .B2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(G54), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n512), .A2(new_n587), .B1(new_n588), .B2(new_n506), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT73), .B1(new_n542), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n521), .A2(new_n592), .A3(G92), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n593), .A3(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT74), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n596), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n586), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n586), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  AND2_X1   g183(.A1(new_n599), .A2(new_n601), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G559), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G860), .B2(new_n602), .ZN(G148));
  OAI21_X1  g186(.A(G868), .B1(new_n609), .B2(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n484), .A2(G123), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT75), .Z(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G111), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G2105), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G135), .B2(new_n474), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(G2096), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n481), .A2(new_n476), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2430), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT76), .B(KEYINPUT14), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT77), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(KEYINPUT77), .B1(new_n632), .B2(new_n633), .ZN(new_n637));
  OAI22_X1  g212(.A1(new_n636), .A2(new_n637), .B1(new_n630), .B2(new_n631), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n642), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n661), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n661), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G25), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n474), .A2(G131), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n475), .A2(G107), .ZN(new_n680));
  OAI21_X1  g255(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n681));
  INV_X1    g256(.A(G119), .ZN(new_n682));
  OAI221_X1 g257(.A(new_n679), .B1(new_n680), .B2(new_n681), .C1(new_n483), .C2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT78), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n678), .B1(new_n685), .B2(new_n677), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT35), .B(G1991), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  MUX2_X1   g267(.A(G23), .B(G288), .S(G16), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n696));
  XOR2_X1   g271(.A(KEYINPUT32), .B(G1981), .Z(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NOR3_X1   g273(.A1(new_n692), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n689), .A2(G24), .ZN(new_n701));
  INV_X1    g276(.A(G290), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n689), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT79), .Z(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  OAI221_X1 g282(.A(new_n688), .B1(KEYINPUT34), .B2(new_n700), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(KEYINPUT34), .B2(new_n700), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT80), .B(KEYINPUT36), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G4), .A2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT81), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n609), .B2(new_n689), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1348), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT30), .B(G28), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(new_n677), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G11), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n717), .B(new_n718), .C1(new_n621), .C2(new_n677), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT87), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n677), .A2(G26), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT28), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n484), .A2(G128), .ZN(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n724));
  INV_X1    g299(.A(G116), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G2105), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G140), .B2(new_n474), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n722), .B1(new_n728), .B2(G29), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT82), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2067), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n689), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n689), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1966), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT88), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n689), .A2(G20), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT23), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n606), .B2(new_n689), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1956), .ZN(new_n739));
  NOR4_X1   g314(.A1(new_n720), .A2(new_n731), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n677), .A2(G32), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n476), .A2(G105), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT26), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n742), .B(new_n744), .C1(G141), .C2(new_n474), .ZN(new_n745));
  INV_X1    g320(.A(G129), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n483), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT85), .Z(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G33), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT83), .Z(new_n753));
  NAND3_X1  g328(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n474), .A2(G139), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n481), .A2(G127), .ZN(new_n758));
  NAND2_X1  g333(.A1(G115), .A2(G2104), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n475), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2072), .ZN(new_n763));
  AND2_X1   g338(.A1(KEYINPUT24), .A2(G34), .ZN(new_n764));
  NOR2_X1   g339(.A1(KEYINPUT24), .A2(G34), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n677), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT84), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G160), .B2(G29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(G2084), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n751), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT86), .ZN(new_n771));
  NOR2_X1   g346(.A1(G5), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G171), .B2(G16), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n773), .A2(G1961), .B1(G1966), .B2(new_n733), .ZN(new_n774));
  INV_X1    g349(.A(new_n773), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n553), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G16), .B2(G19), .ZN(new_n778));
  INV_X1    g353(.A(G1341), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n775), .A2(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n677), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n677), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G2078), .Z(new_n783));
  OAI221_X1 g358(.A(new_n783), .B1(G2084), .B2(new_n768), .C1(new_n778), .C2(new_n779), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n677), .A2(G35), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT89), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G162), .B2(new_n677), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT29), .B(G2090), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n748), .B2(new_n749), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n784), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n771), .A2(new_n774), .A3(new_n780), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(KEYINPUT86), .B2(new_n770), .ZN(new_n794));
  AND4_X1   g369(.A1(new_n711), .A2(new_n715), .A3(new_n740), .A4(new_n794), .ZN(G311));
  NAND4_X1  g370(.A1(new_n711), .A2(new_n715), .A3(new_n740), .A4(new_n794), .ZN(G150));
  XNOR2_X1  g371(.A(new_n552), .B(KEYINPUT91), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n521), .A2(G93), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT90), .B(G55), .Z(new_n800));
  OAI221_X1 g375(.A(new_n798), .B1(new_n525), .B2(new_n799), .C1(new_n512), .C2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n797), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n602), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n808));
  AOI21_X1  g383(.A(G860), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n808), .B2(new_n807), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n801), .A2(G860), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(G145));
  XNOR2_X1  g388(.A(new_n747), .B(new_n728), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G164), .ZN(new_n815));
  INV_X1    g390(.A(new_n761), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n474), .A2(G142), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT93), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT92), .ZN(new_n823));
  OR3_X1    g398(.A1(new_n823), .A2(new_n475), .A3(G118), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n821), .A2(KEYINPUT93), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n823), .B1(new_n475), .B2(G118), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G130), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n820), .B(new_n827), .C1(new_n483), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT94), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n625), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(new_n683), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n683), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(KEYINPUT95), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n831), .B(new_n683), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n819), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n490), .B(G160), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n621), .B(new_n841), .Z(new_n842));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n835), .B1(new_n819), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n817), .A2(KEYINPUT97), .A3(new_n818), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n850));
  INV_X1    g425(.A(new_n842), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n837), .A2(new_n834), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(new_n817), .A3(new_n818), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n840), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n840), .A2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n842), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n840), .B2(new_n846), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT40), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n855), .A2(new_n859), .ZN(G395));
  XNOR2_X1  g435(.A(new_n610), .B(new_n804), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n598), .B(G299), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n598), .B(new_n606), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n864), .B(new_n866), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n861), .B(new_n867), .C1(new_n865), .C2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n869), .A3(KEYINPUT100), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT100), .B1(new_n863), .B2(new_n869), .ZN(new_n871));
  XNOR2_X1  g446(.A(G290), .B(G305), .ZN(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G288), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n863), .A2(new_n869), .A3(KEYINPUT100), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  MUX2_X1   g455(.A(new_n801), .B(new_n880), .S(G868), .Z(G295));
  MUX2_X1   g456(.A(new_n801), .B(new_n880), .S(G868), .Z(G331));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n883));
  NAND2_X1  g458(.A1(G171), .A2(G168), .ZN(new_n884));
  NAND2_X1  g459(.A1(G301), .A2(G286), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n804), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n884), .A2(new_n802), .A3(new_n803), .A4(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(new_n867), .C1(new_n868), .C2(new_n865), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n802), .A2(new_n803), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n885), .A4(new_n884), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n862), .B1(new_n886), .B2(new_n804), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n890), .A2(new_n874), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n887), .A3(new_n895), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n898), .A2(new_n868), .B1(new_n888), .B2(new_n894), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n897), .B(new_n848), .C1(new_n899), .C2(new_n874), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n883), .B1(new_n900), .B2(KEYINPUT43), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n890), .A2(new_n896), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n890), .B(new_n896), .C1(KEYINPUT102), .C2(new_n874), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n901), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n902), .B1(new_n901), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n906), .B1(new_n905), .B2(new_n907), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI22_X1  g488(.A1(new_n909), .A2(new_n910), .B1(KEYINPUT44), .B2(new_n913), .ZN(G397));
  XNOR2_X1  g489(.A(new_n728), .B(G2067), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n501), .A2(new_n503), .ZN(new_n916));
  INV_X1    g491(.A(new_n497), .ZN(new_n917));
  AOI21_X1  g492(.A(G1384), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT45), .ZN(new_n919));
  XOR2_X1   g494(.A(KEYINPUT104), .B(G40), .Z(new_n920));
  AND3_X1   g495(.A1(new_n471), .A2(new_n477), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT105), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n915), .A2(KEYINPUT105), .A3(new_n923), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n747), .B(G1996), .ZN(new_n926));
  AOI211_X1 g501(.A(new_n924), .B(new_n925), .C1(new_n923), .C2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n683), .B(new_n687), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n930));
  NAND2_X1  g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n922), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT57), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n563), .A2(new_n568), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n563), .B2(new_n568), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n918), .A2(new_n940), .ZN(new_n941));
  AOI211_X1 g516(.A(KEYINPUT108), .B(G1384), .C1(new_n916), .C2(new_n917), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT50), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n471), .A2(new_n477), .A3(new_n920), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n918), .ZN(new_n946));
  AOI21_X1  g521(.A(G1956), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT106), .B1(new_n918), .B2(KEYINPUT45), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n944), .B1(KEYINPUT45), .B2(new_n918), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n950), .B(new_n951), .C1(G164), .C2(G1384), .ZN(new_n952));
  XNOR2_X1  g527(.A(KEYINPUT56), .B(G2072), .ZN(new_n953));
  AND4_X1   g528(.A1(new_n948), .A2(new_n949), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n939), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT108), .B1(G164), .B2(G1384), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  INV_X1    g532(.A(new_n503), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n502), .B1(new_n481), .B2(new_n499), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n940), .B(new_n957), .C1(new_n960), .C2(new_n497), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n921), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n956), .A2(new_n961), .A3(new_n921), .A4(KEYINPUT117), .ZN(new_n965));
  AOI21_X1  g540(.A(G2067), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n956), .A2(new_n945), .A3(new_n961), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n957), .B1(new_n960), .B2(new_n497), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n944), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(G1348), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n602), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1956), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n945), .B1(new_n956), .B2(new_n961), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n921), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n949), .A2(new_n948), .A3(new_n952), .A4(new_n953), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n975), .A2(new_n938), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n955), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT118), .Z(new_n979));
  OAI21_X1  g554(.A(KEYINPUT60), .B1(new_n966), .B2(new_n970), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n609), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n982));
  AND3_X1   g557(.A1(new_n981), .A2(new_n971), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n981), .B2(new_n971), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n986));
  AOI21_X1  g561(.A(new_n938), .B1(new_n975), .B2(new_n976), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n977), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT121), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n975), .A2(new_n938), .A3(new_n989), .A4(new_n976), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n955), .A2(KEYINPUT61), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n975), .A2(new_n938), .A3(new_n976), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(KEYINPUT121), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT58), .B(G1341), .Z(new_n995));
  NAND3_X1  g570(.A1(new_n964), .A2(new_n965), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT119), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n964), .A2(new_n999), .A3(new_n965), .A4(new_n995), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n949), .A2(new_n948), .A3(new_n952), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(G1996), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n553), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT59), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n997), .B(new_n1000), .C1(G1996), .C2(new_n1001), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT59), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n553), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n994), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n985), .B1(new_n1008), .B2(KEYINPUT122), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT122), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n1010), .B(new_n994), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n979), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1971), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1001), .A2(KEYINPUT107), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G2090), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n967), .A2(new_n969), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT107), .B1(new_n1001), .B2(new_n1013), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT109), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1001), .A2(new_n1013), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1019), .A2(new_n1024), .A3(G8), .A4(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n962), .A2(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n575), .A2(new_n574), .A3(new_n1034), .A4(new_n579), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT49), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1032), .A2(new_n1037), .A3(KEYINPUT112), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n962), .A3(G8), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n570), .A2(new_n571), .A3(G1976), .A4(new_n572), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(G8), .A3(new_n962), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(G288), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1032), .A2(new_n1045), .A3(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1043), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1031), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n943), .A2(KEYINPUT114), .A3(new_n946), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n973), .B2(new_n974), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1056), .A3(new_n1015), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1053), .B1(new_n1057), .B2(new_n1020), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT115), .B1(new_n1058), .B2(new_n1030), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1020), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n943), .A2(new_n946), .ZN(new_n1062));
  AOI21_X1  g637(.A(G2090), .B1(new_n1062), .B2(new_n1055), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n1063), .B2(new_n1054), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1060), .B(new_n1029), .C1(new_n1064), .C2(new_n1053), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1052), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1961), .B1(new_n967), .B2(new_n969), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1001), .A2(G2078), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n918), .A2(KEYINPUT45), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(G2078), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(G40), .A3(G160), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1070), .B1(new_n919), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n956), .B2(new_n961), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n921), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1072), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1070), .A2(G301), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT126), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT54), .B(new_n1075), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1966), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT116), .B(G2084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n967), .A2(new_n969), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G286), .A2(G8), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1053), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G286), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(KEYINPUT51), .ZN(new_n1097));
  OAI211_X1 g672(.A(G8), .B(new_n1097), .C1(new_n1089), .C2(G286), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT125), .B(KEYINPUT54), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1074), .A2(G171), .ZN(new_n1101));
  AOI21_X1  g676(.A(G301), .B1(new_n1070), .B2(new_n1079), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1066), .A2(new_n1084), .A3(new_n1099), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1012), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1024), .A2(G8), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1106), .A2(new_n1051), .A3(new_n1030), .A4(new_n1019), .ZN(new_n1107));
  OR2_X1    g682(.A1(G288), .A2(G1976), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1035), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1032), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT113), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1043), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT113), .B(new_n1111), .C1(new_n1031), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1031), .A2(new_n1051), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1065), .A2(new_n1059), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1099), .A2(KEYINPUT62), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1093), .A2(new_n1120), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1102), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1112), .A2(new_n1115), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1090), .A2(G286), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1117), .A2(new_n1031), .A3(new_n1051), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(KEYINPUT63), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1019), .A2(G8), .A3(new_n1024), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1029), .B2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1125), .A2(new_n1126), .B1(new_n1116), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1123), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n934), .B1(new_n1105), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n922), .A2(G1996), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT46), .Z(new_n1134));
  OAI21_X1  g709(.A(new_n923), .B1(new_n915), .B2(new_n747), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT47), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n930), .A2(new_n922), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT48), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n929), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n927), .A2(new_n685), .A3(new_n687), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n728), .A2(G2067), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n922), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT127), .B1(new_n1132), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1066), .A2(new_n1084), .A3(new_n1099), .A4(new_n1103), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1005), .A2(new_n1006), .A3(new_n553), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1006), .B1(new_n1005), .B2(new_n553), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1010), .B1(new_n1150), .B2(new_n994), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1008), .A2(KEYINPUT122), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n985), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1147), .B1(new_n1153), .B2(new_n979), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1119), .A2(new_n1102), .A3(new_n1121), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1111), .B1(new_n1031), .B2(new_n1113), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT113), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1158), .A2(new_n1066), .B1(new_n1161), .B2(new_n1114), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n933), .B1(new_n1154), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(new_n1144), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1146), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g742(.A1(G401), .A2(new_n461), .A3(G227), .A4(G229), .ZN(new_n1169));
  OAI21_X1  g743(.A(new_n1169), .B1(new_n849), .B2(new_n854), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1170), .A2(new_n913), .ZN(G308));
  OAI221_X1 g745(.A(new_n1169), .B1(new_n911), .B2(new_n912), .C1(new_n849), .C2(new_n854), .ZN(G225));
endmodule


