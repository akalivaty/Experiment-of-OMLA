//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n208), .B(new_n210), .C1(G113gat), .C2(new_n209), .ZN(new_n211));
  XNOR2_X1  g010(.A(G127gat), .B(G134gat), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n207), .A2(G120gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n209), .A2(G113gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n212), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(G155gat), .B2(G162gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G148gat), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G141gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G155gat), .B(G162gat), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT2), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n229), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n229), .A2(new_n239), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n239), .A3(KEYINPUT81), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(KEYINPUT3), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n252), .A2(new_n211), .B1(new_n219), .B2(new_n220), .ZN(new_n253));
  INV_X1    g052(.A(new_n243), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n251), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n253), .A2(new_n254), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(KEYINPUT83), .A3(new_n256), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n222), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n260), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n268), .B2(new_n251), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n255), .B1(new_n222), .B2(new_n243), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n254), .A3(new_n262), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n272), .A2(KEYINPUT84), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT84), .B1(new_n272), .B2(new_n273), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n249), .B(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n205), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT6), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n270), .A2(new_n205), .A3(new_n276), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n281), .B2(new_n277), .ZN(new_n282));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286));
  INV_X1    g085(.A(G169gat), .ZN(new_n287));
  INV_X1    g086(.A(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n290));
  NOR2_X1   g089(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(KEYINPUT66), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT66), .B1(new_n294), .B2(new_n289), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g095(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n297), .A2(KEYINPUT23), .A3(new_n287), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT24), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n299), .B(new_n304), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n286), .B1(new_n296), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n292), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT70), .B(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n306), .A2(new_n308), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n286), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT68), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n287), .A3(new_n288), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT68), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(KEYINPUT23), .A3(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n325), .A2(KEYINPUT69), .A3(new_n304), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT69), .B1(new_n325), .B2(new_n304), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n316), .B(new_n321), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n302), .A2(new_n303), .B1(new_n289), .B2(KEYINPUT26), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT26), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n323), .A2(new_n332), .A3(new_n324), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n331), .A2(new_n333), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  INV_X1    g133(.A(G183gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n318), .B1(new_n335), .B2(KEYINPUT27), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT28), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(KEYINPUT70), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT27), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n343), .B2(new_n337), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT71), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n336), .B1(new_n317), .B2(KEYINPUT27), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n347), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n334), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n329), .A2(new_n330), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n334), .B(new_n351), .C1(new_n346), .C2(new_n348), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT71), .B1(new_n347), .B2(KEYINPUT28), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n343), .A2(new_n337), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n345), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n357), .A3(new_n339), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n351), .B1(new_n358), .B2(new_n334), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n329), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n330), .A2(KEYINPUT29), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n350), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G218gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G211gat), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G218gat), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT78), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G211gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT22), .B1(new_n371), .B2(G218gat), .ZN(new_n372));
  XOR2_X1   g171(.A(G197gat), .B(G204gat), .Z(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT22), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT77), .B(G211gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n363), .ZN(new_n377));
  INV_X1    g176(.A(new_n373), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n364), .A2(new_n366), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n374), .A2(KEYINPUT79), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT79), .B1(new_n374), .B2(new_n382), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n330), .B(new_n329), .C1(new_n353), .C2(new_n359), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n329), .A2(new_n349), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n361), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT80), .B1(new_n391), .B2(new_n385), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n393), .B(new_n386), .C1(new_n388), .C2(new_n390), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n285), .B(new_n387), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n361), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n329), .B2(new_n349), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n349), .A2(KEYINPUT72), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n400), .A2(new_n352), .B1(new_n312), .B2(new_n328), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n401), .B2(new_n330), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n393), .B1(new_n402), .B2(new_n386), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n391), .A2(KEYINPUT80), .A3(new_n385), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n285), .A4(new_n387), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n387), .B1(new_n392), .B2(new_n394), .ZN(new_n407));
  INV_X1    g206(.A(new_n285), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n282), .A2(new_n397), .A3(new_n406), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(G22gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT31), .B(G50gat), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT29), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n241), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n372), .A2(new_n373), .A3(new_n367), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n381), .B1(new_n377), .B2(new_n378), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n374), .A2(KEYINPUT79), .A3(new_n382), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n418), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n379), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n372), .B2(new_n373), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n254), .B1(new_n428), .B2(new_n240), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n416), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(KEYINPUT85), .B(new_n416), .C1(new_n424), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n241), .A2(new_n417), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n383), .B2(new_n384), .ZN(new_n436));
  INV_X1    g235(.A(new_n416), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT29), .B1(new_n374), .B2(new_n382), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n247), .B1(new_n438), .B2(KEYINPUT3), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n415), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n414), .B(new_n440), .C1(new_n432), .C2(new_n433), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n413), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n240), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n243), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n436), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT85), .B1(new_n447), .B2(new_n416), .ZN(new_n448));
  INV_X1    g247(.A(new_n433), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n441), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n414), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n415), .A3(new_n441), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n412), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n444), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n410), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT36), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT76), .B(KEYINPUT34), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n360), .A2(new_n253), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n222), .B(new_n329), .C1(new_n353), .C2(new_n359), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G227gat), .ZN(new_n462));
  INV_X1    g261(.A(G233gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n464), .B(new_n457), .C1(new_n459), .C2(new_n460), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G43gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n459), .A2(new_n464), .A3(new_n460), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT33), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n471), .A2(KEYINPUT75), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(KEYINPUT75), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(KEYINPUT33), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(KEYINPUT32), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n468), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n466), .ZN(new_n482));
  INV_X1    g281(.A(new_n467), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n476), .A2(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n456), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n480), .ZN(new_n486));
  INV_X1    g285(.A(new_n468), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n476), .A3(new_n480), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT36), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n455), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n455), .A2(new_n485), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n405), .B2(new_n387), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT37), .B1(new_n362), .B2(new_n386), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n392), .B2(new_n394), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n408), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT38), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n272), .A2(new_n273), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n272), .A2(KEYINPUT84), .A3(new_n273), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n248), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n506), .A2(new_n271), .B1(new_n265), .B2(new_n269), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n205), .B(KEYINPUT87), .Z(new_n508));
  OAI211_X1 g307(.A(new_n279), .B(new_n280), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n509), .A2(new_n395), .A3(new_n278), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n496), .B1(new_n362), .B2(new_n385), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n391), .A2(new_n386), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT38), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n499), .A3(new_n408), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT89), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(new_n499), .A3(new_n516), .A4(new_n408), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n501), .A2(new_n510), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n397), .A2(new_n406), .A3(new_n409), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n249), .B1(new_n274), .B2(new_n275), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT39), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n251), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n505), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n250), .B1(new_n523), .B2(new_n249), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT88), .B1(new_n268), .B2(new_n251), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n267), .A2(new_n260), .A3(new_n526), .A4(new_n250), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(KEYINPUT39), .A3(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n522), .B(new_n508), .C1(new_n524), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n507), .A2(new_n508), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n527), .A2(KEYINPUT39), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n525), .B(new_n533), .C1(new_n506), .C2(new_n250), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(KEYINPUT40), .A3(new_n508), .A4(new_n522), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n454), .B1(new_n519), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT90), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n442), .A2(new_n443), .A3(new_n413), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n412), .B1(new_n451), .B2(new_n452), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n481), .B2(new_n484), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT35), .B1(new_n546), .B2(new_n410), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n454), .B1(new_n488), .B2(new_n489), .ZN(new_n550));
  INV_X1    g349(.A(new_n410), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(KEYINPUT92), .A3(KEYINPUT35), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n519), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n509), .B2(new_n278), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n550), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n495), .A2(new_n542), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT16), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(G1gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n562), .B(KEYINPUT95), .ZN(new_n567));
  INV_X1    g366(.A(G1gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G8gat), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n572), .A3(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT96), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n576), .A3(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n580));
  AOI21_X1  g379(.A(G36gat), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G29gat), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n582), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n583));
  OR3_X1    g382(.A1(new_n581), .A2(KEYINPUT15), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT15), .B1(new_n581), .B2(new_n583), .ZN(new_n585));
  XNOR2_X1  g384(.A(G43gat), .B(G50gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n585), .B2(new_n586), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT17), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT97), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n588), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT98), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n588), .A2(KEYINPUT17), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n588), .A2(KEYINPUT17), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n575), .A2(new_n577), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n591), .A2(new_n592), .A3(new_n594), .A4(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT18), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(KEYINPUT98), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n593), .A2(KEYINPUT98), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n603), .A2(new_n604), .B1(new_n597), .B2(new_n598), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(KEYINPUT18), .A3(new_n592), .A4(new_n591), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n594), .B1(new_n588), .B2(new_n574), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n592), .B(KEYINPUT13), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n602), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n611));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G197gat), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT11), .B(G169gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  AND3_X1   g416(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n610), .B2(new_n611), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT105), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G71gat), .B(G78gat), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G57gat), .B(G64gat), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n625), .B1(new_n628), .B2(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G85gat), .A2(G92gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  NAND2_X1  g434(.A1(G99gat), .A2(G106gat), .ZN(new_n636));
  INV_X1    g435(.A(G85gat), .ZN(new_n637));
  INV_X1    g436(.A(G92gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(KEYINPUT8), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT101), .ZN(new_n641));
  XOR2_X1   g440(.A(G99gat), .B(G106gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n640), .B(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n642), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n632), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n642), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n641), .A2(new_n643), .ZN(new_n650));
  INV_X1    g449(.A(new_n632), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n624), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(KEYINPUT10), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n644), .B2(new_n647), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT102), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n622), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n622), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n648), .A2(new_n660), .A3(new_n652), .ZN(new_n661));
  XOR2_X1   g460(.A(G120gat), .B(G148gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT104), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  NAND3_X1  g464(.A1(new_n659), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(new_n659), .B2(new_n661), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n621), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(KEYINPUT105), .A3(new_n666), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT21), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n632), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(G231gat), .A2(G233gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(G127gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n574), .B1(KEYINPUT21), .B2(new_n651), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n236), .ZN(new_n683));
  XOR2_X1   g482(.A(G183gat), .B(G211gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n681), .B(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT102), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT102), .B1(new_n649), .B2(new_n650), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n588), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n656), .A2(new_n589), .A3(new_n657), .ZN(new_n692));
  NAND3_X1  g491(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(G190gat), .B(G218gat), .Z(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT99), .ZN(new_n698));
  XNOR2_X1  g497(.A(G134gat), .B(G162gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n695), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n691), .A2(new_n692), .A3(new_n701), .A4(new_n693), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n696), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n700), .B1(new_n696), .B2(new_n702), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n620), .A2(new_n673), .A3(new_n688), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n561), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n282), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n568), .ZN(G1324gat));
  INV_X1    g512(.A(new_n707), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n572), .B1(new_n714), .B2(new_n519), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT16), .B(G8gat), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n707), .A2(new_n555), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT42), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(KEYINPUT42), .B2(new_n717), .ZN(G1325gat));
  NOR2_X1   g518(.A1(new_n481), .A2(new_n484), .ZN(new_n720));
  OR3_X1    g519(.A1(new_n707), .A2(G15gat), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n485), .A2(new_n490), .ZN(new_n722));
  OAI21_X1  g521(.A(G15gat), .B1(new_n707), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n714), .A2(new_n454), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT107), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  INV_X1    g527(.A(new_n705), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT92), .B1(new_n552), .B2(KEYINPUT35), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT35), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n548), .B(new_n731), .C1(new_n550), .C2(new_n551), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n559), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n518), .A2(new_n537), .A3(new_n540), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n540), .B1(new_n518), .B2(new_n537), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n492), .B(new_n494), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n729), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n620), .A2(new_n673), .A3(new_n687), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n711), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n582), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT45), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n558), .B1(new_n549), .B2(new_n553), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n491), .B1(new_n539), .B2(new_n541), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n743), .B(new_n705), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n746), .B(KEYINPUT108), .C1(new_n737), .C2(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n748), .B(KEYINPUT44), .C1(new_n560), .C2(new_n729), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n747), .A2(new_n749), .A3(new_n740), .A4(new_n738), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G29gat), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n750), .A2(new_n751), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n742), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n742), .B(KEYINPUT110), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1328gat));
  INV_X1    g558(.A(G36gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n739), .A2(new_n760), .A3(new_n519), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n747), .A2(new_n749), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n765), .A2(new_n519), .A3(new_n738), .ZN(new_n766));
  OAI221_X1 g565(.A(new_n764), .B1(new_n762), .B2(new_n761), .C1(new_n766), .C2(new_n760), .ZN(G1329gat));
  INV_X1    g566(.A(new_n722), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n747), .A2(new_n749), .A3(new_n768), .A4(new_n738), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G43gat), .ZN(new_n770));
  INV_X1    g569(.A(G43gat), .ZN(new_n771));
  INV_X1    g570(.A(new_n720), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n739), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT47), .Z(G1330gat));
  NAND4_X1  g574(.A1(new_n747), .A2(new_n749), .A3(new_n454), .A4(new_n738), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G50gat), .ZN(new_n777));
  INV_X1    g576(.A(G50gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n739), .A2(new_n778), .A3(new_n454), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT48), .Z(G1331gat));
  NOR2_X1   g580(.A1(new_n744), .A2(new_n745), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n620), .A2(new_n687), .A3(new_n729), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n782), .A2(new_n672), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n740), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n519), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT49), .B(G64gat), .Z(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(G1333gat));
  NAND2_X1  g589(.A1(new_n784), .A2(new_n768), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n720), .A2(G71gat), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n791), .A2(G71gat), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n784), .A2(new_n454), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT112), .B(G78gat), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n795), .B(new_n796), .ZN(G1335gat));
  INV_X1    g596(.A(new_n620), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n798), .A2(new_n672), .A3(new_n687), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n765), .A2(new_n740), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G85gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n687), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n705), .B(new_n802), .C1(new_n744), .C2(new_n745), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n805), .A2(new_n637), .A3(new_n740), .A4(new_n673), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(G1336gat));
  NAND3_X1  g606(.A1(new_n765), .A2(new_n519), .A3(new_n799), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n672), .A2(G92gat), .A3(new_n555), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n803), .A2(new_n804), .ZN(new_n813));
  MUX2_X1   g612(.A(new_n805), .B(new_n813), .S(KEYINPUT113), .Z(new_n814));
  AOI22_X1  g613(.A1(new_n814), .A2(new_n810), .B1(new_n808), .B2(G92gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(G1337gat));
  NOR2_X1   g616(.A1(new_n720), .A2(G99gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n805), .A2(new_n673), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n765), .A2(new_n768), .A3(new_n799), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G99gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n820), .A2(new_n821), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(G1338gat));
  NAND3_X1  g624(.A1(new_n765), .A2(new_n454), .A3(new_n799), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G106gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n672), .A2(G106gat), .A3(new_n545), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT53), .B1(new_n805), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n814), .A2(new_n828), .B1(new_n826), .B2(G106gat), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(G1339gat));
  INV_X1    g632(.A(new_n653), .ZN(new_n834));
  OAI211_X1 g633(.A(KEYINPUT10), .B(new_n651), .C1(new_n689), .C2(new_n690), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n660), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n659), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n622), .C1(new_n653), .C2(new_n658), .ZN(new_n839));
  INV_X1    g638(.A(new_n665), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n839), .A2(KEYINPUT115), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT115), .B1(new_n839), .B2(new_n840), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT55), .B(new_n837), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n666), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n844), .B(new_n847), .C1(new_n618), .C2(new_n619), .ZN(new_n848));
  INV_X1    g647(.A(new_n617), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n602), .A2(new_n606), .A3(new_n609), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n592), .B1(new_n605), .B2(new_n591), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n607), .A2(new_n608), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n615), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n671), .A2(new_n669), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n705), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n847), .A2(new_n666), .A3(new_n843), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n705), .A2(new_n850), .A3(new_n853), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n858), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n860), .A2(new_n844), .A3(KEYINPUT116), .A4(new_n847), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n688), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n783), .A2(new_n673), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n711), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n546), .A2(new_n519), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n798), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n454), .B1(new_n863), .B2(new_n864), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n711), .A2(new_n519), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n869), .A2(new_n772), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n620), .A2(new_n207), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n867), .B2(new_n673), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n672), .A2(new_n209), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n871), .B2(new_n875), .ZN(G1341gat));
  NAND3_X1  g675(.A1(new_n865), .A2(new_n866), .A3(new_n687), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n678), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n688), .A2(new_n678), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n871), .B2(new_n881), .ZN(G1342gat));
  INV_X1    g681(.A(G134gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n883), .A3(new_n705), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(KEYINPUT56), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n705), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(G134gat), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT118), .B(new_n883), .C1(new_n871), .C2(new_n705), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n885), .B(new_n886), .C1(new_n889), .C2(new_n890), .ZN(G1343gat));
  NAND2_X1  g690(.A1(new_n722), .A2(new_n454), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n555), .B1(new_n892), .B2(KEYINPUT119), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(KEYINPUT119), .B2(new_n892), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n865), .A2(new_n230), .A3(new_n798), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n870), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n768), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n863), .A2(new_n864), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n454), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n902), .B(new_n545), .C1(new_n863), .C2(new_n864), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n798), .B(new_n899), .C1(new_n901), .C2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n897), .B1(new_n904), .B2(G141gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n905), .B(new_n906), .ZN(G1344gat));
  AND2_X1   g706(.A1(new_n865), .A2(new_n894), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n232), .A3(new_n673), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G148gat), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n901), .A2(new_n903), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n768), .A3(new_n898), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n913), .B2(new_n673), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n857), .A2(new_n858), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n854), .B1(new_n620), .B2(new_n857), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n729), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n864), .B1(new_n917), .B2(new_n687), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n454), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n902), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n900), .A2(KEYINPUT57), .A3(new_n454), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n922), .A2(new_n722), .A3(new_n673), .A4(new_n870), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n910), .B1(new_n923), .B2(G148gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n909), .B1(new_n914), .B2(new_n924), .ZN(G1345gat));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n236), .A3(new_n687), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n913), .A2(new_n687), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n236), .ZN(G1346gat));
  OAI211_X1 g727(.A(new_n705), .B(new_n899), .C1(new_n901), .C2(new_n903), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n237), .B1(new_n929), .B2(KEYINPUT121), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(KEYINPUT121), .B2(new_n929), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n908), .A2(new_n237), .A3(new_n705), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1347gat));
  NAND2_X1  g732(.A1(new_n550), .A2(new_n519), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n740), .B(new_n934), .C1(new_n863), .C2(new_n864), .ZN(new_n935));
  AOI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n798), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n740), .A2(new_n555), .A3(new_n720), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n869), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n620), .A2(new_n287), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  AOI21_X1  g739(.A(G176gat), .B1(new_n935), .B2(new_n673), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n672), .B1(new_n297), .B2(new_n298), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n938), .B2(new_n942), .ZN(G1349gat));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT60), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT27), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G183gat), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n935), .A2(new_n947), .A3(new_n338), .A4(new_n687), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n869), .A2(new_n687), .A3(new_n937), .ZN(new_n949));
  INV_X1    g748(.A(new_n317), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n945), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n944), .A2(KEYINPUT60), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n952), .B(new_n953), .Z(G1350gat));
  NAND3_X1  g753(.A1(new_n935), .A2(new_n318), .A3(new_n705), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n869), .A2(new_n705), .A3(new_n937), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT123), .ZN(G1351gat));
  NOR2_X1   g760(.A1(new_n892), .A2(new_n555), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n900), .A2(new_n711), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n798), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n740), .A2(new_n555), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT57), .B1(new_n918), .B2(new_n454), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n722), .B(new_n965), .C1(new_n903), .C2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n798), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n672), .A2(G204gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n963), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT125), .Z(new_n974));
  OAI21_X1  g773(.A(G204gat), .B1(new_n967), .B2(new_n672), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n971), .B1(new_n963), .B2(new_n972), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT124), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n376), .A3(new_n687), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n922), .A2(new_n722), .A3(new_n687), .A4(new_n965), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT63), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n365), .B1(KEYINPUT126), .B2(new_n981), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  OAI21_X1  g785(.A(G218gat), .B1(new_n967), .B2(new_n729), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n963), .A2(new_n363), .A3(new_n705), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n987), .A2(KEYINPUT127), .A3(new_n988), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1355gat));
endmodule


