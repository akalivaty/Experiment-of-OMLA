//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  INV_X1    g000(.A(G57gat), .ZN(new_n202));
  INV_X1    g001(.A(G64gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205));
  AND2_X1   g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(KEYINPUT9), .ZN(new_n207));
  NOR2_X1   g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT95), .ZN(new_n209));
  NAND2_X1  g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(new_n211), .C1(new_n209), .C2(new_n210), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT96), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n203), .B1(new_n213), .B2(new_n202), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n215), .A2(G71gat), .A3(G78gat), .ZN(new_n216));
  OAI221_X1 g015(.A(new_n214), .B1(new_n213), .B2(new_n205), .C1(new_n216), .C2(new_n206), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT21), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(new_n217), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT98), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT98), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n227), .A3(new_n217), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n229), .A2(KEYINPUT21), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT16), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n231), .A2(G1gat), .ZN(new_n236));
  OAI21_X1  g035(.A(G8gat), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G8gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n234), .B(new_n238), .C1(G1gat), .C2(new_n231), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT92), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT92), .B1(new_n237), .B2(new_n239), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(G183gat), .B1(new_n230), .B2(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n240), .A2(new_n241), .ZN(new_n244));
  INV_X1    g043(.A(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n229), .A2(KEYINPUT21), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT97), .ZN(new_n249));
  INV_X1    g048(.A(G231gat), .ZN(new_n250));
  INV_X1    g049(.A(G233gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT97), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n243), .A2(new_n253), .A3(new_n247), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n249), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n224), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n256), .A2(new_n257), .A3(new_n224), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n221), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n220), .A3(new_n258), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT100), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT103), .ZN(new_n266));
  INV_X1    g065(.A(G50gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G43gat), .ZN(new_n268));
  INV_X1    g067(.A(G43gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G50gat), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT15), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT91), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .A4(KEYINPUT15), .ZN(new_n274));
  OR2_X1    g073(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(G29gat), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT14), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(G29gat), .B2(G36gat), .ZN(new_n279));
  INV_X1    g078(.A(G29gat), .ZN(new_n280));
  INV_X1    g079(.A(G36gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT14), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n274), .A2(new_n277), .A3(new_n279), .A4(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n268), .A2(new_n270), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT15), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n273), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT88), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n282), .A2(new_n279), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n277), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n282), .B2(new_n279), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n271), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT90), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT90), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n293), .B(new_n271), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G85gat), .A2(G92gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT7), .ZN(new_n297));
  NAND2_X1  g096(.A1(G99gat), .A2(G106gat), .ZN(new_n298));
  INV_X1    g097(.A(G85gat), .ZN(new_n299));
  INV_X1    g098(.A(G92gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(KEYINPUT8), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n301), .A2(KEYINPUT101), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(KEYINPUT101), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G99gat), .B(G106gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n301), .B(KEYINPUT101), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n308), .B2(new_n297), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT102), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n295), .B(new_n310), .C1(new_n311), .C2(KEYINPUT17), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n294), .ZN(new_n313));
  INV_X1    g112(.A(new_n286), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT17), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT102), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n312), .B1(new_n319), .B2(new_n310), .ZN(new_n320));
  NAND2_X1  g119(.A1(G232gat), .A2(G233gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT99), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT41), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n266), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G190gat), .B(G218gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n265), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n312), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n311), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n310), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT103), .B1(new_n335), .B2(new_n324), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n266), .A3(new_n325), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n327), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n339));
  XOR2_X1   g138(.A(G134gat), .B(G162gat), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n329), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n329), .B2(new_n338), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G141gat), .B(G148gat), .Z(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  INV_X1    g145(.A(G162gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(KEYINPUT2), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G141gat), .B(G148gat), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n349), .B(new_n348), .C1(new_n353), .C2(KEYINPUT2), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT74), .B1(new_n355), .B2(KEYINPUT3), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n352), .A2(new_n354), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G127gat), .B(G134gat), .Z(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G113gat), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n366), .B2(new_n367), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n361), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n361), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(KEYINPUT70), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n364), .A3(G120gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n363), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(new_n377), .A3(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n355), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n372), .A3(new_n378), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n363), .A2(new_n365), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT1), .B1(new_n387), .B2(KEYINPUT69), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n373), .B1(new_n388), .B2(new_n368), .ZN(new_n389));
  INV_X1    g188(.A(new_n378), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n381), .A2(new_n382), .A3(new_n386), .A4(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n355), .B1(new_n389), .B2(new_n390), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n382), .B1(new_n394), .B2(new_n384), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT5), .B1(new_n395), .B2(KEYINPUT75), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT75), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n397), .B(new_n382), .C1(new_n394), .C2(new_n384), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n393), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n392), .A2(new_n386), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(KEYINPUT5), .A3(new_n382), .A4(new_n381), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n381), .ZN(new_n409));
  INV_X1    g208(.A(new_n382), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n382), .A3(new_n384), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT39), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n382), .B1(new_n400), .B2(new_n381), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT39), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n406), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT40), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT83), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n420), .A3(KEYINPUT40), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n408), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n417), .A2(KEYINPUT40), .ZN(new_n423));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(new_n203), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(new_n300), .ZN(new_n426));
  AND2_X1   g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT67), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT66), .ZN(new_n430));
  AND2_X1   g229(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT27), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n245), .ZN(new_n435));
  NAND2_X1  g234(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT66), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G190gat), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI211_X1 g239(.A(KEYINPUT28), .B(G190gat), .C1(new_n435), .C2(new_n436), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n428), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G169gat), .ZN(new_n443));
  INV_X1    g242(.A(G176gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT68), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT26), .Z(new_n446));
  NAND2_X1  g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT65), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n446), .A2(new_n448), .B1(G183gat), .B2(G190gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n441), .ZN(new_n450));
  AOI21_X1  g249(.A(G190gat), .B1(new_n433), .B2(new_n437), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n450), .B(KEYINPUT67), .C1(new_n451), .C2(new_n429), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n442), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT73), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR3_X1   g255(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n448), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n459), .A2(KEYINPUT64), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(KEYINPUT64), .ZN(new_n461));
  NAND3_X1  g260(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(G183gat), .B2(G190gat), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT25), .B1(new_n463), .B2(new_n459), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n465), .A2(KEYINPUT25), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n453), .A2(new_n454), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n454), .B1(new_n453), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n427), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT72), .B(KEYINPUT22), .Z(new_n471));
  NAND2_X1  g270(.A1(G211gat), .A2(G218gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G218gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n223), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n472), .ZN(new_n476));
  XNOR2_X1  g275(.A(G197gat), .B(G204gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n472), .B(new_n475), .C1(new_n479), .C2(new_n471), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n453), .A2(new_n467), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n427), .A2(KEYINPUT29), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n470), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(KEYINPUT73), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n453), .A2(new_n454), .A3(new_n467), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n484), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n453), .A2(new_n467), .A3(new_n427), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n482), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n426), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n481), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n482), .A3(new_n485), .ZN(new_n495));
  INV_X1    g294(.A(new_n426), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n497), .A3(KEYINPUT30), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n494), .A2(new_n499), .A3(new_n495), .A4(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n422), .A2(new_n423), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(G50gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G78gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(G106gat), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT82), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n360), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(KEYINPUT79), .A3(new_n482), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT29), .B1(new_n478), .B2(new_n480), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(KEYINPUT78), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n358), .B1(new_n512), .B2(KEYINPUT78), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n355), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT29), .B1(new_n356), .B2(new_n359), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n481), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G228gat), .A2(G233gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G22gat), .ZN(new_n522));
  OR3_X1    g321(.A1(new_n517), .A2(KEYINPUT81), .A3(new_n481), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n512), .A2(KEYINPUT80), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n358), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n512), .A2(KEYINPUT80), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n355), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n520), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT81), .B1(new_n517), .B2(new_n481), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n523), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n521), .A2(new_n522), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n522), .B1(new_n521), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n508), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n521), .A2(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G22gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n521), .A2(new_n522), .A3(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n507), .B(KEYINPUT82), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n493), .A2(new_n482), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n470), .A2(new_n481), .A3(new_n485), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT37), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n494), .A2(new_n544), .A3(new_n495), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT38), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n543), .A2(new_n545), .A3(new_n546), .A4(new_n426), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n547), .A2(KEYINPUT84), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n426), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n544), .B1(new_n494), .B2(new_n495), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT38), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(KEYINPUT84), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n399), .A2(new_n401), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n405), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT6), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n407), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n408), .A2(KEYINPUT6), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n497), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n503), .B(new_n540), .C1(new_n553), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT76), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n561), .A3(new_n556), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n406), .B1(new_n399), .B2(new_n401), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT76), .B1(new_n563), .B2(KEYINPUT6), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n564), .A3(new_n407), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n558), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n501), .ZN(new_n567));
  INV_X1    g366(.A(new_n540), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n483), .A2(new_n391), .ZN(new_n569));
  NAND2_X1  g368(.A1(G227gat), .A2(G233gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n453), .A2(new_n379), .A3(new_n467), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT32), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G15gat), .B(G43gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G99gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n573), .B(KEYINPUT32), .C1(new_n575), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n569), .A2(new_n572), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n570), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT34), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n453), .A2(new_n379), .A3(new_n467), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n379), .B1(new_n453), .B2(new_n467), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n587), .B(new_n570), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT71), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n584), .A2(new_n592), .A3(new_n587), .A4(new_n570), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n586), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n583), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n591), .A2(new_n593), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(new_n582), .A3(new_n580), .A4(new_n586), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n597), .A3(KEYINPUT36), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n597), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n567), .A2(new_n568), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n560), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n595), .A2(new_n597), .A3(KEYINPUT85), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT85), .B1(new_n595), .B2(new_n597), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT35), .B1(new_n557), .B2(new_n558), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n501), .A2(new_n540), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT86), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n540), .A2(new_n595), .A3(new_n597), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT35), .B1(new_n567), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n501), .A2(new_n540), .A3(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT86), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT85), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n583), .A2(new_n594), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n596), .A2(new_n586), .B1(new_n580), .B2(new_n582), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n595), .A2(new_n597), .A3(KEYINPUT85), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n609), .A2(new_n611), .A3(new_n620), .ZN(new_n621));
  AOI211_X1 g420(.A(new_n264), .B(new_n344), .C1(new_n603), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n237), .A2(new_n239), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n331), .B2(new_n332), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n242), .A2(new_n315), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(KEYINPUT18), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n244), .A2(new_n295), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n626), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n627), .B(KEYINPUT13), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n630), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT11), .B(G169gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G197gat), .ZN(new_n640));
  XOR2_X1   g439(.A(G113gat), .B(G141gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT87), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n645), .A3(new_n635), .A4(new_n637), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n648), .A2(KEYINPUT94), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(KEYINPUT94), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n305), .A2(KEYINPUT104), .ZN(new_n655));
  OAI22_X1  g454(.A1(new_n307), .A2(new_n309), .B1(new_n225), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n225), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n308), .A2(new_n305), .A3(new_n297), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n304), .A2(new_n306), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n229), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n654), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n660), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n654), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT106), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n362), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n662), .A2(KEYINPUT105), .A3(new_n663), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT105), .B1(new_n662), .B2(new_n663), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n653), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n665), .A2(new_n654), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n675), .A3(new_n670), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n652), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n622), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n566), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n232), .ZN(G1324gat));
  OAI21_X1  g480(.A(G8gat), .B1(new_n679), .B2(new_n501), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT16), .B(G8gat), .Z(new_n683));
  NAND4_X1  g482(.A1(new_n622), .A2(new_n678), .A3(new_n502), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT107), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n685), .A2(new_n689), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n679), .ZN(new_n692));
  INV_X1    g491(.A(new_n601), .ZN(new_n693));
  INV_X1    g492(.A(new_n598), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n692), .A2(G15gat), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(G15gat), .B1(new_n692), .B2(new_n619), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n679), .A2(new_n540), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n621), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n609), .A2(new_n620), .A3(new_n611), .A4(KEYINPUT108), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n603), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n344), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n344), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n603), .B2(new_n621), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT44), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n678), .A2(new_n264), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n566), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n710), .A2(new_n715), .ZN(new_n718));
  INV_X1    g517(.A(new_n566), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(new_n280), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(G1328gat));
  NAND2_X1  g521(.A1(new_n275), .A2(new_n276), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n723), .A3(new_n502), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT46), .Z(new_n725));
  NOR2_X1   g524(.A1(new_n716), .A2(new_n501), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n723), .ZN(G1329gat));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  AOI21_X1  g527(.A(G43gat), .B1(new_n718), .B2(new_n619), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n695), .A2(G43gat), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n728), .B(new_n730), .C1(new_n716), .C2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n712), .A2(new_n714), .A3(new_n731), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT47), .B1(new_n733), .B2(new_n729), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1330gat));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  AOI21_X1  g535(.A(G50gat), .B1(new_n718), .B2(new_n568), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n568), .A2(G50gat), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n736), .B(new_n738), .C1(new_n716), .C2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n712), .A2(new_n714), .A3(new_n739), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT48), .B1(new_n741), .B2(new_n737), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1331gat));
  NOR2_X1   g542(.A1(new_n264), .A2(new_n344), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n705), .A2(new_n652), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n677), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n566), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n202), .ZN(G1332gat));
  NAND2_X1  g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n502), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n746), .A2(KEYINPUT109), .A3(new_n750), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n752), .A2(new_n753), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n753), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n751), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1333gat));
  AND2_X1   g557(.A1(new_n745), .A2(new_n677), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(G71gat), .A3(new_n695), .ZN(new_n760));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n746), .B2(new_n606), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT50), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n760), .A2(new_n765), .A3(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n759), .A2(new_n568), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g568(.A1(new_n261), .A2(new_n263), .ZN(new_n770));
  INV_X1    g569(.A(new_n677), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n770), .A2(new_n651), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n708), .A2(new_n719), .A3(new_n711), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(G85gat), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n770), .A2(new_n651), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n705), .A2(new_n344), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n344), .A4(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n782), .A2(new_n299), .A3(new_n719), .A4(new_n677), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n776), .A2(new_n783), .ZN(G1336gat));
  NAND4_X1  g583(.A1(new_n708), .A2(new_n502), .A3(new_n711), .A4(new_n772), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n502), .A2(new_n300), .A3(new_n677), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT52), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n786), .A2(new_n790), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1337gat));
  NAND3_X1  g594(.A1(new_n713), .A2(new_n695), .A3(new_n772), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G99gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n606), .A2(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n677), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1338gat));
  NAND4_X1  g599(.A1(new_n708), .A2(new_n568), .A3(new_n711), .A4(new_n772), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n540), .A2(new_n771), .A3(G106gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT114), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n782), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n802), .B(new_n805), .C1(new_n807), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n502), .A2(new_n566), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n662), .A2(new_n654), .A3(new_n663), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n674), .A2(KEYINPUT54), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n670), .B1(new_n664), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  INV_X1    g620(.A(new_n676), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n651), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n633), .A2(new_n634), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n627), .B1(new_n625), .B2(new_n626), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n642), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT115), .B(new_n642), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n677), .B(new_n831), .C1(new_n649), .C2(new_n650), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n344), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n329), .A2(new_n338), .A3(new_n341), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n631), .A2(new_n637), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT94), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n645), .A4(new_n635), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n648), .A2(KEYINPUT94), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(new_n838), .B1(new_n829), .B2(new_n830), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n329), .A2(new_n338), .ZN(new_n840));
  INV_X1    g639(.A(new_n341), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND4_X1   g641(.A1(new_n834), .A2(new_n839), .A3(new_n823), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n815), .B1(new_n833), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n344), .A2(new_n823), .A3(new_n839), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n651), .A2(new_n823), .B1(new_n839), .B2(new_n677), .ZN(new_n846));
  OAI211_X1 g645(.A(KEYINPUT116), .B(new_n845), .C1(new_n846), .C2(new_n344), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n264), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n770), .A2(new_n709), .A3(new_n652), .A4(new_n771), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n814), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n610), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n364), .A3(new_n651), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n540), .A3(new_n619), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n652), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT117), .ZN(G1340gat));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n362), .A3(new_n677), .ZN(new_n859));
  OAI21_X1  g658(.A(G120gat), .B1(new_n855), .B2(new_n771), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  AOI21_X1  g660(.A(G127gat), .B1(new_n853), .B2(new_n770), .ZN(new_n862));
  INV_X1    g661(.A(G127gat), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n855), .A2(new_n863), .A3(new_n264), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n862), .A2(new_n864), .ZN(G1342gat));
  NOR3_X1   g664(.A1(new_n852), .A2(G134gat), .A3(new_n709), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n855), .B2(new_n709), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n867), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G1343gat));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n695), .A2(new_n540), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n850), .A2(new_n873), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n874), .A2(G141gat), .A3(new_n652), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(KEYINPUT118), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n540), .B1(new_n848), .B2(new_n849), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n695), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n813), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n833), .A2(new_n843), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n849), .B1(new_n882), .B2(new_n770), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n568), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n884), .B2(KEYINPUT57), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n652), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n875), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n876), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n887), .B(new_n875), .C1(KEYINPUT118), .C2(new_n872), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(new_n874), .ZN(new_n892));
  INV_X1    g691(.A(G148gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n677), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n885), .A3(new_n677), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n893), .A2(KEYINPUT59), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n877), .A2(new_n878), .ZN(new_n902));
  INV_X1    g701(.A(new_n881), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n849), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n744), .A2(KEYINPUT120), .A3(new_n652), .A4(new_n771), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n905), .B(new_n906), .C1(new_n882), .C2(new_n770), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n878), .A3(new_n568), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n902), .A2(new_n677), .A3(new_n903), .A4(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n901), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n894), .B1(new_n900), .B2(new_n910), .ZN(G1345gat));
  NOR3_X1   g710(.A1(new_n886), .A2(new_n346), .A3(new_n264), .ZN(new_n912));
  AOI21_X1  g711(.A(G155gat), .B1(new_n892), .B2(new_n770), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(G1346gat));
  NOR3_X1   g713(.A1(new_n886), .A2(new_n347), .A3(new_n709), .ZN(new_n915));
  AOI21_X1  g714(.A(G162gat), .B1(new_n892), .B2(new_n344), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1347gat));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n848), .A2(new_n849), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n566), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n922), .A3(new_n566), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n610), .A2(new_n501), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n924), .A2(new_n443), .A3(new_n651), .A4(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n719), .A2(new_n501), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n606), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n848), .B2(new_n849), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n568), .B1(new_n929), .B2(new_n930), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n652), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n918), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n922), .B1(new_n919), .B2(new_n566), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT121), .B(new_n719), .C1(new_n848), .C2(new_n849), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n443), .B(new_n925), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n918), .B(new_n935), .C1(new_n939), .C2(new_n652), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n936), .A2(new_n941), .ZN(G1348gat));
  OAI211_X1 g741(.A(new_n677), .B(new_n925), .C1(new_n937), .C2(new_n938), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(new_n444), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n932), .A2(G176gat), .A3(new_n677), .A4(new_n933), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT125), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n943), .A2(new_n444), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n951), .A2(new_n952), .A3(new_n948), .A4(new_n947), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(G1349gat));
  NAND4_X1  g753(.A1(new_n924), .A2(new_n438), .A3(new_n770), .A4(new_n925), .ZN(new_n955));
  OAI21_X1  g754(.A(G183gat), .B1(new_n934), .B2(new_n264), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n959), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n932), .A2(new_n344), .A3(new_n933), .ZN(new_n962));
  NAND2_X1  g761(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n962), .A2(G190gat), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g763(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n924), .A2(new_n439), .A3(new_n925), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n966), .B(new_n967), .C1(new_n709), .C2(new_n968), .ZN(G1351gat));
  NOR2_X1   g768(.A1(new_n928), .A2(new_n695), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n902), .A2(new_n908), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n652), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n937), .A2(new_n938), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n873), .A2(new_n502), .ZN(new_n974));
  OR3_X1    g773(.A1(new_n973), .A2(G197gat), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n975), .B2(new_n652), .ZN(G1352gat));
  NOR2_X1   g775(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  XOR2_X1   g776(.A(KEYINPUT127), .B(G204gat), .Z(new_n978));
  NOR2_X1   g777(.A1(new_n771), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n902), .A2(new_n677), .A3(new_n908), .ZN(new_n982));
  INV_X1    g781(.A(new_n970), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n977), .A2(new_n985), .A3(new_n979), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n981), .A2(new_n984), .A3(new_n986), .ZN(G1353gat));
  NAND3_X1  g786(.A1(new_n977), .A2(new_n223), .A3(new_n770), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n902), .A2(new_n770), .A3(new_n908), .A4(new_n970), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  AOI21_X1  g792(.A(G218gat), .B1(new_n977), .B2(new_n344), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n971), .A2(new_n474), .A3(new_n709), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


