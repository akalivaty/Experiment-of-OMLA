//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G77), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT65), .B(G244), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n218), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n215), .B1(new_n209), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n216), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n248), .A2(new_n249), .B1(new_n216), .B2(G68), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n216), .A2(new_n246), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n250), .A2(KEYINPUT80), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n250), .A2(KEYINPUT80), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n247), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT11), .Z(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n260), .A2(new_n257), .A3(G13), .A4(G20), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT74), .B1(new_n259), .B2(new_n261), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n266));
  INV_X1    g0066(.A(new_n247), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n257), .A2(G20), .ZN(new_n268));
  XOR2_X1   g0068(.A(new_n268), .B(KEYINPUT69), .Z(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n264), .A2(G68), .A3(new_n267), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n259), .A2(new_n261), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G68), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n266), .B(new_n271), .C1(KEYINPUT12), .C2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n256), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT81), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT78), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G97), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  AND2_X1   g0087(.A1(G232), .A2(G1698), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT78), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n287), .A2(new_n290), .A3(G226), .A4(new_n282), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n284), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT79), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT79), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n292), .A2(new_n298), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  INV_X1    g0101(.A(new_n215), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n293), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(KEYINPUT66), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT66), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n257), .C1(G41), .C2(G45), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n308), .A2(new_n294), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(G238), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n278), .B1(new_n300), .B2(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n292), .A2(new_n298), .A3(new_n295), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n298), .B1(new_n292), .B2(new_n295), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n278), .B(new_n312), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n277), .B(G169), .C1(new_n313), .C2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(G179), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n316), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n277), .B1(new_n323), .B2(G169), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n276), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(G169), .B1(new_n313), .B2(new_n317), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n321), .A4(new_n318), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n275), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n275), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n320), .B2(new_n316), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n269), .A2(new_n251), .ZN(new_n337));
  INV_X1    g0137(.A(new_n272), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n247), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n337), .A2(new_n339), .B1(new_n251), .B2(new_n338), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n341), .A2(new_n248), .B1(new_n342), .B2(new_n252), .ZN(new_n343));
  INV_X1    g0143(.A(new_n203), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n216), .B1(new_n344), .B2(new_n251), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n247), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT67), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n347), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n340), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT9), .ZN(new_n351));
  OR2_X1    g0151(.A1(KEYINPUT3), .A2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  AOI21_X1  g0153(.A(G1698), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G222), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n282), .B1(new_n352), .B2(new_n353), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G223), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n355), .B(new_n357), .C1(new_n219), .C2(new_n287), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n295), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n307), .B1(new_n311), .B2(G226), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G190), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT75), .B(G200), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n361), .A2(new_n365), .B1(new_n366), .B2(KEYINPUT10), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n351), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(KEYINPUT10), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n361), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n350), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n308), .A2(new_n221), .A3(new_n294), .A4(new_n310), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT70), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n306), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n306), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT70), .ZN(new_n381));
  OAI211_X1 g0181(.A(G238), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n206), .B2(new_n287), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n287), .A2(new_n384), .A3(G232), .A4(new_n282), .ZN(new_n385));
  OAI211_X1 g0185(.A(G232), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT71), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n383), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n379), .B(new_n381), .C1(new_n388), .C2(new_n294), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT72), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n377), .B2(new_n306), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n356), .A2(G238), .B1(new_n281), .B2(G107), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n384), .B1(new_n354), .B2(G232), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n386), .A2(KEYINPUT71), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(new_n295), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT72), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n379), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n390), .A2(new_n398), .A3(new_n373), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT76), .ZN(new_n400));
  AOI21_X1  g0200(.A(G179), .B1(new_n390), .B2(new_n398), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n216), .A2(new_n219), .B1(new_n341), .B2(new_n252), .ZN(new_n404));
  INV_X1    g0204(.A(new_n248), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT15), .B(G87), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n404), .A2(KEYINPUT73), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(KEYINPUT73), .B2(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n247), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n264), .A2(G77), .A3(new_n267), .A4(new_n270), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n265), .A2(new_n219), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n401), .B2(KEYINPUT76), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n403), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n397), .B1(new_n396), .B2(new_n379), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n387), .A2(new_n385), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n294), .B1(new_n418), .B2(new_n392), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n377), .A2(new_n378), .A3(new_n306), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n419), .A2(new_n420), .A3(new_n391), .A4(KEYINPUT72), .ZN(new_n421));
  OAI21_X1  g0221(.A(G190), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n390), .A2(new_n398), .A3(new_n365), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n414), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n287), .A2(new_n427), .A3(G20), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n281), .B2(new_n216), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G58), .A2(G68), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n203), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G20), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT82), .ZN(new_n434));
  INV_X1    g0234(.A(new_n252), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G159), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n216), .B1(new_n203), .B2(new_n431), .ZN(new_n438));
  INV_X1    g0238(.A(G159), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n252), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT82), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n430), .A2(KEYINPUT16), .A3(new_n437), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT16), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n427), .B1(new_n287), .B2(G20), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n202), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n433), .A2(new_n436), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(new_n247), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n308), .A2(G232), .A3(new_n294), .A4(new_n310), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n450), .A2(new_n306), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G87), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT84), .ZN(new_n453));
  OAI211_X1 g0253(.A(G223), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n454));
  OAI211_X1 g0254(.A(G226), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n295), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G190), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n269), .A2(new_n341), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(new_n339), .B1(new_n338), .B2(new_n341), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n451), .A2(new_n457), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G200), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n449), .A2(new_n459), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT87), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n461), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n437), .A2(new_n441), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n446), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n267), .B1(new_n469), .B2(KEYINPUT16), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n467), .B1(new_n470), .B2(new_n448), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n462), .A2(new_n330), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(G200), .B2(new_n462), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT87), .ZN(new_n474));
  INV_X1    g0274(.A(new_n465), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n471), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n464), .A2(KEYINPUT17), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n466), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n449), .A2(new_n461), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT83), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n449), .A2(KEYINPUT83), .A3(new_n461), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n458), .A2(G179), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n462), .A2(G169), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g0285(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n486));
  NAND4_X1  g0286(.A1(new_n481), .A2(new_n482), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n449), .A2(KEYINPUT83), .A3(new_n461), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT83), .B1(new_n449), .B2(new_n461), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n483), .A2(new_n484), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n478), .B(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AND4_X1   g0294(.A1(new_n336), .A2(new_n376), .A3(new_n426), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT91), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(KEYINPUT21), .ZN(new_n497));
  OAI211_X1 g0297(.A(G264), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT90), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n287), .A2(KEYINPUT90), .A3(G264), .A4(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G257), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n352), .B2(new_n353), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(new_n282), .B1(new_n281), .B2(G303), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n294), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT88), .ZN(new_n507));
  INV_X1    g0307(.A(G41), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n509));
  INV_X1    g0309(.A(G45), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G1), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT5), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT88), .B1(new_n512), .B2(G41), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(G41), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n509), .B(new_n511), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(G270), .A3(new_n294), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n507), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n512), .B2(G41), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n257), .A2(G45), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n514), .B2(new_n507), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n520), .A3(new_n303), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(G169), .B1(new_n506), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n272), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n261), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n257), .B2(G33), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n267), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n262), .B2(new_n263), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n216), .C1(G33), .C2(new_n205), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n247), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n532), .A2(new_n247), .A3(KEYINPUT20), .A4(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n529), .A2(new_n530), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n497), .B1(new_n523), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n522), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n542));
  INV_X1    g0342(.A(G303), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n287), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n500), .B2(new_n501), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n541), .B(G190), .C1(new_n545), .C2(new_n294), .ZN(new_n546));
  OAI21_X1  g0346(.A(G200), .B1(new_n506), .B2(new_n522), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(new_n539), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n541), .B1(new_n545), .B2(new_n294), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n529), .A2(new_n530), .A3(new_n538), .ZN(new_n550));
  INV_X1    g0350(.A(new_n497), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n549), .A2(G169), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n506), .A2(new_n371), .A3(new_n522), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n550), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n540), .A2(new_n548), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G250), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n556));
  OAI211_X1 g0356(.A(G244), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n531), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT4), .B1(new_n354), .B2(G244), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n295), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n295), .B1(new_n518), .B2(new_n520), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G257), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n521), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n338), .A2(new_n205), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n257), .A2(G33), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n272), .A2(new_n267), .A3(G97), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g0369(.A(G97), .B(G107), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT6), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n571), .A2(new_n205), .A3(G107), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(G20), .B1(G77), .B2(new_n435), .ZN(new_n576));
  OAI21_X1  g0376(.A(G107), .B1(new_n428), .B2(new_n429), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n569), .B1(new_n578), .B2(new_n247), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n561), .A2(G190), .A3(new_n521), .A4(new_n563), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n565), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n216), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT22), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n287), .A2(new_n584), .A3(new_n216), .A4(G87), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT23), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n216), .B2(G107), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n405), .A2(G116), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n587), .B1(new_n586), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n247), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n338), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT25), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n272), .B2(G107), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n272), .A2(G107), .A3(new_n267), .A4(new_n567), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(G257), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n601));
  OAI211_X1 g0401(.A(G250), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n602));
  INV_X1    g0402(.A(G294), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n601), .B(new_n602), .C1(new_n246), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n295), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n515), .A2(G264), .A3(new_n294), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n521), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G200), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(G190), .A3(new_n521), .A4(new_n606), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n594), .A2(new_n600), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n564), .A2(new_n373), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n561), .A2(new_n371), .A3(new_n521), .A4(new_n563), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n573), .B1(new_n571), .B2(new_n570), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n613), .A2(new_n216), .B1(new_n249), .B2(new_n252), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n206), .B1(new_n444), .B2(new_n445), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n247), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n569), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n581), .A2(new_n610), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n607), .A2(new_n373), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n605), .A2(new_n371), .A3(new_n521), .A4(new_n606), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n594), .B2(new_n600), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n406), .B1(new_n262), .B2(new_n263), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT19), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n216), .B1(new_n285), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G87), .B2(new_n207), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n216), .B(G68), .C1(new_n279), .C2(new_n280), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n626), .B1(new_n248), .B2(new_n205), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n247), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n272), .A2(new_n267), .A3(G87), .A4(new_n567), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n625), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(G238), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n635));
  OAI211_X1 g0435(.A(G244), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n636));
  NAND2_X1  g0436(.A1(G33), .A2(G116), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n295), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n294), .A2(G274), .A3(new_n511), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n294), .A2(G250), .A3(new_n519), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(G190), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n642), .B1(new_n295), .B2(new_n638), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(KEYINPUT89), .A3(G190), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n639), .A2(new_n643), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n365), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n634), .A2(new_n646), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n272), .A2(new_n267), .A3(new_n407), .A4(new_n567), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n625), .A2(new_n632), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n371), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n653), .B(new_n654), .C1(G169), .C2(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n620), .A2(new_n624), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n495), .A2(new_n555), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT92), .ZN(G372));
  NAND2_X1  g0459(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT93), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n647), .B2(G169), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n649), .A2(KEYINPUT93), .A3(new_n373), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n634), .A2(new_n644), .A3(new_n650), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n664), .A2(new_n619), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n581), .A2(new_n610), .A3(new_n619), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n586), .A2(new_n591), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT24), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n267), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n598), .A2(new_n599), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n621), .B(new_n622), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(new_n540), .A3(new_n554), .A4(new_n552), .ZN(new_n676));
  INV_X1    g0476(.A(new_n660), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n663), .A2(new_n662), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n625), .A2(new_n632), .A3(new_n633), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n364), .B1(new_n639), .B2(new_n643), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n677), .A2(new_n678), .B1(new_n681), .B2(new_n644), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n669), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT26), .B1(new_n656), .B2(new_n619), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n668), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n495), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n375), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n479), .A2(new_n485), .ZN(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n416), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n329), .B1(new_n334), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n466), .A2(new_n476), .A3(new_n477), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n687), .B1(new_n696), .B2(new_n370), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n686), .A2(new_n697), .ZN(G369));
  NAND3_X1  g0498(.A1(new_n257), .A2(new_n216), .A3(G13), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n550), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n555), .A2(new_n705), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n540), .A2(new_n554), .A3(new_n552), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n675), .A2(new_n704), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n704), .B1(new_n673), .B2(new_n674), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n610), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n711), .B1(new_n675), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n707), .A2(new_n704), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n711), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n210), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n213), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n624), .A2(new_n656), .ZN(new_n726));
  INV_X1    g0526(.A(new_n704), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n669), .A3(new_n555), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT96), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT96), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n657), .A2(new_n730), .A3(new_n555), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n607), .A2(new_n649), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n354), .A2(KEYINPUT4), .A3(G244), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n557), .A2(new_n558), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n531), .A4(new_n556), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n736), .A2(new_n295), .B1(G257), .B2(new_n562), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n733), .A2(new_n553), .A3(KEYINPUT30), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n561), .A2(new_n563), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n607), .A3(new_n649), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT95), .A3(KEYINPUT30), .A4(new_n553), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n604), .A2(new_n295), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n606), .A2(new_n521), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n737), .A3(new_n647), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n541), .B(G179), .C1(new_n545), .C2(new_n294), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n747), .A2(G179), .A3(new_n647), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n549), .A3(new_n564), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n740), .A2(new_n743), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n704), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT31), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n732), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n758), .A2(G330), .ZN(new_n759));
  INV_X1    g0559(.A(new_n683), .ZN(new_n760));
  INV_X1    g0560(.A(new_n664), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(new_n667), .A3(new_n655), .A4(new_n651), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n761), .B(new_n763), .C1(new_n666), .C2(new_n667), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n727), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT29), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n682), .A2(new_n762), .A3(new_n667), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n767), .A2(new_n684), .A3(new_n761), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n704), .B1(new_n768), .B2(new_n683), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n766), .B1(new_n770), .B2(KEYINPUT29), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n759), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n725), .B1(new_n772), .B2(G1), .ZN(G364));
  NOR2_X1   g0573(.A1(new_n708), .A2(G330), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT97), .Z(new_n775));
  AND2_X1   g0575(.A1(new_n216), .A2(G13), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n257), .B1(new_n776), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n720), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n775), .A2(new_n709), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n719), .A2(new_n281), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G355), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G116), .B2(new_n210), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n241), .A2(new_n510), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n719), .A2(new_n287), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n510), .B2(new_n214), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n215), .B1(G20), .B2(new_n373), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n779), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n216), .A2(new_n371), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G190), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n287), .B1(new_n799), .B2(new_n219), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n797), .A2(G190), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT32), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n216), .A2(G179), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n798), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n439), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n803), .A2(new_n201), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n797), .A2(new_n330), .A3(G200), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n800), .B(new_n808), .C1(G68), .C2(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n330), .A2(G179), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n216), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n205), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n801), .A2(new_n332), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n251), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n814), .B(new_n817), .C1(new_n804), .C2(new_n807), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n365), .A2(new_n805), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n330), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(G190), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G87), .A2(new_n820), .B1(new_n821), .B2(G107), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n811), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT98), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G326), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n816), .A2(new_n826), .B1(new_n603), .B2(new_n813), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G322), .B2(new_n802), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n281), .B1(new_n799), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(KEYINPUT33), .B(G317), .Z(new_n831));
  INV_X1    g0631(.A(G329), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n809), .A2(new_n831), .B1(new_n832), .B2(new_n806), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n830), .B(new_n833), .C1(new_n821), .C2(G283), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n820), .B(KEYINPUT99), .Z(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n828), .B(new_n834), .C1(new_n836), .C2(new_n543), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n823), .A2(new_n824), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n825), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n796), .B1(new_n839), .B2(new_n793), .ZN(new_n840));
  INV_X1    g0640(.A(new_n792), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n708), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n781), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  NOR2_X1   g0644(.A1(new_n793), .A2(new_n790), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n779), .B1(G77), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n803), .A2(new_n603), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n814), .B(new_n848), .C1(G303), .C2(new_n815), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n281), .B1(new_n809), .B2(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n799), .A2(new_n527), .B1(new_n806), .B2(new_n829), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(new_n821), .C2(G87), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n849), .B(new_n853), .C1(new_n836), .C2(new_n206), .ZN(new_n854));
  INV_X1    g0654(.A(new_n799), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n810), .A2(G150), .B1(new_n855), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G143), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n803), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G137), .B2(new_n815), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n287), .B1(new_n806), .B2(new_n861), .C1(new_n813), .C2(new_n201), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G68), .B2(new_n821), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n836), .B2(new_n251), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n854), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n847), .B1(new_n865), .B2(new_n793), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n413), .A2(new_n704), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n390), .A2(new_n398), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n399), .A2(KEYINPUT76), .B1(new_n868), .B2(new_n371), .ZN(new_n869));
  OAI211_X1 g0669(.A(KEYINPUT76), .B(new_n371), .C1(new_n417), .C2(new_n421), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n413), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n424), .B(new_n867), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n867), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n403), .A2(new_n415), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n866), .B1(new_n875), .B2(new_n791), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT100), .Z(new_n877));
  INV_X1    g0677(.A(new_n759), .ZN(new_n878));
  INV_X1    g0678(.A(new_n875), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(new_n769), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n779), .B1(new_n878), .B2(new_n881), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(G384));
  AND2_X1   g0686(.A1(new_n729), .A2(new_n731), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n757), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n753), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n704), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n756), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT106), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n756), .A2(new_n890), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT106), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(new_n732), .A3(new_n894), .A4(new_n889), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n325), .A2(new_n328), .ZN(new_n897));
  INV_X1    g0697(.A(new_n275), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n275), .A2(new_n727), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n334), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT102), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n325), .A2(new_n328), .A3(new_n334), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n900), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n899), .A2(new_n903), .A3(new_n334), .A4(new_n901), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n896), .A2(new_n906), .A3(new_n875), .A4(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n464), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n491), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n702), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n481), .A2(new_n482), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n464), .A3(new_n688), .ZN(new_n915));
  INV_X1    g0715(.A(new_n910), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n912), .A2(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n692), .B2(new_n478), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n909), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n443), .B1(new_n468), .B2(new_n446), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n467), .B1(new_n470), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n702), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(new_n695), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n481), .A2(new_n482), .A3(new_n485), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n925), .A2(new_n914), .A3(new_n464), .A4(new_n910), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n464), .B1(new_n921), .B2(new_n490), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT37), .B1(new_n927), .B2(new_n922), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n919), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT40), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n908), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n924), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n924), .B2(new_n929), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n908), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n495), .A2(new_n896), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  INV_X1    g0743(.A(G330), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n495), .A2(new_n771), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n697), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT104), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n416), .A2(new_n704), .ZN(new_n949));
  AOI211_X1 g0749(.A(KEYINPUT101), .B(new_n949), .C1(new_n769), .C2(new_n875), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT101), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n875), .A2(new_n685), .A3(new_n727), .ZN(new_n952));
  INV_X1    g0752(.A(new_n949), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n906), .B(new_n907), .C1(new_n950), .C2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n937), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT39), .B1(new_n919), .B2(new_n930), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n937), .B2(KEYINPUT39), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n329), .A3(new_n727), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n702), .B1(new_n690), .B2(new_n691), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n948), .B(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n945), .A2(new_n962), .B1(new_n257), .B2(new_n776), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n945), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n965), .A2(G116), .A3(new_n217), .A4(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT36), .Z(new_n968));
  NAND3_X1  g0768(.A1(new_n214), .A2(new_n220), .A3(new_n431), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n251), .A2(G68), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n257), .B(G13), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n964), .A2(new_n968), .A3(new_n971), .ZN(G367));
  NAND2_X1  g0772(.A1(new_n679), .A2(new_n704), .ZN(new_n973));
  MUX2_X1   g0773(.A(new_n664), .B(new_n682), .S(new_n973), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n581), .B(new_n619), .C1(new_n579), .C2(new_n727), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n619), .B2(new_n727), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n714), .A2(new_n716), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n619), .B1(new_n976), .B2(new_n675), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n727), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n975), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n984), .B(new_n985), .Z(new_n986));
  INV_X1    g0786(.A(new_n715), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n977), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT107), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n988), .B(KEYINPUT107), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n720), .B(KEYINPUT41), .Z(new_n993));
  NAND2_X1  g0793(.A1(new_n717), .A2(new_n977), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT45), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n717), .A2(new_n977), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(new_n987), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT109), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n709), .B2(KEYINPUT108), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n1000), .B2(new_n709), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n714), .B(new_n716), .Z(new_n1003));
  MUX2_X1   g0803(.A(new_n1001), .B(new_n1002), .S(new_n1003), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n772), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n999), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n993), .B1(new_n1006), .B2(new_n772), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n991), .B1(new_n986), .B2(new_n992), .C1(new_n1007), .C2(new_n778), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n794), .B1(new_n210), .B2(new_n406), .C1(new_n237), .C2(new_n787), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1009), .A2(new_n779), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n857), .A2(new_n816), .B1(new_n803), .B2(new_n342), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n813), .A2(new_n202), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n809), .A2(new_n439), .B1(new_n799), .B2(new_n251), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n806), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n281), .B(new_n1014), .C1(G137), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n820), .A2(G58), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n821), .A2(new_n220), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT46), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n836), .A2(new_n1020), .A3(new_n527), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n543), .A2(new_n803), .B1(new_n816), .B2(new_n829), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n813), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(G107), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n820), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1020), .B1(new_n1025), .B2(new_n527), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n821), .A2(G97), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n809), .A2(new_n603), .B1(new_n799), .B2(new_n850), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n287), .B(new_n1028), .C1(G317), .C2(new_n1015), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1019), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  INV_X1    g0832(.A(new_n793), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1010), .B1(new_n841), .B2(new_n974), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1008), .A2(new_n1034), .ZN(G387));
  NAND2_X1  g0835(.A1(new_n1004), .A2(new_n778), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT110), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n341), .A2(G50), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT50), .Z(new_n1039));
  OAI211_X1 g0839(.A(new_n722), .B(new_n510), .C1(new_n202), .C2(new_n249), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n786), .B1(new_n1039), .B2(new_n1040), .C1(new_n234), .C2(new_n510), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n722), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n782), .A2(new_n1042), .B1(new_n206), .B2(new_n719), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(KEYINPUT111), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n794), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT111), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n779), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n813), .A2(new_n406), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n287), .B1(new_n806), .B2(new_n342), .C1(new_n803), .C2(new_n251), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(G159), .C2(new_n815), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n809), .A2(new_n341), .B1(new_n799), .B2(new_n202), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT112), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n820), .A2(new_n220), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1027), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n810), .A2(G311), .B1(new_n855), .B2(G303), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n802), .A2(G317), .ZN(new_n1056));
  INV_X1    g0856(.A(G322), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1055), .B(new_n1056), .C1(new_n1057), .C2(new_n816), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n820), .A2(G294), .B1(G283), .B2(new_n1023), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT49), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n821), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n281), .B1(new_n826), .B2(new_n806), .C1(new_n1066), .C2(new_n527), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1054), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1047), .B1(new_n1070), .B2(new_n793), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n714), .B2(new_n841), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1004), .A2(new_n772), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n720), .B(KEYINPUT113), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1005), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1037), .B(new_n1072), .C1(new_n1073), .C2(new_n1075), .ZN(G393));
  NAND2_X1  g0876(.A1(new_n999), .A2(new_n1005), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1006), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT114), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n777), .B1(new_n999), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1079), .B2(new_n999), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n794), .B1(new_n205), .B2(new_n210), .C1(new_n244), .C2(new_n787), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n779), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G150), .A2(new_n815), .B1(new_n802), .B2(G159), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n809), .A2(new_n251), .B1(new_n806), .B2(new_n857), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n813), .A2(new_n249), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n287), .B1(new_n799), .B2(new_n341), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G68), .A2(new_n820), .B1(new_n821), .B2(G87), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1086), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1092), .A2(KEYINPUT116), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G311), .A2(new_n802), .B1(new_n815), .B2(G317), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT52), .Z(new_n1095));
  OAI21_X1  g0895(.A(new_n281), .B1(new_n799), .B2(new_n603), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n809), .A2(new_n543), .B1(new_n806), .B2(new_n1057), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(G116), .C2(new_n1023), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G107), .A2(new_n821), .B1(new_n820), .B2(G283), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1092), .A2(KEYINPUT116), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1083), .B1(new_n1102), .B2(new_n793), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n977), .B2(new_n841), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1078), .A2(new_n1081), .A3(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n329), .A2(new_n727), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n958), .B1(new_n955), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n953), .B1(new_n879), .B2(new_n765), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n904), .A2(new_n900), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT102), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n329), .A2(new_n335), .A3(new_n900), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n907), .B(new_n1109), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n931), .A2(new_n1107), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n758), .A2(G330), .A3(new_n875), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n906), .A3(new_n907), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1106), .B1(new_n1108), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n907), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n950), .A2(new_n954), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1107), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n958), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n329), .A2(KEYINPUT102), .A3(new_n335), .A4(new_n900), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n902), .B2(new_n905), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1127), .A2(new_n1117), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(KEYINPUT117), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1125), .A2(new_n1115), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n908), .A2(new_n944), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1120), .A2(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n778), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n780), .B1(new_n341), .B2(new_n845), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1135), .A2(new_n816), .B1(new_n803), .B2(new_n861), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT54), .B(G143), .Z(new_n1137));
  AOI21_X1  g0937(.A(new_n281), .B1(new_n855), .B2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n810), .A2(G137), .B1(new_n1015), .B2(G125), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n1066), .C2(new_n251), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1136), .B(new_n1140), .C1(G159), .C2(new_n1023), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n820), .A2(G150), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT53), .Z(new_n1143));
  OAI22_X1  g0943(.A1(new_n809), .A2(new_n206), .B1(new_n799), .B2(new_n205), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n821), .A2(G68), .B1(new_n1144), .B2(KEYINPUT119), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(KEYINPUT119), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n281), .B1(new_n806), .B2(new_n603), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n527), .A2(new_n803), .B1(new_n816), .B2(new_n850), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1146), .A2(new_n1088), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n835), .A2(G87), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1141), .A2(new_n1143), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1134), .B1(new_n1033), .B2(new_n1151), .C1(new_n958), .C2(new_n791), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1133), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT118), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1115), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1131), .B1(new_n1108), .B2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1108), .A2(new_n1119), .A3(new_n1106), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT117), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1121), .A2(new_n1116), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n908), .B2(new_n944), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1122), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1109), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n944), .B(new_n879), .C1(new_n892), .C2(new_n895), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1118), .B(new_n1164), .C1(new_n1165), .C2(new_n1127), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n495), .A2(G330), .A3(new_n896), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n697), .A3(new_n946), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1154), .B1(new_n1159), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1169), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1132), .A2(KEYINPUT118), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1074), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1159), .B2(new_n1171), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1153), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(G378));
  NOR2_X1   g0979(.A1(G33), .A2(G41), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G50), .B(new_n1180), .C1(new_n281), .C2(new_n508), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n816), .A2(new_n527), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1012), .B(new_n1182), .C1(G107), .C2(new_n802), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n821), .A2(G58), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n809), .A2(new_n205), .B1(new_n799), .B2(new_n406), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n508), .B(new_n281), .C1(new_n806), .C2(new_n850), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1053), .A3(new_n1184), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1181), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1189), .B2(new_n1188), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n810), .A2(G132), .B1(new_n855), .B2(G137), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1135), .B2(new_n803), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n820), .B2(new_n1137), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G150), .A2(new_n1023), .B1(new_n815), .B2(G125), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT120), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1015), .A2(G124), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1180), .B(new_n1200), .C1(new_n1066), .C2(new_n439), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n793), .B1(new_n1191), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n780), .B1(new_n251), .B2(new_n845), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n350), .A2(new_n913), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n376), .B(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1206), .B(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1203), .B(new_n1204), .C1(new_n1209), .C2(new_n791), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1206), .B(new_n1207), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n939), .B2(new_n944), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n961), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1209), .A2(G330), .A3(new_n938), .A4(new_n933), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1213), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1210), .B1(new_n1217), .B2(new_n777), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1120), .A2(new_n1129), .ZN(new_n1220));
  AND4_X1   g1020(.A1(KEYINPUT118), .A2(new_n1173), .A3(new_n1220), .A4(new_n1156), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT118), .B1(new_n1132), .B2(new_n1173), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1170), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1216), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1169), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1074), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1219), .B1(new_n1227), .B2(new_n1230), .ZN(G375));
  INV_X1    g1031(.A(new_n993), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1163), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1171), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n816), .A2(new_n861), .B1(new_n251), .B2(new_n813), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G137), .B2(new_n802), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n799), .A2(new_n342), .B1(new_n806), .B2(new_n1135), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n281), .B(new_n1237), .C1(new_n810), .C2(new_n1137), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1184), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G159), .B2(new_n835), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n835), .A2(G97), .B1(G303), .B2(new_n1015), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT122), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n281), .B1(new_n799), .B2(new_n206), .C1(new_n527), .C2(new_n809), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1048), .B1(G283), .B2(new_n802), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n603), .B2(new_n816), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(G77), .C2(new_n821), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1240), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1247), .A2(KEYINPUT123), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(KEYINPUT123), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n793), .A3(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n779), .C1(G68), .C2(new_n846), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1121), .B2(new_n790), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n777), .B(KEYINPUT121), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1167), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1234), .A2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G390), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n885), .ZN(new_n1258));
  OR4_X1    g1058(.A1(G396), .A2(G387), .A3(G393), .A4(new_n1258), .ZN(new_n1259));
  OR4_X1    g1059(.A1(G378), .A2(new_n1259), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g1060(.A1(new_n703), .A2(G213), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1178), .A2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G407), .B(G213), .C1(G375), .C2(new_n1263), .ZN(G409));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1233), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1233), .A2(new_n1265), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1074), .A3(new_n1171), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1255), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n885), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(G384), .A3(new_n1255), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1262), .A2(G2897), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(KEYINPUT125), .Z(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1270), .A2(new_n1271), .A3(new_n1274), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1219), .C1(new_n1227), .C2(new_n1230), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1210), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1253), .B1(new_n1228), .B2(new_n993), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n1226), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1279), .B1(G378), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1278), .B1(new_n1283), .B2(new_n1261), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G387), .A2(new_n1257), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G393), .B(G396), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G390), .B1(new_n1008), .B2(new_n1034), .ZN(new_n1287));
  OR3_X1    g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1286), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1284), .A2(KEYINPUT61), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT124), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1223), .A2(new_n1232), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1217), .B1(new_n1293), .B2(new_n1253), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1178), .B1(new_n1294), .B2(new_n1280), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1262), .B(new_n1272), .C1(new_n1295), .C2(new_n1279), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1296), .B2(KEYINPUT63), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(KEYINPUT63), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1272), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT57), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1176), .B1(new_n1301), .B2(new_n1223), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1228), .B2(new_n1217), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1178), .B(new_n1218), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1281), .A2(new_n1226), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G378), .B1(new_n1305), .B2(new_n1210), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1261), .B(new_n1299), .C1(new_n1304), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(KEYINPUT124), .A3(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1291), .A2(new_n1297), .A3(new_n1298), .A4(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1261), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1278), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1283), .A2(new_n1314), .A3(new_n1261), .A4(new_n1299), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1290), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1310), .A2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1178), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1299), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(G375), .A2(new_n1178), .A3(new_n1272), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1279), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1321), .B(new_n1322), .C1(KEYINPUT126), .C2(new_n1304), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1325), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1290), .A2(KEYINPUT127), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1331), .A2(new_n1327), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1329), .B1(new_n1330), .B2(new_n1332), .ZN(G402));
endmodule


