

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759;

  OR2_X1 U369 ( .A1(n643), .A2(G902), .ZN(n469) );
  XNOR2_X1 U370 ( .A(n469), .B(G472), .ZN(n616) );
  INV_X1 U371 ( .A(G953), .ZN(n751) );
  NOR2_X2 U372 ( .A1(n444), .A2(n348), .ZN(n443) );
  NOR2_X1 U373 ( .A1(n755), .A2(n759), .ZN(n579) );
  INV_X1 U374 ( .A(n629), .ZN(n660) );
  NOR2_X1 U375 ( .A1(n626), .A2(n390), .ZN(n384) );
  NOR2_X2 U376 ( .A1(n660), .A2(n659), .ZN(n665) );
  OR2_X1 U377 ( .A1(n730), .A2(G902), .ZN(n477) );
  INV_X1 U378 ( .A(KEYINPUT22), .ZN(n383) );
  NAND2_X1 U379 ( .A1(n450), .A2(n449), .ZN(n379) );
  NAND2_X1 U380 ( .A1(n452), .A2(n451), .ZN(n450) );
  NAND2_X1 U381 ( .A1(n395), .A2(n394), .ZN(n367) );
  XNOR2_X1 U382 ( .A(n568), .B(n569), .ZN(n755) );
  NAND2_X1 U383 ( .A1(n461), .A2(n458), .ZN(n457) );
  XNOR2_X1 U384 ( .A(n443), .B(n359), .ZN(n602) );
  NAND2_X1 U385 ( .A1(n456), .A2(KEYINPUT106), .ZN(n454) );
  XNOR2_X1 U386 ( .A(n384), .B(n383), .ZN(n632) );
  NAND2_X1 U387 ( .A1(n445), .A2(n474), .ZN(n444) );
  BUF_X1 U388 ( .A(n626), .Z(n430) );
  XNOR2_X1 U389 ( .A(n613), .B(n475), .ZN(n590) );
  INV_X1 U390 ( .A(n591), .ZN(n445) );
  OR2_X1 U391 ( .A1(n448), .A2(n447), .ZN(n653) );
  XNOR2_X1 U392 ( .A(n567), .B(n566), .ZN(n591) );
  XNOR2_X1 U393 ( .A(n501), .B(KEYINPUT38), .ZN(n448) );
  NOR2_X1 U394 ( .A1(n719), .A2(G902), .ZN(n560) );
  XNOR2_X1 U395 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U396 ( .A(G119), .B(KEYINPUT70), .ZN(n465) );
  XNOR2_X1 U397 ( .A(G116), .B(KEYINPUT3), .ZN(n496) );
  XNOR2_X1 U398 ( .A(n543), .B(n746), .ZN(n730) );
  OR2_X1 U399 ( .A1(n615), .A2(n427), .ZN(n405) );
  XNOR2_X2 U400 ( .A(n747), .B(G146), .ZN(n558) );
  XNOR2_X2 U401 ( .A(n369), .B(n525), .ZN(n747) );
  XNOR2_X2 U402 ( .A(n560), .B(n439), .ZN(n411) );
  XNOR2_X2 U403 ( .A(n477), .B(n476), .ZN(n629) );
  BUF_X1 U404 ( .A(n616), .Z(n427) );
  INV_X1 U405 ( .A(G134), .ZN(n467) );
  XNOR2_X1 U406 ( .A(n393), .B(KEYINPUT0), .ZN(n626) );
  XOR2_X1 U407 ( .A(G478), .B(n510), .Z(n575) );
  NAND2_X1 U408 ( .A1(n404), .A2(n403), .ZN(n402) );
  INV_X1 U409 ( .A(n654), .ZN(n403) );
  NAND2_X1 U410 ( .A1(n406), .A2(n405), .ZN(n404) );
  NAND2_X1 U411 ( .A1(n628), .A2(KEYINPUT105), .ZN(n462) );
  NAND2_X1 U412 ( .A1(n664), .A2(n460), .ZN(n459) );
  INV_X1 U413 ( .A(KEYINPUT105), .ZN(n460) );
  AND2_X1 U414 ( .A1(n420), .A2(n415), .ZN(n414) );
  XOR2_X1 U415 ( .A(KEYINPUT68), .B(G131), .Z(n524) );
  XNOR2_X1 U416 ( .A(n498), .B(n464), .ZN(n526) );
  XNOR2_X1 U417 ( .A(n465), .B(n497), .ZN(n464) );
  INV_X1 U418 ( .A(n590), .ZN(n474) );
  XNOR2_X1 U419 ( .A(n427), .B(KEYINPUT6), .ZN(n554) );
  NOR2_X1 U420 ( .A1(n430), .A2(KEYINPUT34), .ZN(n375) );
  INV_X1 U421 ( .A(n554), .ZN(n627) );
  XNOR2_X1 U422 ( .A(n500), .B(n485), .ZN(n582) );
  INV_X1 U423 ( .A(G469), .ZN(n439) );
  XNOR2_X1 U424 ( .A(n558), .B(n470), .ZN(n643) );
  XNOR2_X1 U425 ( .A(n532), .B(n471), .ZN(n470) );
  XNOR2_X1 U426 ( .A(n530), .B(n428), .ZN(n532) );
  INV_X1 U427 ( .A(n526), .ZN(n471) );
  XNOR2_X1 U428 ( .A(n492), .B(n349), .ZN(n733) );
  XNOR2_X1 U429 ( .A(G143), .B(G104), .ZN(n514) );
  XOR2_X1 U430 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n519) );
  XOR2_X1 U431 ( .A(KEYINPUT91), .B(KEYINPUT79), .Z(n490) );
  XNOR2_X1 U432 ( .A(n526), .B(n425), .ZN(n734) );
  XNOR2_X1 U433 ( .A(n499), .B(G122), .ZN(n425) );
  XOR2_X1 U434 ( .A(KEYINPUT16), .B(KEYINPUT73), .Z(n499) );
  XNOR2_X1 U435 ( .A(n733), .B(n493), .ZN(n557) );
  XNOR2_X1 U436 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n493) );
  XNOR2_X1 U437 ( .A(n546), .B(n544), .ZN(n476) );
  NOR2_X1 U438 ( .A1(n632), .A2(n627), .ZN(n631) );
  INV_X1 U439 ( .A(n575), .ZN(n595) );
  XNOR2_X1 U440 ( .A(n523), .B(n386), .ZN(n594) );
  XNOR2_X1 U441 ( .A(n522), .B(n392), .ZN(n386) );
  INV_X1 U442 ( .A(G475), .ZN(n392) );
  NOR2_X1 U443 ( .A1(n628), .A2(KEYINPUT87), .ZN(n397) );
  XNOR2_X1 U444 ( .A(n506), .B(n380), .ZN(n509) );
  XNOR2_X1 U445 ( .A(n558), .B(n407), .ZN(n719) );
  XNOR2_X1 U446 ( .A(n557), .B(n408), .ZN(n407) );
  XNOR2_X1 U447 ( .A(n559), .B(n409), .ZN(n408) );
  INV_X1 U448 ( .A(G140), .ZN(n409) );
  NOR2_X1 U449 ( .A1(G952), .A2(n751), .ZN(n732) );
  INV_X1 U450 ( .A(n449), .ZN(n378) );
  INV_X1 U451 ( .A(KEYINPUT69), .ZN(n497) );
  AND2_X1 U452 ( .A1(n448), .A2(n447), .ZN(n651) );
  INV_X1 U453 ( .A(n650), .ZN(n447) );
  AND2_X1 U454 ( .A1(n594), .A2(n391), .ZN(n389) );
  INV_X1 U455 ( .A(n659), .ZN(n391) );
  XOR2_X1 U456 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n529) );
  XNOR2_X1 U457 ( .A(n531), .B(n429), .ZN(n428) );
  INV_X1 U458 ( .A(KEYINPUT5), .ZN(n429) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n418) );
  INV_X1 U460 ( .A(KEYINPUT103), .ZN(n401) );
  NOR2_X1 U461 ( .A1(G953), .A2(G237), .ZN(n527) );
  XNOR2_X1 U462 ( .A(G902), .B(KEYINPUT15), .ZN(n486) );
  XOR2_X1 U463 ( .A(G137), .B(KEYINPUT4), .Z(n484) );
  XNOR2_X1 U464 ( .A(n472), .B(n601), .ZN(n381) );
  OR2_X1 U465 ( .A1(G237), .A2(G902), .ZN(n561) );
  INV_X1 U466 ( .A(n592), .ZN(n446) );
  AND2_X1 U467 ( .A1(n459), .A2(n354), .ZN(n458) );
  XNOR2_X1 U468 ( .A(G107), .B(KEYINPUT9), .ZN(n503) );
  XNOR2_X1 U469 ( .A(n435), .B(n434), .ZN(n648) );
  INV_X1 U470 ( .A(KEYINPUT81), .ZN(n434) );
  XNOR2_X1 U471 ( .A(n556), .B(KEYINPUT108), .ZN(n587) );
  AND2_X1 U472 ( .A1(n374), .A2(n372), .ZN(n371) );
  INV_X1 U473 ( .A(KEYINPUT109), .ZN(n475) );
  XNOR2_X1 U474 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U475 ( .A(n517), .B(n387), .ZN(n521) );
  XNOR2_X1 U476 ( .A(n520), .B(n516), .ZN(n387) );
  XNOR2_X1 U477 ( .A(n424), .B(n494), .ZN(n712) );
  XNOR2_X1 U478 ( .A(n495), .B(n734), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n491), .B(n350), .ZN(n495) );
  AND2_X1 U480 ( .A1(n682), .A2(n751), .ZN(n433) );
  XNOR2_X1 U481 ( .A(KEYINPUT32), .B(KEYINPUT67), .ZN(n432) );
  NAND2_X1 U482 ( .A1(n631), .A2(n630), .ZN(n400) );
  NOR2_X1 U483 ( .A1(n595), .A2(n580), .ZN(n703) );
  NOR2_X1 U484 ( .A1(n575), .A2(n594), .ZN(n700) );
  INV_X1 U485 ( .A(n405), .ZN(n690) );
  AND2_X1 U486 ( .A1(n398), .A2(n396), .ZN(n395) );
  NOR2_X1 U487 ( .A1(n397), .A2(n660), .ZN(n396) );
  INV_X1 U488 ( .A(n732), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n726), .B(n423), .ZN(n728) );
  XNOR2_X1 U490 ( .A(n727), .B(KEYINPUT124), .ZN(n423) );
  XNOR2_X1 U491 ( .A(n717), .B(n431), .ZN(n720) );
  XNOR2_X1 U492 ( .A(n719), .B(n718), .ZN(n431) );
  XOR2_X1 U493 ( .A(n351), .B(n536), .Z(n347) );
  OR2_X1 U494 ( .A1(n448), .A2(n446), .ZN(n348) );
  XOR2_X1 U495 ( .A(G104), .B(G107), .Z(n349) );
  XOR2_X1 U496 ( .A(n490), .B(n489), .Z(n350) );
  XOR2_X1 U497 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n351) );
  AND2_X1 U498 ( .A1(n482), .A2(n481), .ZN(n352) );
  AND2_X1 U499 ( .A1(n450), .A2(n377), .ZN(n353) );
  AND2_X1 U500 ( .A1(n633), .A2(n660), .ZN(n354) );
  XOR2_X1 U501 ( .A(G116), .B(G122), .Z(n355) );
  AND2_X1 U502 ( .A1(n628), .A2(KEYINPUT87), .ZN(n356) );
  AND2_X1 U503 ( .A1(n648), .A2(n647), .ZN(n357) );
  AND2_X1 U504 ( .A1(n479), .A2(n757), .ZN(n358) );
  XNOR2_X1 U505 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n359) );
  NOR2_X1 U506 ( .A1(n680), .A2(n410), .ZN(n360) );
  XOR2_X1 U507 ( .A(n643), .B(KEYINPUT62), .Z(n361) );
  XNOR2_X1 U508 ( .A(n486), .B(KEYINPUT90), .ZN(n533) );
  INV_X1 U509 ( .A(KEYINPUT106), .ZN(n463) );
  XOR2_X1 U510 ( .A(n684), .B(KEYINPUT123), .Z(n362) );
  AND2_X2 U511 ( .A1(n440), .A2(n441), .ZN(n363) );
  AND2_X2 U512 ( .A1(n440), .A2(n441), .ZN(n478) );
  NAND2_X1 U513 ( .A1(n642), .A2(n641), .ZN(n440) );
  INV_X1 U514 ( .A(n456), .ZN(n455) );
  NAND2_X1 U515 ( .A1(n455), .A2(n463), .ZN(n449) );
  NOR2_X1 U516 ( .A1(n466), .A2(n533), .ZN(n421) );
  NAND2_X1 U517 ( .A1(n381), .A2(n358), .ZN(n466) );
  XNOR2_X1 U518 ( .A(n347), .B(n539), .ZN(n542) );
  BUF_X1 U519 ( .A(n586), .Z(n364) );
  NAND2_X1 U520 ( .A1(n582), .A2(n650), .ZN(n586) );
  XNOR2_X1 U521 ( .A(n364), .B(n583), .ZN(n365) );
  XNOR2_X1 U522 ( .A(n586), .B(n583), .ZN(n609) );
  XNOR2_X1 U523 ( .A(n366), .B(n362), .ZN(G75) );
  NAND2_X1 U524 ( .A1(n683), .A2(n433), .ZN(n366) );
  NAND2_X1 U525 ( .A1(n638), .A2(n367), .ZN(n419) );
  XNOR2_X1 U526 ( .A(n367), .B(n685), .ZN(G3) );
  NAND2_X1 U527 ( .A1(n421), .A2(n368), .ZN(n639) );
  OR2_X1 U528 ( .A1(n368), .A2(KEYINPUT2), .ZN(n435) );
  NAND2_X1 U529 ( .A1(n368), .A2(n751), .ZN(n738) );
  NAND2_X1 U530 ( .A1(n422), .A2(n368), .ZN(n436) );
  XNOR2_X2 U531 ( .A(n382), .B(KEYINPUT45), .ZN(n368) );
  XNOR2_X1 U532 ( .A(n369), .B(n355), .ZN(n380) );
  XNOR2_X2 U533 ( .A(n502), .B(n467), .ZN(n369) );
  NAND2_X1 U534 ( .A1(n371), .A2(n370), .ZN(n624) );
  NAND2_X1 U535 ( .A1(n410), .A2(KEYINPUT34), .ZN(n370) );
  AND2_X1 U536 ( .A1(n373), .A2(n621), .ZN(n372) );
  NAND2_X1 U537 ( .A1(n430), .A2(KEYINPUT34), .ZN(n373) );
  NAND2_X1 U538 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U539 ( .A(n410), .ZN(n376) );
  XNOR2_X2 U540 ( .A(n620), .B(n619), .ZN(n410) );
  NOR2_X1 U541 ( .A1(n378), .A2(n637), .ZN(n377) );
  NOR2_X1 U542 ( .A1(n379), .A2(n758), .ZN(n636) );
  NAND2_X1 U543 ( .A1(n379), .A2(n483), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n379), .B(n412), .ZN(G12) );
  NAND2_X1 U545 ( .A1(n602), .A2(n700), .ZN(n568) );
  NAND2_X1 U546 ( .A1(n625), .A2(n418), .ZN(n417) );
  NOR2_X1 U547 ( .A1(n419), .A2(n417), .ZN(n416) );
  NAND2_X1 U548 ( .A1(n416), .A2(n385), .ZN(n382) );
  NOR2_X1 U549 ( .A1(n587), .A2(n562), .ZN(n563) );
  INV_X1 U550 ( .A(n708), .ZN(n479) );
  NAND2_X1 U551 ( .A1(n414), .A2(n352), .ZN(n385) );
  NAND2_X1 U552 ( .A1(n388), .A2(n650), .ZN(n567) );
  XNOR2_X1 U553 ( .A(n616), .B(KEYINPUT104), .ZN(n388) );
  NAND2_X1 U554 ( .A1(n595), .A2(n594), .ZN(n652) );
  NAND2_X1 U555 ( .A1(n389), .A2(n595), .ZN(n390) );
  NAND2_X1 U556 ( .A1(n609), .A2(n610), .ZN(n393) );
  OR2_X1 U557 ( .A1(n399), .A2(KEYINPUT87), .ZN(n394) );
  NAND2_X1 U558 ( .A1(n399), .A2(n356), .ZN(n398) );
  XNOR2_X1 U559 ( .A(n631), .B(KEYINPUT86), .ZN(n399) );
  NAND2_X1 U560 ( .A1(n758), .A2(n483), .ZN(n415) );
  XNOR2_X2 U561 ( .A(n400), .B(n432), .ZN(n758) );
  INV_X1 U562 ( .A(n704), .ZN(n406) );
  NOR2_X1 U563 ( .A1(n658), .A2(n410), .ZN(n674) );
  NAND2_X1 U564 ( .A1(n665), .A2(n411), .ZN(n613) );
  XNOR2_X1 U565 ( .A(n411), .B(KEYINPUT1), .ZN(n604) );
  NAND2_X1 U566 ( .A1(n574), .A2(n411), .ZN(n581) );
  INV_X1 U567 ( .A(G110), .ZN(n412) );
  AND2_X1 U568 ( .A1(n357), .A2(n441), .ZN(n649) );
  XNOR2_X2 U569 ( .A(n436), .B(n413), .ZN(n441) );
  INV_X1 U570 ( .A(KEYINPUT75), .ZN(n413) );
  NAND2_X1 U571 ( .A1(n353), .A2(n480), .ZN(n420) );
  NOR2_X1 U572 ( .A1(n466), .A2(n646), .ZN(n422) );
  NOR2_X2 U573 ( .A1(n725), .A2(n732), .ZN(n442) );
  NOR2_X2 U574 ( .A1(n715), .A2(n732), .ZN(n716) );
  NAND2_X1 U575 ( .A1(n635), .A2(KEYINPUT66), .ZN(n481) );
  NAND2_X1 U576 ( .A1(n478), .A2(G210), .ZN(n713) );
  XNOR2_X1 U577 ( .A(n713), .B(n714), .ZN(n715) );
  INV_X1 U578 ( .A(n426), .ZN(n461) );
  NOR2_X1 U579 ( .A1(n632), .A2(n462), .ZN(n426) );
  XNOR2_X1 U580 ( .A(n644), .B(n361), .ZN(n438) );
  XNOR2_X1 U581 ( .A(n488), .B(n502), .ZN(n491) );
  XNOR2_X1 U582 ( .A(n557), .B(KEYINPUT4), .ZN(n494) );
  NAND2_X1 U583 ( .A1(n438), .A2(n437), .ZN(n645) );
  XNOR2_X1 U584 ( .A(n442), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U585 ( .A1(n457), .A2(KEYINPUT106), .ZN(n451) );
  NAND2_X1 U586 ( .A1(n453), .A2(n454), .ZN(n452) );
  INV_X1 U587 ( .A(n457), .ZN(n453) );
  NAND2_X1 U588 ( .A1(n632), .A2(n460), .ZN(n456) );
  NAND2_X1 U589 ( .A1(n466), .A2(n646), .ZN(n647) );
  XNOR2_X1 U590 ( .A(n466), .B(n750), .ZN(n752) );
  XNOR2_X2 U591 ( .A(n468), .B(G128), .ZN(n502) );
  XNOR2_X2 U592 ( .A(G143), .B(KEYINPUT65), .ZN(n468) );
  NAND2_X1 U593 ( .A1(n473), .A2(n600), .ZN(n472) );
  XNOR2_X1 U594 ( .A(n579), .B(n578), .ZN(n473) );
  NAND2_X1 U595 ( .A1(n478), .A2(G475), .ZN(n724) );
  NAND2_X1 U596 ( .A1(n363), .A2(G472), .ZN(n644) );
  NAND2_X1 U597 ( .A1(n363), .A2(G469), .ZN(n717) );
  NAND2_X1 U598 ( .A1(n363), .A2(G478), .ZN(n726) );
  NAND2_X1 U599 ( .A1(n363), .A2(G217), .ZN(n729) );
  INV_X1 U600 ( .A(n758), .ZN(n480) );
  NOR2_X1 U601 ( .A1(n635), .A2(KEYINPUT66), .ZN(n483) );
  AND2_X1 U602 ( .A1(G210), .A2(n561), .ZN(n485) );
  INV_X1 U603 ( .A(KEYINPUT66), .ZN(n637) );
  XNOR2_X1 U604 ( .A(n511), .B(n487), .ZN(n488) );
  XNOR2_X1 U605 ( .A(n565), .B(KEYINPUT110), .ZN(n566) );
  XNOR2_X1 U606 ( .A(n524), .B(n484), .ZN(n525) );
  INV_X1 U607 ( .A(n533), .ZN(n640) );
  XOR2_X2 U608 ( .A(G146), .B(G125), .Z(n511) );
  XOR2_X1 U609 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n487) );
  NAND2_X1 U610 ( .A1(G224), .A2(n751), .ZN(n489) );
  XNOR2_X1 U611 ( .A(G101), .B(G110), .ZN(n492) );
  XNOR2_X1 U612 ( .A(n496), .B(G113), .ZN(n498) );
  NAND2_X1 U613 ( .A1(n712), .A2(n533), .ZN(n500) );
  BUF_X1 U614 ( .A(n582), .Z(n501) );
  XOR2_X1 U615 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n504) );
  XNOR2_X1 U616 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U617 ( .A(n505), .B(KEYINPUT7), .Z(n506) );
  NAND2_X1 U618 ( .A1(G234), .A2(n751), .ZN(n507) );
  XOR2_X1 U619 ( .A(KEYINPUT8), .B(n507), .Z(n540) );
  NAND2_X1 U620 ( .A1(G217), .A2(n540), .ZN(n508) );
  XNOR2_X1 U621 ( .A(n509), .B(n508), .ZN(n727) );
  NOR2_X1 U622 ( .A1(G902), .A2(n727), .ZN(n510) );
  XNOR2_X1 U623 ( .A(n511), .B(G140), .ZN(n512) );
  XNOR2_X1 U624 ( .A(n512), .B(KEYINPUT10), .ZN(n746) );
  XNOR2_X1 U625 ( .A(G113), .B(n524), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n513), .B(G122), .ZN(n517) );
  XOR2_X1 U627 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n515) );
  XNOR2_X1 U628 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U629 ( .A1(G214), .A2(n527), .ZN(n518) );
  XNOR2_X1 U630 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U631 ( .A(n746), .B(n521), .ZN(n722) );
  NOR2_X1 U632 ( .A1(G902), .A2(n722), .ZN(n523) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n522) );
  NAND2_X1 U634 ( .A1(n527), .A2(G210), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U636 ( .A(G101), .B(KEYINPUT74), .ZN(n531) );
  NAND2_X1 U637 ( .A1(G234), .A2(n533), .ZN(n534) );
  XNOR2_X1 U638 ( .A(n534), .B(KEYINPUT20), .ZN(n545) );
  NAND2_X1 U639 ( .A1(n545), .A2(G221), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n535), .B(KEYINPUT21), .ZN(n659) );
  XNOR2_X1 U641 ( .A(KEYINPUT78), .B(KEYINPUT24), .ZN(n536) );
  XOR2_X1 U642 ( .A(G110), .B(G128), .Z(n538) );
  XNOR2_X1 U643 ( .A(G119), .B(G137), .ZN(n537) );
  XNOR2_X1 U644 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U645 ( .A1(G221), .A2(n540), .ZN(n541) );
  XNOR2_X1 U646 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n544) );
  NAND2_X1 U647 ( .A1(n545), .A2(G217), .ZN(n546) );
  NOR2_X1 U648 ( .A1(n659), .A2(n629), .ZN(n553) );
  NAND2_X1 U649 ( .A1(G234), .A2(G237), .ZN(n547) );
  XNOR2_X1 U650 ( .A(n547), .B(KEYINPUT14), .ZN(n550) );
  NAND2_X1 U651 ( .A1(G952), .A2(n550), .ZN(n548) );
  XNOR2_X1 U652 ( .A(KEYINPUT92), .B(n548), .ZN(n678) );
  NOR2_X1 U653 ( .A1(n678), .A2(G953), .ZN(n549) );
  XNOR2_X1 U654 ( .A(n549), .B(KEYINPUT93), .ZN(n607) );
  NAND2_X1 U655 ( .A1(G902), .A2(n550), .ZN(n605) );
  NOR2_X1 U656 ( .A1(G900), .A2(n605), .ZN(n551) );
  NAND2_X1 U657 ( .A1(G953), .A2(n551), .ZN(n552) );
  NAND2_X1 U658 ( .A1(n607), .A2(n552), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n553), .A2(n592), .ZN(n570) );
  NOR2_X1 U660 ( .A1(n554), .A2(n570), .ZN(n555) );
  NAND2_X1 U661 ( .A1(n700), .A2(n555), .ZN(n556) );
  NAND2_X1 U662 ( .A1(n751), .A2(G227), .ZN(n559) );
  INV_X1 U663 ( .A(n604), .ZN(n628) );
  NAND2_X1 U664 ( .A1(G214), .A2(n561), .ZN(n650) );
  NAND2_X1 U665 ( .A1(n628), .A2(n650), .ZN(n562) );
  XNOR2_X1 U666 ( .A(n563), .B(KEYINPUT43), .ZN(n564) );
  NOR2_X1 U667 ( .A1(n501), .A2(n564), .ZN(n708) );
  XOR2_X1 U668 ( .A(KEYINPUT114), .B(KEYINPUT40), .Z(n569) );
  XOR2_X1 U669 ( .A(KEYINPUT111), .B(KEYINPUT30), .Z(n565) );
  XOR2_X1 U670 ( .A(KEYINPUT104), .B(n427), .Z(n633) );
  NOR2_X1 U671 ( .A1(n633), .A2(n570), .ZN(n573) );
  XOR2_X1 U672 ( .A(KEYINPUT28), .B(KEYINPUT113), .Z(n571) );
  XNOR2_X1 U673 ( .A(KEYINPUT112), .B(n571), .ZN(n572) );
  XNOR2_X1 U674 ( .A(n573), .B(n572), .ZN(n574) );
  NOR2_X1 U675 ( .A1(n652), .A2(n653), .ZN(n576) );
  XNOR2_X1 U676 ( .A(n576), .B(KEYINPUT41), .ZN(n680) );
  NOR2_X1 U677 ( .A1(n581), .A2(n680), .ZN(n577) );
  XNOR2_X1 U678 ( .A(n577), .B(KEYINPUT42), .ZN(n759) );
  XNOR2_X1 U679 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n578) );
  INV_X1 U680 ( .A(n594), .ZN(n580) );
  NOR2_X1 U681 ( .A1(n703), .A2(n700), .ZN(n654) );
  INV_X1 U682 ( .A(n581), .ZN(n584) );
  XNOR2_X1 U683 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n583) );
  NAND2_X1 U684 ( .A1(n584), .A2(n365), .ZN(n697) );
  NOR2_X1 U685 ( .A1(n654), .A2(n697), .ZN(n585) );
  XOR2_X1 U686 ( .A(n585), .B(KEYINPUT47), .Z(n599) );
  NOR2_X1 U687 ( .A1(n587), .A2(n364), .ZN(n588) );
  XNOR2_X1 U688 ( .A(n588), .B(KEYINPUT36), .ZN(n589) );
  INV_X1 U689 ( .A(n628), .ZN(n664) );
  NAND2_X1 U690 ( .A1(n589), .A2(n664), .ZN(n707) );
  NOR2_X1 U691 ( .A1(n591), .A2(n590), .ZN(n593) );
  AND2_X1 U692 ( .A1(n593), .A2(n592), .ZN(n596) );
  NOR2_X1 U693 ( .A1(n595), .A2(n594), .ZN(n621) );
  AND2_X1 U694 ( .A1(n596), .A2(n621), .ZN(n597) );
  NAND2_X1 U695 ( .A1(n501), .A2(n597), .ZN(n696) );
  NAND2_X1 U696 ( .A1(n707), .A2(n696), .ZN(n598) );
  NOR2_X1 U697 ( .A1(n599), .A2(n598), .ZN(n600) );
  INV_X1 U698 ( .A(KEYINPUT48), .ZN(n601) );
  NAND2_X1 U699 ( .A1(n602), .A2(n703), .ZN(n603) );
  XOR2_X1 U700 ( .A(KEYINPUT115), .B(n603), .Z(n757) );
  NAND2_X1 U701 ( .A1(n665), .A2(n604), .ZN(n617) );
  INV_X1 U702 ( .A(n427), .ZN(n663) );
  NOR2_X1 U703 ( .A1(n617), .A2(n663), .ZN(n670) );
  INV_X1 U704 ( .A(n605), .ZN(n606) );
  NOR2_X1 U705 ( .A1(G898), .A2(n751), .ZN(n736) );
  NAND2_X1 U706 ( .A1(n606), .A2(n736), .ZN(n608) );
  NAND2_X1 U707 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U708 ( .A(n430), .ZN(n611) );
  NAND2_X1 U709 ( .A1(n670), .A2(n611), .ZN(n612) );
  XNOR2_X1 U710 ( .A(KEYINPUT31), .B(n612), .ZN(n704) );
  NOR2_X1 U711 ( .A1(n430), .A2(n613), .ZN(n614) );
  XNOR2_X1 U712 ( .A(n614), .B(KEYINPUT95), .ZN(n615) );
  XNOR2_X1 U713 ( .A(n617), .B(KEYINPUT107), .ZN(n618) );
  NAND2_X1 U714 ( .A1(n627), .A2(n618), .ZN(n620) );
  INV_X1 U715 ( .A(KEYINPUT33), .ZN(n619) );
  XNOR2_X1 U716 ( .A(KEYINPUT35), .B(KEYINPUT80), .ZN(n622) );
  XNOR2_X1 U717 ( .A(n622), .B(KEYINPUT84), .ZN(n623) );
  XNOR2_X2 U718 ( .A(n624), .B(n623), .ZN(n756) );
  NAND2_X1 U719 ( .A1(KEYINPUT44), .A2(n756), .ZN(n625) );
  NOR2_X1 U720 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U721 ( .A1(n756), .A2(KEYINPUT44), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n636), .A2(n634), .ZN(n638) );
  INV_X1 U723 ( .A(KEYINPUT44), .ZN(n635) );
  XNOR2_X1 U724 ( .A(n639), .B(KEYINPUT82), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  XNOR2_X1 U726 ( .A(n645), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U727 ( .A(KEYINPUT2), .ZN(n646) );
  XNOR2_X1 U728 ( .A(n649), .B(KEYINPUT83), .ZN(n683) );
  XNOR2_X1 U729 ( .A(KEYINPUT121), .B(KEYINPUT52), .ZN(n676) );
  NOR2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n656) );
  NOR2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT120), .ZN(n658) );
  AND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n661), .B(KEYINPUT49), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT50), .ZN(n667) );
  NOR2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U740 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT51), .B(n671), .Z(n672) );
  NOR2_X1 U742 ( .A1(n680), .A2(n672), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U744 ( .A(n676), .B(n675), .Z(n677) );
  NOR2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n679), .B(KEYINPUT122), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n681), .A2(n360), .ZN(n682) );
  INV_X1 U748 ( .A(KEYINPUT53), .ZN(n684) );
  XNOR2_X1 U749 ( .A(G101), .B(KEYINPUT116), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n690), .A2(n700), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(G104), .ZN(G6) );
  XOR2_X1 U752 ( .A(KEYINPUT27), .B(KEYINPUT118), .Z(n688) );
  XNOR2_X1 U753 ( .A(G107), .B(KEYINPUT117), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U755 ( .A(KEYINPUT26), .B(n689), .Z(n692) );
  NAND2_X1 U756 ( .A1(n690), .A2(n703), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n692), .B(n691), .ZN(G9) );
  INV_X1 U758 ( .A(n703), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n693), .A2(n697), .ZN(n695) );
  XNOR2_X1 U760 ( .A(G128), .B(KEYINPUT29), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n695), .B(n694), .ZN(G30) );
  XNOR2_X1 U762 ( .A(G143), .B(n696), .ZN(G45) );
  INV_X1 U763 ( .A(n700), .ZN(n698) );
  NOR2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U765 ( .A(G146), .B(n699), .Z(G48) );
  XOR2_X1 U766 ( .A(G113), .B(KEYINPUT119), .Z(n702) );
  NAND2_X1 U767 ( .A1(n704), .A2(n700), .ZN(n701) );
  XNOR2_X1 U768 ( .A(n702), .B(n701), .ZN(G15) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U770 ( .A(n705), .B(G116), .ZN(G18) );
  XOR2_X1 U771 ( .A(G125), .B(KEYINPUT37), .Z(n706) );
  XNOR2_X1 U772 ( .A(n707), .B(n706), .ZN(G27) );
  XOR2_X1 U773 ( .A(G140), .B(n708), .Z(G42) );
  XOR2_X1 U774 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n710) );
  XNOR2_X1 U775 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n712), .B(n711), .ZN(n714) );
  XNOR2_X1 U778 ( .A(n716), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n718) );
  NOR2_X1 U780 ( .A1(n732), .A2(n720), .ZN(G54) );
  INV_X1 U781 ( .A(KEYINPUT59), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U783 ( .A1(n732), .A2(n728), .ZN(G63) );
  XNOR2_X1 U784 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U785 ( .A1(n732), .A2(n731), .ZN(G66) );
  XNOR2_X1 U786 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n735), .B(KEYINPUT127), .ZN(n737) );
  NOR2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n738), .B(KEYINPUT126), .ZN(n743) );
  XOR2_X1 U790 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n740) );
  NAND2_X1 U791 ( .A1(G224), .A2(G953), .ZN(n739) );
  XNOR2_X1 U792 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U793 ( .A1(n741), .A2(G898), .ZN(n742) );
  NAND2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n745), .B(n744), .ZN(G69) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(n750) );
  XNOR2_X1 U797 ( .A(G227), .B(n750), .ZN(n748) );
  NAND2_X1 U798 ( .A1(G900), .A2(n748), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n749), .A2(G953), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U802 ( .A(n755), .B(G131), .Z(G33) );
  XOR2_X1 U803 ( .A(n756), .B(G122), .Z(G24) );
  XNOR2_X1 U804 ( .A(G134), .B(n757), .ZN(G36) );
  XOR2_X1 U805 ( .A(n758), .B(G119), .Z(G21) );
  XOR2_X1 U806 ( .A(G137), .B(n759), .Z(G39) );
endmodule

