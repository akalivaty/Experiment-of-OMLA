

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  XNOR2_X1 U325 ( .A(KEYINPUT110), .B(KEYINPUT45), .ZN(n372) );
  XNOR2_X1 U326 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U327 ( .A(G36GAT), .B(G190GAT), .Z(n391) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n381) );
  XNOR2_X1 U329 ( .A(n382), .B(n381), .ZN(n546) );
  XOR2_X1 U330 ( .A(n311), .B(n349), .Z(n458) );
  XNOR2_X1 U331 ( .A(n455), .B(KEYINPUT58), .ZN(n456) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(n391), .B(KEYINPUT11), .Z(n294) );
  NAND2_X1 U334 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U335 ( .A(n294), .B(n293), .Z(n302) );
  XOR2_X1 U336 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n296) );
  XNOR2_X1 U337 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n298) );
  INV_X1 U339 ( .A(KEYINPUT79), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n300) );
  XOR2_X1 U341 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XNOR2_X1 U342 ( .A(G218GAT), .B(n422), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT80), .Z(n413) );
  XOR2_X1 U346 ( .A(KEYINPUT73), .B(G92GAT), .Z(n304) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(KEYINPUT74), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U349 ( .A(G85GAT), .B(n305), .ZN(n367) );
  XOR2_X1 U350 ( .A(n413), .B(n367), .Z(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U352 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n309) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G29GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT7), .B(n310), .Z(n349) );
  XOR2_X1 U356 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XOR2_X1 U357 ( .A(n442), .B(KEYINPUT84), .Z(n313) );
  NAND2_X1 U358 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U360 ( .A(KEYINPUT15), .B(KEYINPUT83), .Z(n315) );
  XNOR2_X1 U361 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U363 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U364 ( .A(G1GAT), .B(KEYINPUT70), .Z(n335) );
  XOR2_X1 U365 ( .A(KEYINPUT82), .B(G64GAT), .Z(n319) );
  XNOR2_X1 U366 ( .A(G211GAT), .B(G155GAT), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U368 ( .A(n335), .B(n320), .Z(n322) );
  NAND2_X1 U369 ( .A1(n321), .A2(n322), .ZN(n326) );
  INV_X1 U370 ( .A(n321), .ZN(n324) );
  INV_X1 U371 ( .A(n322), .ZN(n323) );
  NAND2_X1 U372 ( .A1(n324), .A2(n323), .ZN(n325) );
  NAND2_X1 U373 ( .A1(n326), .A2(n325), .ZN(n330) );
  XOR2_X1 U374 ( .A(G8GAT), .B(KEYINPUT81), .Z(n383) );
  XOR2_X1 U375 ( .A(G57GAT), .B(KEYINPUT13), .Z(n354) );
  XOR2_X1 U376 ( .A(n383), .B(n354), .Z(n328) );
  XNOR2_X1 U377 ( .A(G183GAT), .B(G71GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n332) );
  XNOR2_X1 U380 ( .A(G22GAT), .B(G78GAT), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n556) );
  INV_X1 U382 ( .A(n556), .ZN(n588) );
  NAND2_X1 U383 ( .A1(n458), .A2(n588), .ZN(n370) );
  XOR2_X1 U384 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n334) );
  XNOR2_X1 U385 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U387 ( .A(G50GAT), .B(G36GAT), .Z(n337) );
  XOR2_X1 U388 ( .A(G141GAT), .B(G22GAT), .Z(n428) );
  XNOR2_X1 U389 ( .A(n428), .B(n335), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n341) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U394 ( .A(G197GAT), .B(G113GAT), .Z(n343) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G15GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U397 ( .A(n345), .B(n344), .Z(n351) );
  XOR2_X1 U398 ( .A(G8GAT), .B(KEYINPUT68), .Z(n347) );
  XNOR2_X1 U399 ( .A(KEYINPUT67), .B(KEYINPUT71), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U402 ( .A(n351), .B(n350), .Z(n549) );
  INV_X1 U403 ( .A(n549), .ZN(n578) );
  XOR2_X1 U404 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n353) );
  XNOR2_X1 U405 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n352) );
  XOR2_X1 U406 ( .A(n353), .B(n352), .Z(n365) );
  XOR2_X1 U407 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n356) );
  XOR2_X1 U408 ( .A(G176GAT), .B(G64GAT), .Z(n386) );
  XNOR2_X1 U409 ( .A(n354), .B(n386), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U411 ( .A(n357), .B(KEYINPUT76), .Z(n363) );
  XNOR2_X1 U412 ( .A(G106GAT), .B(G78GAT), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n358), .B(G148GAT), .ZN(n424) );
  XOR2_X1 U414 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  XOR2_X1 U415 ( .A(n424), .B(n445), .Z(n360) );
  NAND2_X1 U416 ( .A1(G230GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U418 ( .A(G204GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U421 ( .A(n367), .B(n366), .Z(n584) );
  XOR2_X1 U422 ( .A(KEYINPUT41), .B(n584), .Z(n565) );
  NOR2_X1 U423 ( .A1(n578), .A2(n565), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n368), .B(KEYINPUT46), .ZN(n369) );
  NOR2_X1 U425 ( .A1(n370), .A2(n369), .ZN(n371) );
  XOR2_X1 U426 ( .A(KEYINPUT47), .B(n371), .Z(n380) );
  XNOR2_X1 U427 ( .A(n458), .B(KEYINPUT36), .ZN(n591) );
  NOR2_X1 U428 ( .A1(n588), .A2(n591), .ZN(n373) );
  AND2_X1 U429 ( .A1(n374), .A2(n584), .ZN(n376) );
  INV_X1 U430 ( .A(KEYINPUT111), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  AND2_X1 U432 ( .A1(n377), .A2(n578), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n378), .B(KEYINPUT112), .ZN(n379) );
  NOR2_X1 U434 ( .A1(n380), .A2(n379), .ZN(n382) );
  XOR2_X1 U435 ( .A(n383), .B(G92GAT), .Z(n385) );
  NAND2_X1 U436 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U438 ( .A(n387), .B(n386), .Z(n393) );
  XOR2_X1 U439 ( .A(G211GAT), .B(G218GAT), .Z(n389) );
  XNOR2_X1 U440 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(n390), .ZN(n433) );
  XOR2_X1 U443 ( .A(n433), .B(n391), .Z(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U445 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n395) );
  XNOR2_X1 U446 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U448 ( .A(G169GAT), .B(n396), .ZN(n440) );
  INV_X1 U449 ( .A(n440), .ZN(n397) );
  XOR2_X1 U450 ( .A(n398), .B(n397), .Z(n465) );
  NOR2_X1 U451 ( .A1(n546), .A2(n465), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n399), .B(KEYINPUT54), .ZN(n574) );
  XOR2_X1 U453 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n401) );
  XNOR2_X1 U454 ( .A(G1GAT), .B(G57GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n419) );
  XOR2_X1 U456 ( .A(G85GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT4), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U460 ( .A(G141GAT), .B(G127GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U462 ( .A(n407), .B(n406), .Z(n412) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n409) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U466 ( .A(KEYINPUT90), .B(n410), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U468 ( .A(n414), .B(n413), .Z(n417) );
  XOR2_X1 U469 ( .A(G113GAT), .B(KEYINPUT0), .Z(n441) );
  XNOR2_X1 U470 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n415), .B(KEYINPUT2), .ZN(n423) );
  XNOR2_X1 U472 ( .A(n441), .B(n423), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n575) );
  XOR2_X1 U475 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n421) );
  XNOR2_X1 U476 ( .A(KEYINPUT89), .B(KEYINPUT24), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n432) );
  XOR2_X1 U478 ( .A(n423), .B(n422), .Z(n430) );
  XOR2_X1 U479 ( .A(n424), .B(KEYINPUT22), .Z(n426) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n473) );
  AND2_X1 U486 ( .A1(n575), .A2(n473), .ZN(n435) );
  NAND2_X1 U487 ( .A1(n574), .A2(n435), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n436), .B(KEYINPUT55), .ZN(n454) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n438) );
  XNOR2_X1 U490 ( .A(G43GAT), .B(G99GAT), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U492 ( .A(n440), .B(n439), .Z(n453) );
  XOR2_X1 U493 ( .A(G134GAT), .B(G190GAT), .Z(n444) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U496 ( .A(n446), .B(n445), .Z(n451) );
  XOR2_X1 U497 ( .A(G176GAT), .B(KEYINPUT85), .Z(n448) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(KEYINPUT20), .B(n449), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U502 ( .A(n453), .B(n452), .Z(n474) );
  INV_X1 U503 ( .A(n474), .ZN(n531) );
  NAND2_X1 U504 ( .A1(n454), .A2(n531), .ZN(n570) );
  NOR2_X1 U505 ( .A1(n458), .A2(n570), .ZN(n457) );
  INV_X1 U506 ( .A(G190GAT), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n479) );
  NAND2_X1 U508 ( .A1(n549), .A2(n584), .ZN(n495) );
  INV_X1 U509 ( .A(n458), .ZN(n559) );
  NOR2_X1 U510 ( .A1(n588), .A2(n559), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT16), .ZN(n477) );
  NOR2_X1 U512 ( .A1(n465), .A2(n474), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT93), .ZN(n461) );
  NAND2_X1 U514 ( .A1(n461), .A2(n473), .ZN(n463) );
  XOR2_X1 U515 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n462) );
  XOR2_X1 U516 ( .A(n463), .B(n462), .Z(n469) );
  NOR2_X1 U517 ( .A1(n531), .A2(n473), .ZN(n464) );
  XNOR2_X1 U518 ( .A(KEYINPUT26), .B(n464), .ZN(n576) );
  INV_X1 U519 ( .A(n576), .ZN(n466) );
  INV_X1 U520 ( .A(n465), .ZN(n523) );
  XOR2_X1 U521 ( .A(n523), .B(KEYINPUT27), .Z(n472) );
  NOR2_X1 U522 ( .A1(n466), .A2(n472), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT92), .B(n467), .ZN(n468) );
  NOR2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U525 ( .A(KEYINPUT95), .B(n470), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n471), .A2(n575), .ZN(n476) );
  OR2_X1 U527 ( .A1(n575), .A2(n472), .ZN(n545) );
  XOR2_X1 U528 ( .A(KEYINPUT28), .B(n473), .Z(n527) );
  NOR2_X1 U529 ( .A1(n545), .A2(n527), .ZN(n530) );
  NAND2_X1 U530 ( .A1(n530), .A2(n474), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n476), .A2(n475), .ZN(n491) );
  NAND2_X1 U532 ( .A1(n477), .A2(n491), .ZN(n508) );
  NOR2_X1 U533 ( .A1(n495), .A2(n508), .ZN(n487) );
  INV_X1 U534 ( .A(n575), .ZN(n521) );
  NAND2_X1 U535 ( .A1(n487), .A2(n521), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n482) );
  NAND2_X1 U539 ( .A1(n487), .A2(n523), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n485) );
  NAND2_X1 U543 ( .A1(n487), .A2(n531), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U545 ( .A(G15GAT), .B(n486), .Z(G1326GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n489) );
  NAND2_X1 U547 ( .A1(n487), .A2(n527), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(n490), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U551 ( .A1(n588), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT102), .B(n492), .ZN(n493) );
  NOR2_X1 U553 ( .A1(n493), .A2(n591), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT37), .ZN(n519) );
  NOR2_X1 U555 ( .A1(n519), .A2(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT38), .B(n496), .ZN(n504) );
  NAND2_X1 U557 ( .A1(n521), .A2(n504), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT103), .Z(n500) );
  NAND2_X1 U560 ( .A1(n504), .A2(n523), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n502) );
  NAND2_X1 U563 ( .A1(n531), .A2(n504), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U565 ( .A(G43GAT), .B(n503), .Z(G1330GAT) );
  XOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U567 ( .A1(n504), .A2(n527), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n510) );
  NOR2_X1 U570 ( .A1(n549), .A2(n565), .ZN(n507) );
  XOR2_X1 U571 ( .A(KEYINPUT106), .B(n507), .Z(n520) );
  NOR2_X1 U572 ( .A1(n520), .A2(n508), .ZN(n514) );
  NAND2_X1 U573 ( .A1(n514), .A2(n521), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n523), .A2(n514), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n514), .A2(n531), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U581 ( .A1(n514), .A2(n527), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT108), .Z(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n526) );
  NAND2_X1 U586 ( .A1(n521), .A2(n526), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n526), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n531), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT113), .Z(n534) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n546), .A2(n532), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n549), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  INV_X1 U601 ( .A(n565), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n541), .A2(n551), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n538) );
  NAND2_X1 U606 ( .A1(n541), .A2(n556), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U610 ( .A1(n541), .A2(n559), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n576), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT117), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n549), .A2(n560), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n555) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT118), .Z(n553) );
  NAND2_X1 U620 ( .A1(n560), .A2(n551), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT119), .Z(n558) );
  NAND2_X1 U624 ( .A1(n560), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  INV_X1 U628 ( .A(KEYINPUT120), .ZN(n563) );
  NOR2_X1 U629 ( .A1(n570), .A2(n578), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  NOR2_X1 U632 ( .A1(n570), .A2(n565), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n567) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NOR2_X1 U637 ( .A1(n588), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(n573), .ZN(G1350GAT) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n590) );
  NOR2_X1 U643 ( .A1(n578), .A2(n590), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(KEYINPUT60), .B(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n590), .ZN(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

