//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT0), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n192), .B2(new_n193), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n191), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n204), .A3(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT81), .ZN(new_n210));
  INV_X1    g024(.A(G224), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G953), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n200), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n210), .B2(new_n214), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G107), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(G107), .ZN(new_n224));
  OAI22_X1  g038(.A1(new_n218), .A2(G107), .B1(KEYINPUT74), .B2(KEYINPUT3), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G104), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n224), .A3(KEYINPUT75), .ZN(new_n229));
  OR3_X1    g043(.A1(new_n218), .A2(KEYINPUT75), .A3(G107), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G101), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G119), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT66), .A3(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(G119), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT67), .B1(new_n244), .B2(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n247));
  INV_X1    g061(.A(G113), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n234), .A2(G119), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT5), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n247), .B(new_n251), .C1(new_n244), .C2(new_n250), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n244), .B2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT79), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n232), .A2(new_n246), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G110), .B(G122), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n243), .A2(new_n245), .B1(new_n241), .B2(new_n244), .ZN(new_n257));
  INV_X1    g071(.A(new_n221), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n228), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n225), .A2(new_n224), .ZN(new_n261));
  OAI21_X1  g075(.A(G101), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(G101), .C1(new_n260), .C2(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n255), .B(new_n256), .C1(new_n257), .C2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n255), .B1(new_n257), .B2(new_n266), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n256), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n267), .A2(KEYINPUT6), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n268), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n217), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT7), .B1(new_n211), .B2(G953), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n200), .A2(new_n208), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n200), .B2(new_n208), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n256), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n243), .A2(new_n245), .B1(new_n281), .B2(new_n251), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n226), .A2(new_n231), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND4_X1   g098(.A1(new_n246), .A2(new_n283), .A3(new_n252), .A4(new_n254), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT83), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n246), .A2(new_n253), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n232), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n246), .A2(new_n283), .A3(new_n254), .A4(new_n252), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT83), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n280), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n278), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n273), .A2(new_n293), .A3(new_n295), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n189), .A2(G128), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n193), .A2(G143), .ZN(new_n303));
  INV_X1    g117(.A(G134), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G122), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G116), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n234), .A2(G122), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G107), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n227), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n305), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT13), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n193), .B2(G143), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n189), .A2(KEYINPUT13), .A3(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n303), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G134), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(new_n316), .B2(G134), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n312), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT86), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n312), .B(new_n322), .C1(new_n318), .C2(new_n319), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n304), .B1(new_n302), .B2(new_n303), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n311), .B1(new_n305), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT14), .ZN(new_n326));
  OAI21_X1  g140(.A(G107), .B1(new_n308), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n309), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n323), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT9), .B(G234), .ZN(new_n333));
  INV_X1    g147(.A(G217), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n333), .A2(new_n334), .A3(G953), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n321), .A2(new_n323), .A3(new_n331), .A4(new_n335), .ZN(new_n338));
  AOI21_X1  g152(.A(G902), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT15), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G478), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n301), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G902), .ZN(new_n343));
  INV_X1    g157(.A(new_n338), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n330), .B1(new_n320), .B2(KEYINPUT86), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n335), .B1(new_n345), .B2(new_n323), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n343), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(KEYINPUT87), .A3(new_n340), .A4(G478), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n343), .B(new_n341), .C1(new_n344), .C2(new_n346), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT88), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n338), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(KEYINPUT88), .A3(new_n343), .A4(new_n341), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n342), .A2(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n218), .ZN(new_n356));
  INV_X1    g170(.A(G140), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G125), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n207), .A2(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(G146), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G143), .A3(G214), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G143), .B1(new_n362), .B2(G214), .ZN(new_n365));
  OAI211_X1 g179(.A(KEYINPUT18), .B(G131), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(G214), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n189), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT18), .A2(G131), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n361), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G131), .B1(new_n364), .B2(new_n365), .ZN(new_n372));
  INV_X1    g186(.A(G131), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n373), .A3(new_n363), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT17), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT17), .B(G131), .C1(new_n364), .C2(new_n365), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT16), .ZN(new_n378));
  OR3_X1    g192(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n187), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n379), .A3(G146), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n356), .B(new_n371), .C1(new_n376), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n378), .A2(G146), .A3(new_n379), .ZN(new_n386));
  AOI21_X1  g200(.A(G146), .B1(new_n378), .B2(new_n379), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(new_n377), .C1(new_n375), .C2(KEYINPUT17), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n356), .B1(new_n389), .B2(new_n371), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n343), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G475), .ZN(new_n392));
  NAND2_X1  g206(.A1(G234), .A2(G237), .ZN(new_n393));
  INV_X1    g207(.A(G953), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(G952), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT21), .B(G898), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(G902), .A3(G953), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT89), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n358), .A2(new_n359), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n360), .B1(new_n405), .B2(KEYINPUT19), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n406), .A3(new_n187), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT71), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n378), .A2(new_n379), .A3(new_n409), .A4(G146), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n375), .A2(new_n407), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n371), .ZN(new_n412));
  INV_X1    g226(.A(new_n356), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n384), .ZN(new_n415));
  NOR2_X1   g229(.A1(G475), .A2(G902), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n401), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n416), .ZN(new_n418));
  AOI211_X1 g232(.A(KEYINPUT20), .B(new_n418), .C1(new_n414), .C2(new_n384), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n392), .B(new_n400), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n299), .A2(new_n300), .A3(new_n354), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G221), .ZN(new_n423));
  INV_X1    g237(.A(new_n333), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(new_n343), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n304), .B2(G137), .ZN(new_n428));
  INV_X1    g242(.A(G137), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT11), .A3(G134), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n304), .A2(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G131), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n428), .A2(new_n430), .A3(new_n373), .A4(new_n431), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(KEYINPUT64), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n436), .A3(G131), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AND4_X1   g252(.A1(new_n204), .A2(new_n188), .A3(new_n190), .A4(G128), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT76), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n201), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n188), .A2(KEYINPUT76), .A3(KEYINPUT1), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(G128), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n439), .B1(new_n443), .B2(new_n191), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n283), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n206), .B1(new_n226), .B2(new_n231), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n438), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT12), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n394), .A2(G227), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT72), .ZN(new_n450));
  XOR2_X1   g264(.A(G110), .B(G140), .Z(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n201), .A2(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n439), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n283), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n444), .B2(new_n283), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n438), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n263), .A2(new_n199), .A3(new_n265), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n444), .B2(new_n283), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n435), .A2(new_n437), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n206), .A2(KEYINPUT10), .A3(new_n226), .A4(new_n231), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n459), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n448), .A2(new_n452), .A3(new_n458), .A4(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n438), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n452), .B1(new_n467), .B2(new_n464), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n465), .B1(new_n468), .B2(KEYINPUT78), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n447), .A2(KEYINPUT12), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n457), .B1(new_n456), .B2(new_n438), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n452), .A4(new_n464), .ZN(new_n474));
  AOI211_X1 g288(.A(G469), .B(G902), .C1(new_n469), .C2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n448), .A2(new_n464), .A3(new_n458), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n452), .B(KEYINPUT73), .Z(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n467), .A2(new_n452), .A3(new_n464), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(G469), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(G469), .A2(G902), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n426), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n422), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n334), .B1(G234), .B2(new_n343), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT22), .B(G137), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n394), .A2(G221), .A3(G234), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n193), .A2(G119), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n236), .A2(G128), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT69), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G110), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G110), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT69), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n491), .A4(new_n492), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n236), .B2(G128), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n492), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G110), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n490), .B1(new_n509), .B2(new_n388), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n495), .A2(new_n502), .B1(G110), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n381), .A2(new_n382), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT70), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n493), .A2(new_n494), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n505), .A2(new_n506), .A3(new_n496), .A4(new_n492), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n515), .A2(new_n516), .B1(new_n402), .B2(new_n187), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n517), .A2(new_n408), .A3(new_n410), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n489), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  AOI211_X1 g334(.A(new_n488), .B(new_n518), .C1(new_n510), .C2(new_n513), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT25), .B1(new_n522), .B2(new_n343), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n509), .A2(new_n388), .A3(new_n490), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT70), .B1(new_n511), .B2(new_n512), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n488), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n514), .A2(new_n519), .A3(new_n489), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n527), .A2(KEYINPUT25), .A3(new_n343), .A4(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n485), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n522), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n485), .A2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n362), .A2(G210), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT27), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT26), .B(G101), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n304), .A2(G137), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n429), .A2(G134), .ZN(new_n543));
  OAI21_X1  g357(.A(G131), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n434), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT68), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n434), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n206), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n435), .A2(new_n437), .A3(new_n199), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n257), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT28), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n549), .A2(new_n550), .A3(new_n257), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(KEYINPUT65), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT65), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n435), .A2(new_n199), .A3(new_n557), .A4(new_n437), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n454), .A2(new_n545), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n257), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n541), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT30), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n562), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n551), .A2(new_n541), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT31), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n559), .B1(new_n550), .B2(KEYINPUT65), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT30), .B1(new_n574), .B2(new_n558), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT31), .B(new_n572), .C1(new_n575), .C2(new_n569), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n565), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n579));
  NOR2_X1   g393(.A1(G472), .A2(G902), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n572), .B1(new_n575), .B2(new_n569), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n564), .B1(new_n584), .B2(new_n576), .ZN(new_n585));
  INV_X1    g399(.A(new_n580), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT32), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n549), .A2(new_n550), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n562), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n555), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n541), .A2(KEYINPUT29), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n541), .B1(new_n571), .B2(new_n551), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n555), .A2(new_n563), .A3(new_n541), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI221_X1 g410(.A(new_n343), .B1(new_n591), .B2(new_n592), .C1(new_n593), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n537), .B1(new_n588), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n484), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND3_X1  g415(.A1(new_n527), .A2(new_n343), .A3(new_n528), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT25), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n529), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n535), .B1(new_n605), .B2(new_n485), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n426), .C1(new_n475), .C2(new_n482), .ZN(new_n607));
  OAI21_X1  g421(.A(G472), .B1(new_n585), .B2(G902), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n578), .A2(new_n580), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n273), .A2(new_n293), .A3(new_n295), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n295), .B1(new_n273), .B2(new_n293), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n300), .B(new_n400), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n338), .B2(KEYINPUT90), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n352), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n337), .B(new_n338), .C1(KEYINPUT90), .C2(new_n615), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(G478), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G478), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n343), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n339), .B2(new_n620), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n392), .B1(new_n417), .B2(new_n419), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n614), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n611), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NAND2_X1  g443(.A1(new_n342), .A2(new_n348), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n351), .A2(new_n353), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n392), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n356), .B1(new_n411), .B2(new_n371), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n416), .B1(new_n385), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT20), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(KEYINPUT91), .A3(new_n419), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n415), .A2(new_n401), .A3(new_n416), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT91), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n638), .B1(new_n417), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n633), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n614), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n611), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  OAI21_X1  g460(.A(new_n300), .B1(new_n612), .B2(new_n613), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n354), .A2(new_n421), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(G902), .B1(new_n469), .B2(new_n474), .ZN(new_n650));
  INV_X1    g464(.A(G469), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n482), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n425), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n608), .A2(new_n609), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n526), .B(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n534), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n531), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n649), .A2(new_n654), .A3(new_n655), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  OR2_X1    g477(.A1(new_n398), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n395), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n632), .A2(new_n641), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT92), .B1(new_n666), .B2(new_n647), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n419), .B1(new_n636), .B2(KEYINPUT91), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n635), .A2(new_n639), .A3(KEYINPUT20), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n392), .B(new_n665), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n354), .ZN(new_n671));
  INV_X1    g485(.A(new_n300), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n297), .B2(new_n298), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT92), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n482), .B1(new_n650), .B2(new_n651), .ZN(new_n676));
  INV_X1    g490(.A(new_n485), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n604), .B2(new_n529), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n658), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n676), .A2(new_n679), .A3(new_n425), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n588), .A2(new_n598), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n667), .A2(new_n675), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  INV_X1    g497(.A(new_n624), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n660), .A2(new_n672), .A3(new_n354), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT94), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT93), .B(KEYINPUT38), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n299), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n582), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n541), .B1(new_n590), .B2(new_n551), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n343), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G472), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n579), .B1(new_n578), .B2(new_n580), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n585), .A2(KEYINPUT32), .A3(new_n586), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n685), .A2(new_n686), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n690), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n665), .B(KEYINPUT39), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n654), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT40), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n189), .ZN(G45));
  AND4_X1   g518(.A1(new_n624), .A2(new_n619), .A3(new_n622), .A4(new_n665), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n680), .A2(new_n681), .A3(new_n673), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  NAND2_X1  g521(.A1(new_n469), .A2(new_n474), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n343), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT95), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n650), .B2(new_n651), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n709), .A2(new_n711), .A3(G469), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n425), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n599), .A3(new_n626), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n714), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n599), .A2(new_n719), .A3(new_n426), .A4(new_n643), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  OAI211_X1 g535(.A(new_n354), .B(new_n421), .C1(new_n678), .C2(new_n658), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n588), .B2(new_n598), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n715), .A2(new_n673), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  INV_X1    g539(.A(new_n614), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n573), .A2(new_n577), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n541), .B1(new_n555), .B2(new_n590), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n580), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n606), .A2(new_n729), .A3(new_n608), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n632), .A2(KEYINPUT96), .A3(new_n624), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT96), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n354), .B2(new_n684), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n715), .A2(new_n726), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  AND4_X1   g550(.A1(new_n608), .A2(new_n660), .A3(new_n705), .A4(new_n729), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n719), .A2(new_n737), .A3(new_n426), .A4(new_n673), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT97), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n478), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n476), .A2(KEYINPUT97), .A3(new_n477), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(G469), .A3(new_n479), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n481), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n426), .B1(new_n744), .B2(new_n475), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n297), .A2(new_n300), .A3(new_n298), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n599), .A3(new_n705), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n747), .A2(new_n599), .A3(KEYINPUT42), .A4(new_n705), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NAND3_X1  g567(.A1(new_n747), .A2(new_n599), .A3(new_n671), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT98), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT98), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n747), .A2(new_n599), .A3(new_n756), .A4(new_n671), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND2_X1  g573(.A1(new_n742), .A2(new_n479), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT97), .B1(new_n476), .B2(new_n477), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT45), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n478), .B2(new_n479), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n651), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n481), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n652), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n426), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n700), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n623), .A2(new_n684), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT43), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT43), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n610), .B(new_n660), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n775), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n746), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n782), .B2(new_n783), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n772), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT47), .B(new_n426), .C1(new_n770), .C2(new_n771), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n537), .A2(new_n705), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n681), .A2(new_n746), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT100), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(KEYINPUT100), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  INV_X1    g615(.A(new_n719), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n776), .A2(new_n537), .A3(new_n425), .A4(new_n672), .ZN(new_n804));
  INV_X1    g618(.A(new_n697), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n689), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n719), .A2(new_n426), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n809), .A2(KEYINPUT109), .A3(new_n300), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT109), .B1(new_n809), .B2(new_n300), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n689), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT110), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT110), .ZN(new_n814));
  INV_X1    g628(.A(new_n395), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n777), .A2(new_n815), .A3(new_n778), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT107), .Z(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n730), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(KEYINPUT50), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n819), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n425), .B1(new_n802), .B2(KEYINPUT108), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(KEYINPUT108), .B2(new_n802), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n818), .B(new_n786), .C1(new_n793), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n809), .A2(new_n746), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n805), .A2(new_n606), .A3(new_n815), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n623), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n684), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n660), .A2(new_n608), .A3(new_n729), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n817), .A2(KEYINPUT112), .A3(new_n826), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT112), .B1(new_n817), .B2(new_n826), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n832), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT51), .B1(new_n822), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n599), .B1(new_n835), .B2(new_n836), .ZN(new_n843));
  XOR2_X1   g657(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n818), .A2(new_n673), .A3(new_n715), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(G952), .A3(new_n394), .ZN(new_n847));
  INV_X1    g661(.A(new_n625), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n829), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n842), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT105), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n738), .A2(new_n682), .A3(new_n706), .ZN(new_n854));
  OAI21_X1  g668(.A(G469), .B1(new_n762), .B2(G902), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n425), .B1(new_n855), .B2(new_n652), .ZN(new_n856));
  INV_X1    g670(.A(new_n665), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n660), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n697), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n734), .A2(new_n673), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT103), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n745), .A2(new_n660), .A3(new_n857), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n647), .B1(new_n731), .B2(new_n733), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT103), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n697), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n854), .A2(new_n866), .A3(KEYINPUT52), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT52), .B1(new_n854), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n680), .A2(new_n681), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n746), .A2(new_n632), .A3(new_n670), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n871), .A2(new_n872), .B1(new_n737), .B2(new_n747), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n752), .A2(new_n758), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n676), .A2(new_n537), .A3(new_n425), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n632), .A2(new_n684), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n614), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n877), .A3(new_n655), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT101), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n878), .A2(new_n661), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n878), .B2(new_n661), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n484), .A2(new_n599), .B1(new_n611), .B2(new_n626), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n715), .B(new_n599), .C1(new_n626), .C2(new_n643), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n724), .A4(new_n735), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT102), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n354), .A2(new_n624), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n673), .A2(new_n400), .A3(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n889), .A2(new_n607), .A3(new_n610), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n660), .A2(new_n609), .A3(new_n608), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n422), .A2(new_n891), .A3(new_n483), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT101), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n878), .A2(new_n661), .A3(new_n879), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n716), .A2(new_n724), .A3(new_n720), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n730), .A2(new_n734), .A3(new_n726), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n809), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n681), .A2(new_n606), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n654), .A2(new_n673), .A3(new_n354), .A4(new_n421), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n655), .A2(new_n654), .A3(new_n606), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n848), .A2(new_n673), .A3(new_n400), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n899), .A2(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n895), .A2(new_n896), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n752), .A2(new_n758), .A3(new_n873), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT102), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n870), .B1(new_n887), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n853), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n869), .A2(KEYINPUT104), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT104), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n868), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n887), .A2(new_n908), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n874), .A2(new_n886), .A3(KEYINPUT102), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n869), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(KEYINPUT105), .A3(KEYINPUT53), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n911), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n909), .A2(KEYINPUT106), .A3(new_n910), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT106), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n920), .B2(KEYINPUT53), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n905), .A2(new_n906), .A3(new_n910), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n912), .A2(new_n914), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n822), .A2(new_n841), .A3(KEYINPUT51), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n852), .A2(new_n923), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT115), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(G952), .A2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT116), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n933), .B2(new_n934), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n808), .B1(new_n935), .B2(new_n938), .ZN(G75));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n343), .B1(new_n927), .B2(new_n930), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(G210), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n271), .A2(new_n272), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n217), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT55), .Z(new_n947));
  AND2_X1   g761(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n944), .A2(new_n947), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n394), .A2(G952), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(G51));
  NOR2_X1   g765(.A1(new_n942), .A2(new_n766), .ZN(new_n952));
  INV_X1    g766(.A(new_n708), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT106), .B1(new_n909), .B2(new_n910), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n920), .A2(new_n925), .A3(KEYINPUT53), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n930), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT54), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n931), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n481), .B(KEYINPUT57), .Z(new_n959));
  AOI21_X1  g773(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT117), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n952), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n959), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n957), .B2(new_n931), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT117), .B1(new_n964), .B2(new_n953), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n950), .B1(new_n962), .B2(new_n965), .ZN(G54));
  INV_X1    g780(.A(KEYINPUT118), .ZN(new_n967));
  NAND2_X1  g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n956), .A2(G902), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n415), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n950), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n941), .A2(KEYINPUT118), .A3(new_n415), .A4(new_n969), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT119), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT119), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n972), .A2(new_n973), .A3(new_n977), .A4(new_n974), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(G60));
  NAND2_X1  g793(.A1(new_n617), .A2(new_n618), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n923), .A2(new_n931), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n621), .B(KEYINPUT59), .Z(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n980), .A2(new_n982), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n950), .B(new_n983), .C1(new_n958), .C2(new_n984), .ZN(G63));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT60), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n956), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n532), .ZN(new_n989));
  INV_X1    g803(.A(new_n950), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n657), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n956), .A2(new_n992), .A3(new_n987), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT120), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n991), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT121), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n989), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n988), .A2(KEYINPUT121), .A3(new_n532), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n999), .A2(KEYINPUT61), .A3(new_n990), .A4(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n993), .B(KEYINPUT120), .ZN(new_n1002));
  OAI22_X1  g816(.A1(new_n997), .A2(KEYINPUT61), .B1(new_n1001), .B2(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n396), .B2(new_n211), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n886), .B2(G953), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n945), .B1(G898), .B2(new_n394), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G69));
  NAND2_X1  g821(.A1(new_n567), .A2(new_n568), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n404), .A2(new_n406), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G900), .A2(G953), .ZN(new_n1011));
  INV_X1    g825(.A(new_n788), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n774), .A2(new_n899), .A3(new_n860), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n854), .B(KEYINPUT122), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n752), .A2(new_n758), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT124), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1014), .A2(new_n800), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1010), .B(new_n1011), .C1(new_n1018), .C2(G953), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1015), .B1(new_n702), .B2(new_n699), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n746), .B1(new_n625), .B2(new_n876), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n599), .A2(new_n1022), .A3(new_n654), .A4(new_n700), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1021), .A2(new_n788), .A3(new_n800), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1025));
  OAI21_X1  g839(.A(KEYINPUT123), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1023), .B1(new_n785), .B2(new_n787), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1027), .B1(new_n798), .B2(new_n799), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT123), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1025), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1021), .ZN(new_n1031));
  AOI21_X1  g845(.A(G953), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1019), .B1(new_n1032), .B2(new_n1010), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n394), .B1(G227), .B2(G900), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1033), .B(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  OAI21_X1  g851(.A(new_n1037), .B1(new_n1018), .B2(new_n905), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n571), .A2(new_n551), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT125), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1040), .A2(new_n541), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n950), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1040), .A2(new_n541), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1026), .A2(new_n1031), .A3(new_n886), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1043), .B1(new_n1044), .B2(new_n1037), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT126), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g861(.A(KEYINPUT126), .B(new_n1043), .C1(new_n1044), .C2(new_n1037), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n922), .B(new_n1037), .C1(new_n691), .C2(new_n593), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT127), .Z(new_n1051));
  NOR2_X1   g865(.A1(new_n1049), .A2(new_n1051), .ZN(G57));
endmodule


