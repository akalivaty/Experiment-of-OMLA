

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XOR2_X1 U324 ( .A(n456), .B(KEYINPUT41), .Z(n565) );
  INV_X1 U325 ( .A(KEYINPUT47), .ZN(n399) );
  XNOR2_X1 U326 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U327 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n427) );
  XNOR2_X1 U328 ( .A(n402), .B(n401), .ZN(n410) );
  XNOR2_X1 U329 ( .A(n428), .B(n427), .ZN(n449) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n453) );
  XNOR2_X1 U331 ( .A(n453), .B(KEYINPUT58), .ZN(n454) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n293) );
  XNOR2_X1 U334 ( .A(G134GAT), .B(G106GAT), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n309) );
  XOR2_X1 U336 ( .A(G50GAT), .B(G162GAT), .Z(n332) );
  XOR2_X1 U337 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n295) );
  XNOR2_X1 U338 ( .A(KEYINPUT9), .B(KEYINPUT77), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U340 ( .A(n332), .B(n296), .Z(n298) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U343 ( .A(KEYINPUT72), .B(G85GAT), .Z(n300) );
  XNOR2_X1 U344 ( .A(G99GAT), .B(KEYINPUT71), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U346 ( .A(G92GAT), .B(n301), .Z(n384) );
  XOR2_X1 U347 ( .A(n302), .B(n384), .Z(n307) );
  XOR2_X1 U348 ( .A(G29GAT), .B(G43GAT), .Z(n304) );
  XNOR2_X1 U349 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n368) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n305), .B(G218GAT), .ZN(n414) );
  XNOR2_X1 U353 ( .A(n368), .B(n414), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n556) );
  XOR2_X1 U356 ( .A(G176GAT), .B(G183GAT), .Z(n311) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n320) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n313) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n422) );
  XOR2_X1 U362 ( .A(n422), .B(G71GAT), .Z(n315) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U365 ( .A(G15GAT), .B(G127GAT), .Z(n346) );
  XOR2_X1 U366 ( .A(n316), .B(n346), .Z(n318) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G190GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U370 ( .A(KEYINPUT82), .B(G134GAT), .Z(n322) );
  XNOR2_X1 U371 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U373 ( .A(G113GAT), .B(n323), .Z(n436) );
  XOR2_X2 U374 ( .A(n324), .B(n436), .Z(n530) );
  XOR2_X1 U375 ( .A(G211GAT), .B(KEYINPUT24), .Z(n326) );
  XNOR2_X1 U376 ( .A(G218GAT), .B(KEYINPUT86), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(G197GAT), .B(KEYINPUT21), .Z(n413) );
  XOR2_X1 U379 ( .A(n327), .B(n413), .Z(n335) );
  XOR2_X1 U380 ( .A(G148GAT), .B(G204GAT), .Z(n329) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n385) );
  XOR2_X1 U383 ( .A(n385), .B(KEYINPUT22), .Z(n331) );
  NAND2_X1 U384 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U388 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n337) );
  XNOR2_X1 U389 ( .A(KEYINPUT23), .B(KEYINPUT83), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n344) );
  XNOR2_X1 U392 ( .A(G22GAT), .B(G155GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n340), .B(G78GAT), .ZN(n358) );
  XOR2_X1 U394 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n342) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(KEYINPUT84), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n435) );
  XNOR2_X1 U397 ( .A(n358), .B(n435), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n465) );
  XNOR2_X1 U399 ( .A(G71GAT), .B(G57GAT), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n345), .B(KEYINPUT13), .ZN(n382) );
  XNOR2_X1 U401 ( .A(n382), .B(n346), .ZN(n348) );
  AND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U404 ( .A(n349), .B(KEYINPUT80), .Z(n351) );
  XOR2_X1 U405 ( .A(KEYINPUT68), .B(G1GAT), .Z(n364) );
  XNOR2_X1 U406 ( .A(n364), .B(G64GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U408 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n353) );
  XNOR2_X1 U409 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT78), .B(G211GAT), .Z(n357) );
  XNOR2_X1 U413 ( .A(G8GAT), .B(G183GAT), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n421) );
  XNOR2_X1 U415 ( .A(n358), .B(n421), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n583) );
  XNOR2_X1 U417 ( .A(n583), .B(KEYINPUT110), .ZN(n569) );
  XOR2_X1 U418 ( .A(G113GAT), .B(G36GAT), .Z(n362) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G50GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n366) );
  AND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U424 ( .A(KEYINPUT66), .B(n367), .Z(n370) );
  XNOR2_X1 U425 ( .A(n368), .B(KEYINPUT30), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n406) );
  XOR2_X1 U427 ( .A(G197GAT), .B(G141GAT), .Z(n372) );
  XNOR2_X1 U428 ( .A(G15GAT), .B(G22GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U430 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n374) );
  XNOR2_X1 U431 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U433 ( .A(n376), .B(n375), .Z(n405) );
  XNOR2_X1 U434 ( .A(n406), .B(n405), .ZN(n560) );
  XOR2_X1 U435 ( .A(G176GAT), .B(G64GAT), .Z(n412) );
  XOR2_X1 U436 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n378) );
  XNOR2_X1 U437 ( .A(G120GAT), .B(G78GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n412), .B(n379), .ZN(n381) );
  NAND2_X1 U440 ( .A1(G230GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U445 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n389) );
  XNOR2_X1 U446 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  NAND2_X1 U448 ( .A1(n391), .A2(n390), .ZN(n395) );
  INV_X1 U449 ( .A(n390), .ZN(n393) );
  INV_X1 U450 ( .A(n391), .ZN(n392) );
  NAND2_X1 U451 ( .A1(n393), .A2(n392), .ZN(n394) );
  NAND2_X1 U452 ( .A1(n395), .A2(n394), .ZN(n456) );
  NOR2_X1 U453 ( .A1(n560), .A2(n565), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n396), .B(KEYINPUT46), .ZN(n397) );
  NOR2_X1 U455 ( .A1(n569), .A2(n397), .ZN(n398) );
  INV_X1 U456 ( .A(n556), .ZN(n545) );
  NAND2_X1 U457 ( .A1(n398), .A2(n545), .ZN(n402) );
  XOR2_X1 U458 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n400) );
  XNOR2_X1 U459 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n404) );
  XOR2_X1 U460 ( .A(KEYINPUT36), .B(n556), .Z(n588) );
  INV_X1 U461 ( .A(n583), .ZN(n489) );
  NOR2_X1 U462 ( .A1(n588), .A2(n489), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n407) );
  XOR2_X1 U464 ( .A(n406), .B(n405), .Z(n575) );
  NOR2_X1 U465 ( .A1(n407), .A2(n575), .ZN(n408) );
  NAND2_X1 U466 ( .A1(n456), .A2(n408), .ZN(n409) );
  NAND2_X1 U467 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n411), .B(KEYINPUT48), .ZN(n528) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n426) );
  XOR2_X1 U470 ( .A(n414), .B(KEYINPUT93), .Z(n416) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U473 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n418) );
  XNOR2_X1 U474 ( .A(G204GAT), .B(G92GAT), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U476 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(n426), .B(n425), .Z(n519) );
  INV_X1 U480 ( .A(n519), .ZN(n460) );
  NAND2_X1 U481 ( .A1(n528), .A2(n460), .ZN(n428) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n434) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G148GAT), .Z(n430) );
  XNOR2_X1 U484 ( .A(G127GAT), .B(G155GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U486 ( .A(G29GAT), .B(G162GAT), .Z(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n448) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n438) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n446) );
  XOR2_X1 U492 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n440) );
  XNOR2_X1 U493 ( .A(KEYINPUT88), .B(KEYINPUT6), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n442) );
  XNOR2_X1 U496 ( .A(G1GAT), .B(G57GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U500 ( .A(n448), .B(n447), .Z(n471) );
  INV_X1 U501 ( .A(n471), .ZN(n517) );
  NAND2_X1 U502 ( .A1(n449), .A2(n517), .ZN(n572) );
  NOR2_X1 U503 ( .A1(n465), .A2(n572), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U505 ( .A1(n530), .A2(n451), .ZN(n452) );
  XNOR2_X1 U506 ( .A(KEYINPUT122), .B(n452), .ZN(n570) );
  AND2_X1 U507 ( .A1(n556), .A2(n570), .ZN(n455) );
  INV_X1 U508 ( .A(n456), .ZN(n579) );
  NOR2_X1 U509 ( .A1(n579), .A2(n560), .ZN(n491) );
  INV_X1 U510 ( .A(n530), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n465), .B(KEYINPUT65), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n457), .B(KEYINPUT28), .ZN(n532) );
  XNOR2_X1 U513 ( .A(n519), .B(KEYINPUT27), .ZN(n467) );
  NOR2_X1 U514 ( .A1(n467), .A2(n517), .ZN(n529) );
  NAND2_X1 U515 ( .A1(n532), .A2(n529), .ZN(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT95), .B(n458), .Z(n459) );
  NOR2_X1 U517 ( .A1(n461), .A2(n459), .ZN(n473) );
  NAND2_X1 U518 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U519 ( .A(KEYINPUT96), .B(n462), .Z(n463) );
  NOR2_X1 U520 ( .A1(n465), .A2(n463), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n464), .Z(n469) );
  NAND2_X1 U522 ( .A1(n530), .A2(n465), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT26), .ZN(n573) );
  NOR2_X1 U524 ( .A1(n573), .A2(n467), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n487) );
  XOR2_X1 U528 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n475) );
  NAND2_X1 U529 ( .A1(n545), .A2(n583), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n487), .A2(n476), .ZN(n477) );
  XOR2_X1 U532 ( .A(KEYINPUT97), .B(n477), .Z(n502) );
  NAND2_X1 U533 ( .A1(n491), .A2(n502), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT98), .ZN(n485) );
  NOR2_X1 U535 ( .A1(n485), .A2(n517), .ZN(n480) );
  XNOR2_X1 U536 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U539 ( .A1(n485), .A2(n519), .ZN(n482) );
  XOR2_X1 U540 ( .A(G8GAT), .B(n482), .Z(G1325GAT) );
  NOR2_X1 U541 ( .A1(n485), .A2(n530), .ZN(n484) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n532), .A2(n485), .ZN(n486) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n486), .Z(G1327GAT) );
  NOR2_X1 U546 ( .A1(n588), .A2(n487), .ZN(n488) );
  NAND2_X1 U547 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n490), .ZN(n516) );
  NAND2_X1 U549 ( .A1(n516), .A2(n491), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n492), .B(KEYINPUT38), .ZN(n500) );
  NOR2_X1 U551 ( .A1(n517), .A2(n500), .ZN(n496) );
  XOR2_X1 U552 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n494) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n500), .A2(n519), .ZN(n497) );
  XOR2_X1 U557 ( .A(G36GAT), .B(n497), .Z(G1329GAT) );
  NOR2_X1 U558 ( .A1(n500), .A2(n530), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(n498), .Z(n499) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n532), .A2(n500), .ZN(n501) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  NOR2_X1 U563 ( .A1(n565), .A2(n575), .ZN(n515) );
  NAND2_X1 U564 ( .A1(n515), .A2(n502), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(KEYINPUT102), .ZN(n511) );
  NOR2_X1 U566 ( .A1(n511), .A2(n517), .ZN(n505) );
  XNOR2_X1 U567 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n511), .A2(n519), .ZN(n507) );
  XOR2_X1 U571 ( .A(KEYINPUT104), .B(n507), .Z(n508) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n511), .A2(n530), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n513) );
  NOR2_X1 U577 ( .A1(n532), .A2(n511), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n525) );
  NOR2_X1 U581 ( .A1(n517), .A2(n525), .ZN(n518) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n525), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n530), .A2(n525), .ZN(n522) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n532), .A2(n525), .ZN(n526) );
  XOR2_X1 U592 ( .A(n527), .B(n526), .Z(G1339GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n529), .ZN(n548) );
  NOR2_X1 U594 ( .A1(n530), .A2(n548), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(n531), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n544) );
  NOR2_X1 U597 ( .A1(n560), .A2(n544), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  NOR2_X1 U601 ( .A1(n565), .A2(n544), .ZN(n538) );
  XNOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n542) );
  INV_X1 U606 ( .A(n544), .ZN(n540) );
  NAND2_X1 U607 ( .A1(n540), .A2(n569), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U609 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  NOR2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n573), .A2(n548), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n575), .A2(n557), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  INV_X1 U617 ( .A(n565), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n557), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  XOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U622 ( .A1(n557), .A2(n583), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(KEYINPUT120), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  INV_X1 U627 ( .A(n570), .ZN(n566) );
  NOR2_X1 U628 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(G169GAT), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT123), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n564) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U633 ( .A(n564), .B(n563), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U635 ( .A(n568), .B(n567), .Z(G1349GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT125), .B(n574), .ZN(n587) );
  INV_X1 U641 ( .A(n587), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U646 ( .A1(n584), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

