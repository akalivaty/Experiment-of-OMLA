//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT90), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G237), .ZN(new_n203));
  INV_X1    g017(.A(G953), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G214), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT64), .A2(G143), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT18), .A2(G131), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n203), .A2(new_n204), .A3(G143), .A4(G214), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n202), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n209), .ZN(new_n215));
  INV_X1    g029(.A(G214), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n216), .A2(G237), .A3(G953), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n211), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT89), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n222), .A3(new_n219), .ZN(new_n223));
  AOI211_X1 g037(.A(new_n192), .B(new_n214), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n223), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n202), .A2(new_n213), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT90), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n218), .A2(G131), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n210), .B2(new_n212), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n197), .B(KEYINPUT19), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n229), .A2(new_n231), .B1(new_n232), .B2(G146), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT16), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n193), .A3(G125), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT80), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT80), .B1(new_n199), .B2(KEYINPUT16), .ZN(new_n238));
  INV_X1    g052(.A(new_n235), .ZN(new_n239));
  OAI211_X1 g053(.A(G146), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n187), .B(new_n191), .C1(new_n228), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n223), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n222), .B1(new_n218), .B2(new_n219), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n226), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n192), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n225), .A2(KEYINPUT90), .A3(new_n226), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n242), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT91), .B1(new_n249), .B2(new_n190), .ZN(new_n250));
  OR3_X1    g064(.A1(new_n229), .A2(KEYINPUT17), .A3(new_n231), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n231), .A2(KEYINPUT17), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n197), .B2(new_n234), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n236), .B1(new_n255), .B2(new_n235), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT81), .A3(G146), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n240), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n200), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n247), .A2(new_n248), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n190), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n243), .A2(new_n250), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT20), .ZN(new_n267));
  NOR2_X1   g081(.A1(G475), .A2(G902), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT92), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT92), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n266), .A2(new_n271), .A3(new_n267), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n268), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G475), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n263), .A2(new_n264), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n191), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n265), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n204), .A2(G952), .ZN(new_n285));
  INV_X1    g099(.A(G234), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n203), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT21), .B(G898), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT96), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT77), .B(G902), .Z(new_n292));
  AOI211_X1 g106(.A(new_n204), .B(new_n292), .C1(G234), .C2(G237), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G478), .ZN(new_n296));
  NOR2_X1   g110(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G116), .B(G122), .ZN(new_n302));
  INV_X1    g116(.A(G107), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT14), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G122), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G116), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n303), .B1(new_n308), .B2(KEYINPUT14), .ZN(new_n309));
  AOI22_X1  g123(.A1(KEYINPUT94), .A2(new_n304), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n208), .A2(G128), .A3(new_n209), .ZN(new_n311));
  INV_X1    g125(.A(G134), .ZN(new_n312));
  INV_X1    g126(.A(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G143), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n311), .B2(new_n314), .ZN(new_n317));
  OAI221_X1 g131(.A(new_n310), .B1(KEYINPUT94), .B2(new_n304), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n315), .B(KEYINPUT93), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n302), .B(new_n303), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n311), .A2(KEYINPUT13), .A3(new_n314), .ZN(new_n321));
  OAI21_X1  g135(.A(G134), .B1(new_n311), .B2(KEYINPUT13), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n318), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT9), .B(G234), .ZN(new_n325));
  INV_X1    g139(.A(G217), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(G953), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n318), .B(new_n327), .C1(new_n319), .C2(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n301), .B1(new_n331), .B2(new_n292), .ZN(new_n332));
  INV_X1    g146(.A(new_n292), .ZN(new_n333));
  AOI211_X1 g147(.A(new_n333), .B(new_n300), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n277), .A2(new_n284), .A3(new_n295), .A4(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT86), .B(G469), .Z(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G140), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n204), .A2(G227), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n189), .B2(G107), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n303), .A2(KEYINPUT3), .A3(G104), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G101), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n303), .B2(G104), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n189), .A2(KEYINPUT82), .A3(G107), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n345), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n189), .A2(G107), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n303), .A2(G104), .ZN(new_n352));
  OAI21_X1  g166(.A(G101), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT84), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n356));
  AOI21_X1  g170(.A(G146), .B1(new_n208), .B2(new_n209), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n200), .A2(G143), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT1), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G143), .B2(new_n200), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n357), .A2(new_n358), .B1(new_n313), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n208), .A2(G146), .A3(new_n209), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n200), .A2(G143), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n313), .A2(KEYINPUT1), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n356), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n350), .A2(new_n367), .A3(new_n353), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n355), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT85), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n355), .A2(new_n366), .A3(new_n371), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G128), .B1(new_n357), .B2(new_n359), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n362), .A2(new_n363), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n362), .A2(new_n377), .A3(new_n363), .A4(new_n364), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n365), .A2(KEYINPUT83), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n354), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT10), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n303), .A2(KEYINPUT3), .A3(G104), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n303), .B2(G104), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n348), .B(new_n349), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n387));
  AND2_X1   g201(.A1(KEYINPUT0), .A2(G128), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n362), .A2(new_n363), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT0), .B(G128), .ZN(new_n390));
  AND2_X1   g204(.A1(KEYINPUT64), .A2(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(KEYINPUT64), .A2(G143), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n200), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n358), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n385), .A2(new_n397), .A3(G101), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n387), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n382), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n373), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n312), .A2(G137), .ZN(new_n402));
  INV_X1    g216(.A(G137), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT66), .B1(new_n403), .B2(G134), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT11), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT66), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n312), .B2(G137), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT11), .ZN(new_n409));
  OAI21_X1  g223(.A(G131), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(KEYINPUT11), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n405), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n230), .A4(new_n402), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(KEYINPUT67), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(G131), .C1(new_n406), .C2(new_n409), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n401), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n373), .A2(new_n400), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n341), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n374), .A2(new_n375), .B1(new_n365), .B2(KEYINPUT83), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n354), .B1(new_n422), .B2(new_n378), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n361), .A2(new_n365), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n381), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n417), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n417), .B(KEYINPUT12), .C1(new_n423), .C2(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n430), .A2(new_n420), .A3(new_n341), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n292), .B(new_n337), .C1(new_n421), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n420), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n340), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n418), .A2(new_n420), .A3(new_n341), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(KEYINPUT2), .A2(G113), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT2), .A2(G113), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT69), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT2), .A3(G113), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n447));
  XNOR2_X1  g261(.A(G116), .B(G119), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n450));
  INV_X1    g264(.A(new_n448), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n451), .B1(new_n446), .B2(new_n452), .ZN(new_n453));
  AOI211_X1 g267(.A(KEYINPUT70), .B(new_n441), .C1(new_n443), .C2(new_n445), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n449), .A2(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n398), .A3(new_n387), .ZN(new_n456));
  INV_X1    g270(.A(G119), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G116), .ZN(new_n458));
  OAI21_X1  g272(.A(G113), .B1(new_n458), .B2(KEYINPUT5), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(KEYINPUT5), .B2(new_n448), .ZN(new_n460));
  INV_X1    g274(.A(new_n441), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n444), .B1(KEYINPUT2), .B2(G113), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n442), .A2(KEYINPUT69), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n448), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT71), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n355), .A3(new_n368), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n456), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  OAI21_X1  g285(.A(G125), .B1(new_n389), .B2(new_n395), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n361), .A2(new_n195), .A3(new_n365), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n390), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n357), .B2(new_n358), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n362), .A2(new_n363), .A3(new_n388), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT87), .B1(new_n478), .B2(G125), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n480));
  INV_X1    g294(.A(G224), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(G953), .ZN(new_n482));
  OAI22_X1  g296(.A1(new_n474), .A2(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n449), .A2(new_n450), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n381), .B1(new_n484), .B2(new_n460), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n467), .A2(new_n354), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n469), .B(KEYINPUT8), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n470), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n472), .A2(new_n473), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT87), .ZN(new_n491));
  INV_X1    g305(.A(new_n479), .ZN(new_n492));
  INV_X1    g306(.A(new_n482), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n491), .A2(KEYINPUT7), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n456), .A2(new_n468), .ZN(new_n496));
  INV_X1    g310(.A(new_n469), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n491), .A2(new_n493), .A3(new_n492), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n482), .B1(new_n474), .B2(new_n479), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n503), .A3(new_n497), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n495), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n495), .A2(new_n505), .A3(new_n507), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n440), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n325), .B2(G902), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n438), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n336), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n455), .A2(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n414), .A2(new_n416), .A3(new_n396), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n465), .A2(new_n466), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT70), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n446), .A2(new_n452), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n451), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n312), .A2(G137), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n524), .B(G131), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n424), .A2(new_n413), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n515), .A2(new_n516), .A3(new_n523), .A4(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n455), .A2(KEYINPUT72), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n522), .B1(new_n517), .B2(new_n521), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n516), .A2(new_n528), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT65), .B1(new_n389), .B2(new_n395), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT65), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n476), .A2(new_n537), .A3(new_n477), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n414), .A2(new_n536), .A3(new_n416), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n528), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n534), .A2(new_n535), .B1(new_n540), .B2(new_n455), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n531), .B1(new_n541), .B2(new_n530), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n543));
  NAND3_X1  g357(.A1(new_n203), .A2(new_n204), .A3(G210), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT26), .B(G101), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n516), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n424), .A2(new_n413), .A3(new_n527), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n389), .A2(new_n395), .A3(KEYINPUT65), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n537), .B1(new_n476), .B2(new_n477), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n417), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n455), .B(new_n550), .C1(new_n555), .C2(KEYINPUT30), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n547), .B1(new_n556), .B2(new_n529), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n549), .A2(KEYINPUT29), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n531), .A2(KEYINPUT76), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n534), .A2(new_n535), .ZN(new_n560));
  INV_X1    g374(.A(new_n529), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT28), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n531), .A2(KEYINPUT76), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n547), .A2(KEYINPUT29), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n292), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G472), .B1(new_n558), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G472), .A2(G902), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT30), .B1(new_n539), .B2(new_n528), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n516), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n571));
  INV_X1    g385(.A(new_n455), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n529), .A2(KEYINPUT74), .A3(new_n547), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT31), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n529), .A2(new_n547), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT74), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n529), .A2(KEYINPUT74), .A3(new_n547), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n580), .A2(new_n556), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n556), .A3(new_n582), .ZN(new_n586));
  AOI22_X1  g400(.A1(KEYINPUT31), .A2(new_n586), .B1(new_n542), .B2(new_n548), .ZN(new_n587));
  AOI211_X1 g401(.A(KEYINPUT32), .B(new_n569), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n589), .B1(new_n592), .B2(new_n568), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n567), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n313), .A2(G119), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n457), .A2(G128), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT24), .B(G110), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n313), .A2(KEYINPUT79), .A3(G119), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT79), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT78), .B1(new_n596), .B2(KEYINPUT23), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT23), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n595), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n599), .B1(new_n607), .B2(G110), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n262), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n597), .A2(new_n598), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n607), .B2(G110), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n240), .A3(new_n201), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT22), .B(G137), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n204), .A2(G221), .A3(G234), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n609), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n609), .B2(new_n612), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(KEYINPUT25), .A3(new_n292), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n612), .ZN(new_n620));
  INV_X1    g434(.A(new_n615), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n609), .A2(new_n612), .A3(new_n615), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n292), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT25), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n326), .B1(new_n292), .B2(G234), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(G902), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n627), .A2(new_n628), .B1(new_n629), .B2(new_n618), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n514), .A2(new_n594), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  AOI22_X1  g446(.A1(new_n269), .A2(KEYINPUT92), .B1(new_n273), .B2(new_n275), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n283), .B1(new_n633), .B2(new_n272), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n511), .A2(new_n295), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n324), .A2(KEYINPUT97), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n331), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n329), .A2(new_n636), .A3(KEYINPUT33), .A4(new_n330), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(G478), .A3(new_n292), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n331), .A2(new_n292), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n296), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n634), .A2(new_n635), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n569), .B1(new_n585), .B2(new_n587), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n592), .A2(new_n292), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(G472), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n438), .A2(new_n630), .A3(new_n512), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NAND3_X1  g466(.A1(new_n266), .A2(new_n268), .A3(new_n274), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n283), .B1(new_n276), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n335), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n635), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n648), .A3(new_n649), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n592), .B2(new_n292), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n513), .A2(new_n662), .A3(new_n646), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n627), .A2(new_n628), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n620), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n629), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n336), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NOR2_X1   g486(.A1(new_n513), .A2(new_n668), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n288), .B1(new_n293), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n656), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n594), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n675), .B(KEYINPUT39), .Z(new_n679));
  NAND3_X1  g493(.A1(new_n438), .A2(new_n512), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n509), .A2(new_n510), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n668), .A2(new_n439), .A3(new_n655), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n681), .A2(new_n634), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n548), .B1(new_n560), .B2(new_n561), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n586), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n688), .B2(G902), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n588), .B2(new_n593), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n686), .B(new_n690), .C1(KEYINPUT40), .C2(new_n680), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n215), .ZN(G45));
  AOI211_X1 g506(.A(new_n644), .B(new_n675), .C1(new_n277), .C2(new_n284), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n594), .A2(new_n693), .A3(new_n673), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  INV_X1    g509(.A(new_n630), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n592), .A2(new_n568), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT32), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n646), .A2(new_n589), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n696), .B1(new_n700), .B2(new_n567), .ZN(new_n701));
  INV_X1    g515(.A(new_n420), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n419), .B1(new_n373), .B2(new_n400), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n340), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n430), .A2(new_n420), .A3(new_n341), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n333), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n432), .B(new_n512), .C1(new_n706), .C2(new_n437), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n701), .A2(KEYINPUT99), .A3(new_n645), .A4(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n645), .A2(new_n594), .A3(new_n630), .A4(new_n708), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT99), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n594), .A2(new_n630), .A3(new_n657), .A4(new_n708), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  INV_X1    g531(.A(KEYINPUT100), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n708), .A2(new_n718), .A3(new_n511), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n682), .A2(new_n439), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT100), .B1(new_n720), .B2(new_n707), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n594), .A3(new_n669), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  XNOR2_X1  g538(.A(new_n568), .B(KEYINPUT101), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n564), .A2(new_n548), .B1(KEYINPUT31), .B2(new_n586), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(new_n726), .B2(new_n585), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n662), .A2(new_n696), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n277), .A2(new_n284), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n720), .A2(new_n707), .A3(new_n294), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n655), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NOR3_X1   g546(.A1(new_n662), .A2(new_n668), .A3(new_n727), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n722), .A2(new_n693), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  AND3_X1   g549(.A1(new_n495), .A2(new_n505), .A3(new_n507), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n507), .B1(new_n495), .B2(new_n505), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n736), .A2(new_n737), .A3(new_n440), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n438), .A2(new_n738), .A3(new_n512), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n438), .A2(new_n738), .A3(KEYINPUT102), .A4(new_n512), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n693), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n698), .A2(new_n744), .A3(new_n699), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT103), .B1(new_n588), .B2(new_n593), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n567), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n743), .A2(new_n747), .A3(KEYINPUT42), .A4(new_n630), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n594), .A2(new_n630), .A3(new_n741), .A4(new_n742), .ZN(new_n750));
  INV_X1    g564(.A(new_n693), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n748), .A2(new_n752), .A3(KEYINPUT104), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT104), .B1(new_n748), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  INV_X1    g570(.A(new_n676), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n750), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n312), .ZN(G36));
  NAND2_X1  g573(.A1(new_n434), .A2(new_n435), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n437), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT46), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n432), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n512), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n679), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT105), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n664), .A2(new_n667), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n729), .A2(new_n644), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT43), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  OAI221_X1 g590(.A(new_n773), .B1(new_n646), .B2(new_n662), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n772), .A2(new_n780), .A3(new_n738), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  XNOR2_X1  g597(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n770), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n693), .A2(new_n696), .A3(new_n738), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n785), .A2(new_n594), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT108), .B(G140), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G42));
  AND2_X1   g603(.A1(new_n775), .A2(new_n288), .ZN(new_n790));
  INV_X1    g604(.A(new_n738), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n707), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n747), .A2(new_n630), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT48), .Z(new_n796));
  INV_X1    g610(.A(new_n690), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n630), .A2(new_n797), .A3(new_n288), .A4(new_n792), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n644), .B1(new_n277), .B2(new_n284), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n285), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n790), .A2(new_n728), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n722), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT117), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n796), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT118), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n706), .A2(new_n437), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n807), .A2(new_n766), .A3(new_n512), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n791), .B1(new_n785), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n707), .A2(new_n439), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT114), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n684), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT115), .Z(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n802), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n802), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT50), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n798), .A2(new_n634), .A3(new_n644), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT116), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n793), .A2(new_n733), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n816), .A2(new_n818), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT51), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n733), .A2(new_n693), .A3(new_n741), .A4(new_n742), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n750), .B2(new_n757), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n631), .A2(new_n670), .ZN(new_n828));
  INV_X1    g642(.A(new_n635), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n648), .A2(new_n649), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT109), .B1(new_n634), .B2(new_n644), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT109), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n641), .A2(new_n300), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n331), .A2(new_n292), .A3(new_n301), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n332), .B2(new_n334), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n799), .A2(new_n832), .B1(new_n634), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n830), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n828), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n838), .A2(new_n675), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n773), .A2(new_n842), .A3(new_n654), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n739), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT111), .B1(new_n844), .B2(new_n594), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n594), .A3(KEYINPUT111), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n827), .A2(new_n841), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT113), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n634), .A2(new_n720), .A3(new_n335), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n438), .A2(new_n512), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n773), .A3(new_n675), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n690), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n734), .A2(new_n677), .A3(new_n694), .A4(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n734), .A2(new_n677), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n858), .A2(new_n856), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n748), .A2(new_n752), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n723), .A2(new_n716), .A3(new_n731), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n712), .B2(new_n709), .ZN(new_n862));
  AND4_X1   g676(.A1(KEYINPUT53), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n850), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n799), .A2(new_n832), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n634), .A2(new_n838), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n831), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n830), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n631), .A3(new_n670), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n844), .A2(new_n594), .A3(KEYINPUT111), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n845), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n871), .A2(new_n873), .A3(new_n826), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n860), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n748), .A2(new_n752), .A3(KEYINPUT104), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n874), .A2(new_n876), .A3(new_n877), .A4(new_n862), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n855), .B(KEYINPUT52), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT112), .B(new_n865), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n723), .A2(new_n716), .A3(new_n731), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n713), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n849), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n755), .A3(new_n857), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT112), .B1(new_n885), .B2(new_n865), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n824), .B(new_n864), .C1(new_n881), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n865), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n859), .A2(new_n865), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n806), .A2(new_n823), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n643), .A2(new_n512), .A3(new_n439), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n684), .A2(new_n630), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n807), .A2(new_n766), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT49), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n797), .A3(new_n898), .A4(new_n634), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G75));
  OAI21_X1  g714(.A(new_n864), .B1(new_n881), .B2(new_n886), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n333), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n508), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n499), .A2(new_n504), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n502), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n904), .B2(new_n905), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n204), .A2(G952), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n887), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n764), .B(KEYINPUT57), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n915), .A2(new_n916), .B1(new_n421), .B2(new_n431), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n902), .A2(new_n763), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n266), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n911), .ZN(G60));
  XOR2_X1   g738(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n925));
  NOR2_X1   g739(.A1(new_n296), .A2(new_n282), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n887), .B2(new_n891), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n638), .A2(new_n639), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT121), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n930), .A2(new_n928), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n914), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n934), .ZN(new_n936));
  AOI211_X1 g750(.A(KEYINPUT120), .B(new_n936), .C1(new_n913), .C2(new_n887), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n932), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n911), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n930), .B1(new_n892), .B2(new_n928), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(KEYINPUT121), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT60), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n901), .A2(new_n666), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n901), .A2(new_n944), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n939), .B(new_n945), .C1(new_n946), .C2(new_n618), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n947), .A2(KEYINPUT122), .A3(new_n949), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  NOR2_X1   g767(.A1(new_n883), .A2(new_n871), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(G953), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT124), .Z(new_n956));
  AOI21_X1  g770(.A(new_n204), .B1(new_n290), .B2(G224), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n906), .B1(G898), .B2(new_n204), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G69));
  OAI211_X1 g775(.A(new_n858), .B(new_n694), .C1(new_n757), .C2(new_n750), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n794), .A2(new_n851), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n772), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n755), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n966), .A2(new_n782), .A3(new_n967), .A4(new_n787), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n782), .A2(new_n787), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT126), .B1(new_n969), .B2(new_n965), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n204), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n570), .A2(new_n571), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n232), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(G900), .B2(G953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n691), .A2(new_n694), .A3(new_n858), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT62), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n680), .A2(new_n791), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n868), .A2(new_n701), .A3(new_n978), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n969), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n973), .B1(new_n980), .B2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n204), .B1(G227), .B2(G900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n975), .A2(new_n985), .A3(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  INV_X1    g803(.A(new_n586), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n890), .B(new_n989), .C1(new_n990), .C2(new_n557), .ZN(new_n991));
  INV_X1    g805(.A(new_n989), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n980), .B2(new_n954), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n556), .A2(new_n529), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n547), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n939), .B(new_n991), .C1(new_n993), .C2(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n968), .A2(new_n954), .A3(new_n970), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(KEYINPUT127), .A3(new_n989), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n994), .A2(new_n547), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n989), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n996), .B1(new_n1000), .B2(new_n1003), .ZN(G57));
endmodule


