

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775;

  NAND2_X1 U374 ( .A1(n693), .A2(n692), .ZN(n616) );
  OR2_X1 U375 ( .A1(n405), .A2(n438), .ZN(n402) );
  NOR2_X1 U376 ( .A1(n664), .A2(n665), .ZN(n626) );
  NAND2_X1 U377 ( .A1(n555), .A2(n653), .ZN(n541) );
  AND2_X2 U378 ( .A1(n404), .A2(n435), .ZN(n403) );
  XNOR2_X2 U379 ( .A(n409), .B(n534), .ZN(n555) );
  INV_X2 U380 ( .A(G143), .ZN(n425) );
  XNOR2_X2 U381 ( .A(n610), .B(KEYINPUT33), .ZN(n685) );
  NOR2_X2 U382 ( .A1(n722), .A2(n545), .ZN(n546) );
  XNOR2_X2 U383 ( .A(n493), .B(n454), .ZN(n426) );
  AND2_X1 U384 ( .A1(n399), .A2(n398), .ZN(n397) );
  XNOR2_X1 U385 ( .A(n628), .B(n495), .ZN(n635) );
  XNOR2_X1 U386 ( .A(n737), .B(n736), .ZN(n738) );
  XNOR2_X1 U387 ( .A(n386), .B(n466), .ZN(n747) );
  XNOR2_X1 U388 ( .A(n741), .B(KEYINPUT122), .ZN(n742) );
  XNOR2_X1 U389 ( .A(G137), .B(G134), .ZN(n449) );
  INV_X1 U390 ( .A(n671), .ZN(n628) );
  XNOR2_X1 U391 ( .A(n458), .B(G125), .ZN(n524) );
  INV_X1 U392 ( .A(G146), .ZN(n458) );
  NAND2_X2 U393 ( .A1(n392), .A2(n389), .ZN(n551) );
  OR2_X1 U394 ( .A1(n426), .A2(n390), .ZN(n389) );
  AND2_X1 U395 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U396 ( .A1(n457), .A2(n391), .ZN(n390) );
  AND2_X1 U397 ( .A1(n419), .A2(n418), .ZN(n383) );
  NAND2_X1 U398 ( .A1(n403), .A2(n402), .ZN(n693) );
  XNOR2_X1 U399 ( .A(KEYINPUT87), .B(KEYINPUT48), .ZN(n577) );
  INV_X1 U400 ( .A(G237), .ZN(n531) );
  AND2_X1 U401 ( .A1(G953), .A2(G902), .ZN(n474) );
  XNOR2_X1 U402 ( .A(n488), .B(G113), .ZN(n489) );
  NOR2_X1 U403 ( .A1(G953), .A2(G237), .ZN(n500) );
  XNOR2_X1 U404 ( .A(n451), .B(n408), .ZN(n407) );
  INV_X1 U405 ( .A(G107), .ZN(n408) );
  XNOR2_X1 U406 ( .A(n406), .B(G140), .ZN(n497) );
  INV_X1 U407 ( .A(G131), .ZN(n406) );
  XNOR2_X1 U408 ( .A(KEYINPUT4), .B(KEYINPUT67), .ZN(n448) );
  XNOR2_X1 U409 ( .A(n521), .B(n524), .ZN(n433) );
  XOR2_X1 U410 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n521) );
  INV_X1 U411 ( .A(n628), .ZN(n437) );
  XNOR2_X1 U412 ( .A(KEYINPUT16), .B(G110), .ZN(n525) );
  XNOR2_X1 U413 ( .A(G140), .B(KEYINPUT24), .ZN(n460) );
  XNOR2_X1 U414 ( .A(n354), .B(n524), .ZN(n496) );
  XOR2_X1 U415 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n464) );
  NOR2_X1 U416 ( .A1(n725), .A2(n428), .ZN(n427) );
  OR2_X1 U417 ( .A1(n635), .A2(n429), .ZN(n428) );
  BUF_X1 U418 ( .A(n555), .Z(n584) );
  XNOR2_X1 U419 ( .A(n378), .B(KEYINPUT74), .ZN(n570) );
  NOR2_X1 U420 ( .A1(n415), .A2(n553), .ZN(n414) );
  NAND2_X1 U421 ( .A1(n437), .A2(KEYINPUT64), .ZN(n436) );
  XNOR2_X1 U422 ( .A(n470), .B(n469), .ZN(n471) );
  INV_X1 U423 ( .A(KEYINPUT44), .ZN(n412) );
  INV_X1 U424 ( .A(n569), .ZN(n654) );
  NAND2_X1 U425 ( .A1(n395), .A2(G902), .ZN(n393) );
  XOR2_X1 U426 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n499) );
  XNOR2_X1 U427 ( .A(G113), .B(G104), .ZN(n527) );
  XNOR2_X1 U428 ( .A(G902), .B(KEYINPUT15), .ZN(n697) );
  NAND2_X1 U429 ( .A1(n400), .A2(n397), .ZN(n396) );
  INV_X1 U430 ( .A(KEYINPUT86), .ZN(n384) );
  INV_X1 U431 ( .A(n733), .ZN(n440) );
  NAND2_X1 U432 ( .A1(G234), .A2(G237), .ZN(n473) );
  XNOR2_X1 U433 ( .A(n584), .B(KEYINPUT38), .ZN(n569) );
  XNOR2_X1 U434 ( .A(n444), .B(KEYINPUT30), .ZN(n415) );
  XNOR2_X1 U435 ( .A(n529), .B(n489), .ZN(n491) );
  XOR2_X1 U436 ( .A(G104), .B(G110), .Z(n452) );
  XNOR2_X1 U437 ( .A(n407), .B(n497), .ZN(n453) );
  XNOR2_X1 U438 ( .A(n522), .B(n523), .ZN(n431) );
  XOR2_X1 U439 ( .A(KEYINPUT41), .B(n565), .Z(n684) );
  NOR2_X1 U440 ( .A1(n658), .A2(n657), .ZN(n565) );
  XNOR2_X1 U441 ( .A(n496), .B(n465), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n536), .B(KEYINPUT36), .ZN(n423) );
  XNOR2_X1 U443 ( .A(n606), .B(n605), .ZN(n692) );
  OR2_X1 U444 ( .A1(n613), .A2(n556), .ZN(n557) );
  AND2_X1 U445 ( .A1(n436), .A2(n599), .ZN(n435) );
  XNOR2_X1 U446 ( .A(n573), .B(KEYINPUT105), .ZN(n725) );
  AND2_X1 U447 ( .A1(n411), .A2(n623), .ZN(n624) );
  XOR2_X1 U448 ( .A(n356), .B(n459), .Z(n353) );
  XOR2_X1 U449 ( .A(KEYINPUT10), .B(KEYINPUT68), .Z(n354) );
  AND2_X1 U450 ( .A1(n380), .A2(n519), .ZN(n355) );
  XOR2_X1 U451 ( .A(G110), .B(G128), .Z(n356) );
  INV_X1 U452 ( .A(n457), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U454 ( .A(G902), .ZN(n391) );
  XOR2_X1 U455 ( .A(KEYINPUT85), .B(KEYINPUT35), .Z(n357) );
  XOR2_X1 U456 ( .A(n709), .B(n708), .Z(n358) );
  XOR2_X1 U457 ( .A(n706), .B(KEYINPUT59), .Z(n359) );
  XOR2_X1 U458 ( .A(n703), .B(n702), .Z(n360) );
  NOR2_X1 U459 ( .A1(n607), .A2(KEYINPUT44), .ZN(n361) );
  XNOR2_X1 U460 ( .A(KEYINPUT119), .B(KEYINPUT56), .ZN(n362) );
  XNOR2_X1 U461 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n363) );
  XOR2_X1 U462 ( .A(n711), .B(KEYINPUT90), .Z(n364) );
  OR2_X1 U463 ( .A1(n697), .A2(n696), .ZN(n365) );
  AND2_X1 U464 ( .A1(n705), .A2(G953), .ZN(n749) );
  INV_X1 U465 ( .A(n749), .ZN(n375) );
  INV_X2 U466 ( .A(G953), .ZN(n519) );
  INV_X1 U467 ( .A(n645), .ZN(n366) );
  XNOR2_X1 U468 ( .A(n396), .B(n644), .ZN(n750) );
  INV_X1 U469 ( .A(n584), .ZN(n556) );
  NOR2_X1 U470 ( .A1(n367), .A2(n616), .ZN(n617) );
  NOR2_X1 U471 ( .A1(n388), .A2(n640), .ZN(n367) );
  NOR2_X1 U472 ( .A1(n641), .A2(n412), .ZN(n639) );
  NAND2_X1 U473 ( .A1(n638), .A2(n712), .ZN(n641) );
  BUF_X1 U474 ( .A(n541), .Z(n368) );
  XNOR2_X1 U475 ( .A(n368), .B(KEYINPUT19), .ZN(n369) );
  XNOR2_X1 U476 ( .A(n541), .B(KEYINPUT19), .ZN(n590) );
  NAND2_X1 U477 ( .A1(n403), .A2(n402), .ZN(n370) );
  XNOR2_X1 U478 ( .A(n629), .B(KEYINPUT94), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n493), .B(n492), .ZN(n709) );
  BUF_X1 U480 ( .A(n611), .Z(n629) );
  XNOR2_X1 U481 ( .A(n434), .B(n591), .ZN(n611) );
  NAND2_X1 U482 ( .A1(n611), .A2(n594), .ZN(n597) );
  XNOR2_X1 U483 ( .A(n371), .B(n362), .ZN(G51) );
  NAND2_X1 U484 ( .A1(n377), .A2(n375), .ZN(n371) );
  XNOR2_X1 U485 ( .A(n372), .B(n363), .ZN(G60) );
  NAND2_X1 U486 ( .A1(n374), .A2(n375), .ZN(n372) );
  XNOR2_X1 U487 ( .A(n373), .B(n364), .ZN(G57) );
  NAND2_X1 U488 ( .A1(n376), .A2(n375), .ZN(n373) );
  XNOR2_X1 U489 ( .A(n707), .B(n359), .ZN(n374) );
  XNOR2_X1 U490 ( .A(n710), .B(n358), .ZN(n376) );
  XNOR2_X1 U491 ( .A(n704), .B(n360), .ZN(n377) );
  XNOR2_X1 U492 ( .A(n695), .B(KEYINPUT83), .ZN(n381) );
  NAND2_X1 U493 ( .A1(n414), .A2(n623), .ZN(n378) );
  INV_X1 U494 ( .A(n762), .ZN(n382) );
  NAND2_X1 U495 ( .A1(n379), .A2(n365), .ZN(n699) );
  NAND2_X1 U496 ( .A1(n381), .A2(n382), .ZN(n379) );
  XNOR2_X1 U497 ( .A(n691), .B(KEYINPUT118), .ZN(n380) );
  XNOR2_X1 U498 ( .A(n624), .B(KEYINPUT98), .ZN(n625) );
  NAND2_X1 U499 ( .A1(n383), .A2(n420), .ZN(n424) );
  XNOR2_X1 U500 ( .A(n421), .B(KEYINPUT69), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n385), .B(n384), .ZN(n649) );
  NAND2_X1 U502 ( .A1(n441), .A2(n440), .ZN(n385) );
  NAND2_X1 U503 ( .A1(n388), .A2(n361), .ZN(n620) );
  OR2_X2 U504 ( .A1(n388), .A2(KEYINPUT66), .ZN(n619) );
  NAND2_X1 U505 ( .A1(n639), .A2(n387), .ZN(n643) );
  INV_X1 U506 ( .A(n388), .ZN(n387) );
  XNOR2_X1 U507 ( .A(n388), .B(G122), .ZN(n773) );
  XNOR2_X2 U508 ( .A(n615), .B(n357), .ZN(n388) );
  NAND2_X1 U509 ( .A1(n426), .A2(n395), .ZN(n394) );
  XNOR2_X2 U510 ( .A(n551), .B(KEYINPUT1), .ZN(n664) );
  NAND2_X1 U511 ( .A1(n643), .A2(n642), .ZN(n398) );
  NAND2_X1 U512 ( .A1(n622), .A2(n621), .ZN(n399) );
  NAND2_X1 U513 ( .A1(n401), .A2(KEYINPUT44), .ZN(n400) );
  NAND2_X1 U514 ( .A1(n618), .A2(n617), .ZN(n401) );
  XNOR2_X2 U515 ( .A(n761), .B(n450), .ZN(n493) );
  XNOR2_X2 U516 ( .A(n413), .B(n449), .ZN(n761) );
  XNOR2_X2 U517 ( .A(n511), .B(n448), .ZN(n413) );
  NAND2_X1 U518 ( .A1(n405), .A2(KEYINPUT64), .ZN(n404) );
  XNOR2_X2 U519 ( .A(n637), .B(KEYINPUT103), .ZN(n405) );
  OR2_X2 U520 ( .A1(n700), .A2(n694), .ZN(n409) );
  XNOR2_X1 U521 ( .A(n410), .B(n755), .ZN(n700) );
  XNOR2_X1 U522 ( .A(n432), .B(n431), .ZN(n410) );
  NAND2_X1 U523 ( .A1(n685), .A2(n411), .ZN(n612) );
  XNOR2_X1 U524 ( .A(n413), .B(n433), .ZN(n432) );
  NAND2_X1 U525 ( .A1(n417), .A2(n416), .ZN(n420) );
  NOR2_X1 U526 ( .A1(n560), .A2(KEYINPUT73), .ZN(n416) );
  INV_X1 U527 ( .A(n561), .ZN(n417) );
  NAND2_X1 U528 ( .A1(n560), .A2(KEYINPUT73), .ZN(n418) );
  NAND2_X1 U529 ( .A1(n561), .A2(KEYINPUT73), .ZN(n419) );
  INV_X1 U530 ( .A(n422), .ZN(n730) );
  NAND2_X1 U531 ( .A1(n424), .A2(n422), .ZN(n421) );
  NAND2_X1 U532 ( .A1(n423), .A2(n581), .ZN(n422) );
  XNOR2_X2 U533 ( .A(n425), .B(G128), .ZN(n511) );
  XNOR2_X1 U534 ( .A(n426), .B(KEYINPUT120), .ZN(n736) );
  XNOR2_X1 U535 ( .A(n427), .B(KEYINPUT107), .ZN(n578) );
  INV_X1 U536 ( .A(n537), .ZN(n429) );
  XNOR2_X1 U537 ( .A(n430), .B(n760), .ZN(n706) );
  XNOR2_X1 U538 ( .A(n496), .B(n497), .ZN(n760) );
  XNOR2_X1 U539 ( .A(n502), .B(n504), .ZN(n430) );
  NAND2_X1 U540 ( .A1(n590), .A2(n446), .ZN(n434) );
  NAND2_X1 U541 ( .A1(n628), .A2(n598), .ZN(n438) );
  NAND2_X1 U542 ( .A1(n439), .A2(n559), .ZN(n560) );
  XNOR2_X1 U543 ( .A(n439), .B(G143), .ZN(G45) );
  XNOR2_X1 U544 ( .A(n558), .B(KEYINPUT109), .ZN(n439) );
  XNOR2_X1 U545 ( .A(n442), .B(n577), .ZN(n441) );
  NAND2_X1 U546 ( .A1(n443), .A2(n576), .ZN(n442) );
  NAND2_X1 U547 ( .A1(n671), .A2(n653), .ZN(n444) );
  XNOR2_X2 U548 ( .A(n494), .B(G472), .ZN(n671) );
  AND2_X2 U549 ( .A1(n601), .A2(n664), .ZN(n637) );
  BUF_X1 U550 ( .A(n700), .Z(n703) );
  AND2_X1 U551 ( .A1(G214), .A2(n500), .ZN(n445) );
  OR2_X1 U552 ( .A1(n589), .A2(n588), .ZN(n446) );
  INV_X1 U553 ( .A(KEYINPUT66), .ZN(n607) );
  XNOR2_X1 U554 ( .A(n501), .B(n445), .ZN(n502) );
  INV_X1 U555 ( .A(G469), .ZN(n455) );
  XNOR2_X1 U556 ( .A(n743), .B(n742), .ZN(n744) );
  INV_X1 U557 ( .A(KEYINPUT65), .ZN(n447) );
  XNOR2_X1 U558 ( .A(n447), .B(G101), .ZN(n523) );
  XNOR2_X1 U559 ( .A(n523), .B(G146), .ZN(n450) );
  NAND2_X1 U560 ( .A1(G227), .A2(n519), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U562 ( .A(KEYINPUT70), .ZN(n456) );
  XNOR2_X1 U563 ( .A(G119), .B(G137), .ZN(n459) );
  XOR2_X1 U564 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n461) );
  XNOR2_X1 U565 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n353), .B(n462), .ZN(n466) );
  NAND2_X1 U567 ( .A1(G234), .A2(n519), .ZN(n463) );
  XNOR2_X1 U568 ( .A(n464), .B(n463), .ZN(n514) );
  NAND2_X1 U569 ( .A1(G221), .A2(n514), .ZN(n465) );
  NOR2_X1 U570 ( .A1(G902), .A2(n747), .ZN(n472) );
  NAND2_X1 U571 ( .A1(n697), .A2(G234), .ZN(n467) );
  XNOR2_X1 U572 ( .A(n467), .B(KEYINPUT20), .ZN(n481) );
  AND2_X1 U573 ( .A1(n481), .A2(G217), .ZN(n468) );
  XNOR2_X1 U574 ( .A(n468), .B(KEYINPUT25), .ZN(n470) );
  XNOR2_X1 U575 ( .A(KEYINPUT75), .B(KEYINPUT96), .ZN(n469) );
  XNOR2_X2 U576 ( .A(n472), .B(n471), .ZN(n667) );
  XNOR2_X1 U577 ( .A(n473), .B(KEYINPUT14), .ZN(n476) );
  NAND2_X1 U578 ( .A1(n476), .A2(n474), .ZN(n587) );
  XNOR2_X1 U579 ( .A(KEYINPUT106), .B(n587), .ZN(n475) );
  NOR2_X1 U580 ( .A1(G900), .A2(n475), .ZN(n479) );
  NAND2_X1 U581 ( .A1(G952), .A2(n476), .ZN(n683) );
  NOR2_X1 U582 ( .A1(G953), .A2(n683), .ZN(n478) );
  INV_X1 U583 ( .A(KEYINPUT93), .ZN(n477) );
  XNOR2_X1 U584 ( .A(n478), .B(n477), .ZN(n589) );
  NOR2_X1 U585 ( .A1(n479), .A2(n589), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n480), .B(KEYINPUT79), .ZN(n552) );
  NAND2_X1 U587 ( .A1(n481), .A2(G221), .ZN(n483) );
  INV_X1 U588 ( .A(KEYINPUT21), .ZN(n482) );
  XNOR2_X1 U589 ( .A(n483), .B(n482), .ZN(n668) );
  NAND2_X1 U590 ( .A1(n552), .A2(n668), .ZN(n484) );
  NOR2_X1 U591 ( .A1(n667), .A2(n484), .ZN(n537) );
  INV_X1 U592 ( .A(KEYINPUT71), .ZN(n485) );
  XNOR2_X1 U593 ( .A(n485), .B(KEYINPUT3), .ZN(n487) );
  XNOR2_X1 U594 ( .A(G119), .B(G116), .ZN(n486) );
  XNOR2_X1 U595 ( .A(n487), .B(n486), .ZN(n529) );
  XOR2_X1 U596 ( .A(KEYINPUT5), .B(G131), .Z(n488) );
  NAND2_X1 U597 ( .A1(G210), .A2(n500), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U599 ( .A1(n709), .A2(n391), .ZN(n494) );
  INV_X1 U600 ( .A(KEYINPUT6), .ZN(n495) );
  XNOR2_X1 U601 ( .A(G143), .B(G122), .ZN(n498) );
  XNOR2_X1 U602 ( .A(n499), .B(n498), .ZN(n501) );
  INV_X1 U603 ( .A(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n527), .B(n503), .ZN(n504) );
  NAND2_X1 U605 ( .A1(n706), .A2(n391), .ZN(n506) );
  XNOR2_X1 U606 ( .A(KEYINPUT13), .B(G475), .ZN(n505) );
  XNOR2_X1 U607 ( .A(n506), .B(n505), .ZN(n564) );
  XOR2_X1 U608 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n508) );
  XNOR2_X1 U609 ( .A(G116), .B(G134), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n508), .B(n507), .ZN(n513) );
  XOR2_X1 U611 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n509) );
  XNOR2_X2 U612 ( .A(G122), .B(G107), .ZN(n526) );
  XOR2_X1 U613 ( .A(n509), .B(n526), .Z(n510) );
  XNOR2_X1 U614 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U615 ( .A(n513), .B(n512), .Z(n516) );
  NAND2_X1 U616 ( .A1(n514), .A2(G217), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n516), .B(n515), .ZN(n741) );
  NOR2_X1 U618 ( .A1(n741), .A2(G902), .ZN(n518) );
  INV_X1 U619 ( .A(G478), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n518), .B(n517), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n564), .A2(n562), .ZN(n573) );
  NAND2_X1 U622 ( .A1(n519), .A2(G224), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n520), .B(KEYINPUT76), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n526), .B(n525), .ZN(n528) );
  XNOR2_X1 U625 ( .A(n528), .B(n527), .ZN(n530) );
  XNOR2_X1 U626 ( .A(n530), .B(n529), .ZN(n755) );
  INV_X1 U627 ( .A(n697), .ZN(n694) );
  NAND2_X1 U628 ( .A1(n391), .A2(n531), .ZN(n535) );
  NAND2_X1 U629 ( .A1(n535), .A2(G210), .ZN(n533) );
  INV_X1 U630 ( .A(KEYINPUT92), .ZN(n532) );
  XNOR2_X1 U631 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U632 ( .A1(n535), .A2(G214), .ZN(n653) );
  NOR2_X1 U633 ( .A1(n578), .A2(n368), .ZN(n536) );
  AND2_X1 U634 ( .A1(n671), .A2(n537), .ZN(n538) );
  XNOR2_X1 U635 ( .A(n538), .B(KEYINPUT28), .ZN(n540) );
  INV_X1 U636 ( .A(n551), .ZN(n539) );
  NAND2_X1 U637 ( .A1(n540), .A2(n539), .ZN(n567) );
  INV_X1 U638 ( .A(n567), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n542), .A2(n369), .ZN(n544) );
  INV_X1 U640 ( .A(KEYINPUT78), .ZN(n543) );
  XNOR2_X2 U641 ( .A(n544), .B(n543), .ZN(n722) );
  INV_X1 U642 ( .A(KEYINPUT47), .ZN(n545) );
  XNOR2_X1 U643 ( .A(n546), .B(KEYINPUT81), .ZN(n549) );
  AND2_X1 U644 ( .A1(n564), .A2(n562), .ZN(n718) );
  NOR2_X1 U645 ( .A1(n573), .A2(n718), .ZN(n659) );
  NOR2_X1 U646 ( .A1(KEYINPUT47), .A2(n659), .ZN(n547) );
  NAND2_X1 U647 ( .A1(n722), .A2(n547), .ZN(n548) );
  NAND2_X1 U648 ( .A1(n549), .A2(n548), .ZN(n561) );
  INV_X1 U649 ( .A(KEYINPUT97), .ZN(n550) );
  XNOR2_X1 U650 ( .A(n668), .B(n550), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n667), .A2(n592), .ZN(n665) );
  NOR2_X1 U652 ( .A1(n551), .A2(n665), .ZN(n623) );
  INV_X1 U653 ( .A(n552), .ZN(n553) );
  INV_X1 U654 ( .A(n564), .ZN(n554) );
  NAND2_X1 U655 ( .A1(n554), .A2(n562), .ZN(n613) );
  NOR2_X1 U656 ( .A1(n570), .A2(n557), .ZN(n558) );
  NAND2_X1 U657 ( .A1(KEYINPUT47), .A2(n659), .ZN(n559) );
  NAND2_X1 U658 ( .A1(n654), .A2(n653), .ZN(n658) );
  INV_X1 U659 ( .A(n562), .ZN(n563) );
  AND2_X1 U660 ( .A1(n564), .A2(n563), .ZN(n593) );
  INV_X1 U661 ( .A(n593), .ZN(n657) );
  INV_X1 U662 ( .A(n684), .ZN(n566) );
  NOR2_X1 U663 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U664 ( .A(n568), .B(KEYINPUT42), .ZN(n775) );
  NOR2_X1 U665 ( .A1(n570), .A2(n569), .ZN(n572) );
  INV_X1 U666 ( .A(KEYINPUT39), .ZN(n571) );
  XNOR2_X1 U667 ( .A(n572), .B(n571), .ZN(n586) );
  AND2_X1 U668 ( .A1(n573), .A2(n586), .ZN(n574) );
  XNOR2_X1 U669 ( .A(n574), .B(KEYINPUT40), .ZN(n774) );
  NOR2_X1 U670 ( .A1(n775), .A2(n774), .ZN(n575) );
  XNOR2_X1 U671 ( .A(KEYINPUT46), .B(n575), .ZN(n576) );
  INV_X1 U672 ( .A(n664), .ZN(n581) );
  INV_X1 U673 ( .A(n578), .ZN(n579) );
  NAND2_X1 U674 ( .A1(n579), .A2(n653), .ZN(n580) );
  NOR2_X1 U675 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U676 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n582) );
  XNOR2_X1 U677 ( .A(n583), .B(n582), .ZN(n585) );
  NOR2_X1 U678 ( .A1(n585), .A2(n584), .ZN(n733) );
  NAND2_X1 U679 ( .A1(n586), .A2(n718), .ZN(n732) );
  NAND2_X1 U680 ( .A1(n649), .A2(n732), .ZN(n762) );
  NOR2_X1 U681 ( .A1(n587), .A2(G898), .ZN(n588) );
  INV_X1 U682 ( .A(KEYINPUT0), .ZN(n591) );
  AND2_X1 U683 ( .A1(n593), .A2(n592), .ZN(n594) );
  INV_X1 U684 ( .A(KEYINPUT72), .ZN(n595) );
  XNOR2_X1 U685 ( .A(n595), .B(KEYINPUT22), .ZN(n596) );
  XNOR2_X2 U686 ( .A(n597), .B(n596), .ZN(n601) );
  INV_X1 U687 ( .A(KEYINPUT64), .ZN(n598) );
  INV_X1 U688 ( .A(n667), .ZN(n599) );
  NOR2_X1 U689 ( .A1(n664), .A2(n667), .ZN(n600) );
  NAND2_X1 U690 ( .A1(n600), .A2(n635), .ZN(n603) );
  INV_X1 U691 ( .A(n601), .ZN(n602) );
  OR2_X1 U692 ( .A1(n603), .A2(n602), .ZN(n606) );
  INV_X1 U693 ( .A(KEYINPUT77), .ZN(n604) );
  XNOR2_X1 U694 ( .A(n604), .B(KEYINPUT32), .ZN(n605) );
  XNOR2_X2 U695 ( .A(n616), .B(KEYINPUT89), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n621), .A2(n607), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n626), .B(KEYINPUT104), .ZN(n609) );
  INV_X1 U698 ( .A(n635), .ZN(n608) );
  NAND2_X1 U699 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U700 ( .A(n612), .B(KEYINPUT34), .ZN(n614) );
  NOR2_X2 U701 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U702 ( .A1(n619), .A2(n620), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n625), .A2(n628), .ZN(n714) );
  INV_X1 U704 ( .A(n626), .ZN(n627) );
  OR2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n674) );
  INV_X1 U706 ( .A(n674), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n629), .A2(n630), .ZN(n632) );
  XNOR2_X1 U708 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n632), .B(n631), .ZN(n727) );
  NAND2_X1 U710 ( .A1(n714), .A2(n727), .ZN(n634) );
  INV_X1 U711 ( .A(n659), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n638) );
  AND2_X1 U713 ( .A1(n635), .A2(n667), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n712) );
  INV_X1 U715 ( .A(KEYINPUT88), .ZN(n640) );
  OR2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U717 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n644) );
  INV_X1 U718 ( .A(n750), .ZN(n645) );
  NOR2_X1 U719 ( .A1(n762), .A2(n645), .ZN(n646) );
  NOR2_X1 U720 ( .A1(n646), .A2(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U721 ( .A1(KEYINPUT2), .A2(n732), .ZN(n647) );
  XOR2_X1 U722 ( .A(KEYINPUT80), .B(n647), .Z(n648) );
  AND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n650), .A2(n366), .ZN(n698) );
  INV_X1 U725 ( .A(n698), .ZN(n651) );
  NOR2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n690) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U728 ( .A(KEYINPUT115), .B(n655), .Z(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U732 ( .A(KEYINPUT116), .B(n662), .Z(n663) );
  NAND2_X1 U733 ( .A1(n663), .A2(n685), .ZN(n680) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n666), .B(KEYINPUT50), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U737 ( .A(KEYINPUT49), .B(n669), .Z(n670) );
  NOR2_X1 U738 ( .A1(n437), .A2(n670), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n677) );
  XOR2_X1 U741 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n676) );
  XNOR2_X1 U742 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n678), .A2(n684), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U745 ( .A(KEYINPUT52), .B(n681), .Z(n682) );
  NOR2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n687) );
  AND2_X1 U747 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT117), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n355), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U752 ( .A(n692), .B(G119), .ZN(G21) );
  XNOR2_X1 U753 ( .A(n370), .B(G110), .ZN(G12) );
  NAND2_X1 U754 ( .A1(n750), .A2(n694), .ZN(n695) );
  INV_X1 U755 ( .A(KEYINPUT2), .ZN(n696) );
  AND2_X2 U756 ( .A1(n699), .A2(n698), .ZN(n735) );
  NAND2_X1 U757 ( .A1(n735), .A2(G210), .ZN(n704) );
  XNOR2_X1 U758 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n701) );
  XNOR2_X1 U759 ( .A(n701), .B(KEYINPUT55), .ZN(n702) );
  INV_X1 U760 ( .A(G952), .ZN(n705) );
  NAND2_X1 U761 ( .A1(n735), .A2(G475), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n735), .A2(G472), .ZN(n710) );
  XOR2_X1 U763 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n708) );
  XNOR2_X1 U764 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n711) );
  XNOR2_X1 U765 ( .A(G101), .B(n712), .ZN(G3) );
  NOR2_X1 U766 ( .A1(n725), .A2(n714), .ZN(n713) );
  XOR2_X1 U767 ( .A(G104), .B(n713), .Z(G6) );
  INV_X1 U768 ( .A(n718), .ZN(n728) );
  NOR2_X1 U769 ( .A1(n728), .A2(n714), .ZN(n716) );
  XNOR2_X1 U770 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n715) );
  XNOR2_X1 U771 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U772 ( .A(G107), .B(n717), .ZN(G9) );
  XOR2_X1 U773 ( .A(G128), .B(KEYINPUT29), .Z(n720) );
  NAND2_X1 U774 ( .A1(n718), .A2(n722), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(G30) );
  INV_X1 U776 ( .A(n725), .ZN(n721) );
  NAND2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U778 ( .A(n723), .B(KEYINPUT112), .ZN(n724) );
  XNOR2_X1 U779 ( .A(G146), .B(n724), .ZN(G48) );
  NOR2_X1 U780 ( .A1(n725), .A2(n727), .ZN(n726) );
  XOR2_X1 U781 ( .A(G113), .B(n726), .Z(G15) );
  NOR2_X1 U782 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U783 ( .A(G116), .B(n729), .Z(G18) );
  XNOR2_X1 U784 ( .A(G125), .B(n730), .ZN(n731) );
  XNOR2_X1 U785 ( .A(n731), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U786 ( .A(G134), .B(n732), .ZN(G36) );
  XNOR2_X1 U787 ( .A(n733), .B(G140), .ZN(n734) );
  XNOR2_X1 U788 ( .A(n734), .B(KEYINPUT113), .ZN(G42) );
  BUF_X2 U789 ( .A(n735), .Z(n745) );
  NAND2_X1 U790 ( .A1(n745), .A2(G469), .ZN(n739) );
  XOR2_X1 U791 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n737) );
  XNOR2_X1 U792 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n749), .A2(n740), .ZN(G54) );
  NAND2_X1 U794 ( .A1(n745), .A2(G478), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n749), .A2(n744), .ZN(G63) );
  NAND2_X1 U796 ( .A1(n745), .A2(G217), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(n747), .ZN(n748) );
  NOR2_X1 U798 ( .A1(n749), .A2(n748), .ZN(G66) );
  NAND2_X1 U799 ( .A1(n366), .A2(n519), .ZN(n754) );
  NAND2_X1 U800 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U801 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U802 ( .A1(n752), .A2(G898), .ZN(n753) );
  NAND2_X1 U803 ( .A1(n754), .A2(n753), .ZN(n759) );
  XNOR2_X1 U804 ( .A(n755), .B(G101), .ZN(n757) );
  NOR2_X1 U805 ( .A1(n519), .A2(G898), .ZN(n756) );
  NOR2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n759), .B(n758), .ZN(G69) );
  XOR2_X1 U808 ( .A(n761), .B(n760), .Z(n766) );
  INV_X1 U809 ( .A(n766), .ZN(n763) );
  XOR2_X1 U810 ( .A(n763), .B(n762), .Z(n764) );
  NOR2_X1 U811 ( .A1(G953), .A2(n764), .ZN(n765) );
  XNOR2_X1 U812 ( .A(KEYINPUT123), .B(n765), .ZN(n772) );
  XOR2_X1 U813 ( .A(n766), .B(G227), .Z(n767) );
  XNOR2_X1 U814 ( .A(n767), .B(KEYINPUT124), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U816 ( .A1(G953), .A2(n769), .ZN(n770) );
  XOR2_X1 U817 ( .A(KEYINPUT125), .B(n770), .Z(n771) );
  NAND2_X1 U818 ( .A1(n772), .A2(n771), .ZN(G72) );
  XNOR2_X1 U819 ( .A(KEYINPUT126), .B(n773), .ZN(G24) );
  XOR2_X1 U820 ( .A(n774), .B(G131), .Z(G33) );
  XOR2_X1 U821 ( .A(G137), .B(n775), .Z(G39) );
endmodule

