//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G116), .B(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n195), .A2(new_n202), .A3(KEYINPUT66), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n193), .A2(new_n194), .A3(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT76), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT76), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G104), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n207), .A2(KEYINPUT3), .A3(G107), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G101), .ZN(new_n220));
  XOR2_X1   g034(.A(KEYINPUT77), .B(G101), .Z(new_n221));
  NAND4_X1  g035(.A1(new_n213), .A2(new_n215), .A3(new_n221), .A4(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n216), .B1(new_n212), .B2(KEYINPUT3), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n215), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n206), .B(new_n220), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n212), .A2(KEYINPUT78), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n207), .A2(G107), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT78), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n208), .A2(new_n210), .A3(new_n230), .A4(new_n211), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  OAI21_X1  g047(.A(G113), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n233), .A2(new_n202), .A3(new_n222), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n227), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(G110), .B(G122), .Z(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n227), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n241), .A2(KEYINPUT82), .A3(new_n243), .A4(KEYINPUT6), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n227), .A2(new_n238), .A3(new_n242), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n242), .B1(new_n227), .B2(new_n238), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n247), .A3(new_n240), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n244), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(KEYINPUT1), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n260), .A3(G143), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n256), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n258), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  OR2_X1    g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n266), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT65), .B1(new_n253), .B2(new_n269), .ZN(new_n270));
  AND4_X1   g084(.A1(KEYINPUT65), .A2(new_n269), .A3(new_n264), .A4(new_n258), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n263), .B1(G125), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G224), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n252), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT7), .B1(new_n274), .B2(G953), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n273), .B(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n240), .B(KEYINPUT8), .Z(new_n281));
  NAND2_X1  g095(.A1(new_n233), .A2(new_n222), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n202), .A3(new_n237), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n236), .B1(KEYINPUT83), .B2(new_n234), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(KEYINPUT83), .B2(new_n234), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n200), .B2(new_n201), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n281), .B(new_n283), .C1(new_n286), .C2(new_n282), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n280), .A2(new_n243), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n188), .B1(new_n278), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n243), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT82), .B1(new_n246), .B2(new_n247), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n276), .B1(new_n292), .B2(new_n244), .ZN(new_n293));
  INV_X1    g107(.A(new_n188), .ZN(new_n294));
  INV_X1    g108(.A(new_n288), .ZN(new_n295));
  NOR4_X1   g109(.A1(new_n293), .A2(G902), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n278), .A2(new_n188), .A3(new_n288), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT84), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT80), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT81), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT9), .B(G234), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT74), .ZN(new_n306));
  OAI21_X1  g120(.A(G221), .B1(new_n306), .B2(G902), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n307), .B(KEYINPUT75), .Z(new_n308));
  INV_X1    g122(.A(new_n262), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n282), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n233), .A2(new_n262), .A3(new_n222), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n313));
  INV_X1    g127(.A(G134), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G137), .ZN(new_n315));
  INV_X1    g129(.A(G137), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT11), .A3(G134), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(G137), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G131), .ZN(new_n320));
  INV_X1    g134(.A(G131), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n315), .A2(new_n317), .A3(new_n321), .A4(new_n318), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT12), .B1(new_n312), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n233), .A2(new_n262), .A3(new_n222), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n262), .B1(new_n233), .B2(new_n222), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT12), .B(new_n323), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT79), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n311), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n265), .B2(new_n266), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n253), .A2(KEYINPUT65), .A3(new_n269), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n253), .A2(new_n269), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n333), .A2(new_n334), .B1(new_n335), .B2(new_n267), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n336), .B(new_n220), .C1(new_n223), .C2(new_n226), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n320), .A2(new_n322), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n262), .A4(new_n222), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n331), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G140), .ZN(new_n342));
  INV_X1    g156(.A(G227), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G953), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n342), .B(new_n344), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT12), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n327), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n329), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n331), .A2(new_n337), .A3(new_n339), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n323), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n340), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n346), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G469), .ZN(new_n359));
  XOR2_X1   g173(.A(KEYINPUT70), .B(G902), .Z(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G902), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n340), .B1(new_n324), .B2(new_n328), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n365), .A2(new_n346), .B1(new_n347), .B2(new_n355), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n366), .B2(G469), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n308), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G475), .ZN(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT73), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n260), .ZN(new_n372));
  INV_X1    g186(.A(G140), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT71), .B1(new_n373), .B2(G125), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT71), .ZN(new_n375));
  INV_X1    g189(.A(G125), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G140), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n374), .A2(new_n377), .B1(G125), .B2(new_n373), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n372), .B1(new_n260), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G237), .ZN(new_n380));
  INV_X1    g194(.A(G953), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G214), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n257), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT18), .A2(G131), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(G131), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n382), .B(G143), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n321), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT16), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n376), .B2(G140), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n260), .B(new_n393), .C1(new_n378), .C2(new_n392), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n378), .B2(new_n392), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G146), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n383), .A2(KEYINPUT17), .A3(G131), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n391), .A2(new_n394), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G113), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n207), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n386), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n386), .B2(new_n398), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n369), .B1(new_n403), .B2(new_n363), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n387), .A2(new_n389), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT19), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n371), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n406), .B2(new_n378), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n396), .B(new_n405), .C1(new_n408), .C2(G146), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n400), .B1(new_n409), .B2(new_n386), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n369), .B(new_n363), .C1(new_n410), .C2(new_n401), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(KEYINPUT20), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(KEYINPUT20), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n404), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n415));
  XNOR2_X1  g229(.A(G128), .B(G143), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT13), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n254), .A2(KEYINPUT13), .A3(G143), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(new_n314), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n417), .A2(new_n419), .B1(new_n314), .B2(new_n416), .ZN(new_n420));
  INV_X1    g234(.A(G122), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G116), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n191), .A2(G122), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n425));
  XNOR2_X1  g239(.A(G116), .B(G122), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n425), .A2(new_n428), .A3(new_n211), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n211), .B1(new_n425), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n420), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n432));
  OAI211_X1 g246(.A(G107), .B(new_n432), .C1(new_n424), .C2(KEYINPUT14), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n416), .B(new_n314), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT14), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n426), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n438), .A2(KEYINPUT86), .A3(G107), .A4(new_n432), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n425), .A2(new_n428), .A3(new_n211), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n435), .A2(new_n436), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G217), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n306), .A2(new_n443), .A3(G953), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n431), .B2(new_n441), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n415), .B(new_n361), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n361), .B1(new_n446), .B2(new_n447), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT87), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT15), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n451), .A2(KEYINPUT88), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(KEYINPUT88), .ZN(new_n453));
  OAI21_X1  g267(.A(G478), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(KEYINPUT87), .B2(KEYINPUT89), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n448), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n449), .B2(KEYINPUT89), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n414), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G952), .ZN(new_n460));
  AOI211_X1 g274(.A(G953), .B(new_n460), .C1(G234), .C2(G237), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n381), .B(new_n361), .C1(G234), .C2(G237), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT21), .B(G898), .Z(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n304), .A2(new_n368), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT23), .B1(new_n254), .B2(G119), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n254), .A2(G119), .ZN(new_n471));
  MUX2_X1   g285(.A(KEYINPUT23), .B(new_n470), .S(new_n471), .Z(new_n472));
  XNOR2_X1  g286(.A(G119), .B(G128), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT24), .B(G110), .Z(new_n474));
  OAI22_X1  g288(.A1(new_n472), .A2(G110), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n396), .A3(new_n372), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n396), .A2(new_n394), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n472), .A2(G110), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(KEYINPUT72), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(KEYINPUT72), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT22), .B(G137), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n381), .A2(G221), .A3(G234), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n476), .B(new_n485), .C1(new_n480), .C2(new_n481), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n361), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT25), .A4(new_n361), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n443), .B1(new_n361), .B2(G234), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n487), .A2(new_n488), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n494), .A2(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n314), .A2(G137), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n316), .A2(G134), .ZN(new_n501));
  OAI21_X1  g315(.A(G131), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n322), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n336), .A2(new_n323), .B1(new_n262), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n504), .A2(KEYINPUT64), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n262), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n338), .B2(new_n272), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT64), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT30), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n206), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n206), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT26), .B(G101), .Z(new_n514));
  NAND3_X1  g328(.A1(new_n380), .A2(new_n381), .A3(G210), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  INV_X1    g334(.A(new_n518), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n508), .A2(new_n206), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT28), .B1(new_n504), .B2(new_n512), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G472), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n511), .A2(KEYINPUT31), .A3(new_n513), .A4(new_n518), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n363), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT32), .B1(new_n530), .B2(KEYINPUT68), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n513), .A2(new_n523), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n525), .B1(new_n535), .B2(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n518), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n505), .B1(new_n504), .B2(KEYINPUT64), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT30), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n512), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n513), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(new_n518), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n361), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(KEYINPUT29), .A3(new_n518), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n536), .A2(KEYINPUT69), .A3(KEYINPUT29), .A4(new_n518), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G472), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n499), .B1(new_n534), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n469), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(new_n221), .Z(G3));
  NAND2_X1  g369(.A1(new_n252), .A2(new_n277), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n363), .A3(new_n288), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n294), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n302), .B1(new_n558), .B2(new_n298), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(new_n466), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n493), .A2(new_n494), .B1(new_n497), .B2(new_n496), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n527), .A2(new_n361), .A3(new_n529), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G472), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n530), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n308), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n362), .A2(new_n367), .ZN(new_n567));
  AND4_X1   g381(.A1(new_n561), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n450), .A2(new_n570), .A3(new_n448), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n446), .B2(new_n447), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n572), .B(KEYINPUT33), .C1(new_n446), .C2(new_n447), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n360), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n571), .B1(new_n577), .B2(new_n570), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n571), .C1(new_n577), .C2(new_n570), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n414), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT92), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT34), .B(G104), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G6));
  INV_X1    g402(.A(new_n404), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n412), .A2(new_n590), .A3(new_n413), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n412), .B2(new_n413), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n458), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n569), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G107), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G9));
  NOR2_X1   g411(.A1(new_n486), .A2(KEYINPUT36), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n482), .B(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n493), .A2(new_n494), .B1(new_n497), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n469), .A2(new_n565), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT95), .B(G110), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G12));
  INV_X1    g420(.A(new_n533), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n552), .B1(new_n607), .B2(new_n531), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n608), .A2(new_n559), .A3(new_n368), .A4(new_n601), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT96), .B(G900), .Z(new_n610));
  AOI21_X1  g424(.A(new_n461), .B1(new_n463), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n594), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n254), .ZN(G30));
  XOR2_X1   g429(.A(new_n611), .B(KEYINPUT39), .Z(new_n616));
  NAND2_X1  g430(.A1(new_n368), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT97), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n600), .B1(new_n619), .B2(KEYINPUT40), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n544), .A2(new_n521), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n363), .B1(new_n535), .B2(new_n518), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n534), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n414), .A2(new_n458), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n625), .B(new_n626), .C1(new_n618), .C2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n300), .B(KEYINPUT38), .ZN(new_n629));
  OR4_X1    g443(.A1(new_n302), .A2(new_n620), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G143), .ZN(G45));
  INV_X1    g445(.A(new_n414), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n582), .A2(new_n632), .A3(new_n612), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n609), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G146), .ZN(G48));
  NAND2_X1  g451(.A1(new_n358), .A2(new_n361), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G469), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n639), .A2(new_n566), .A3(new_n362), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n560), .A2(new_n553), .A3(new_n584), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT41), .B(G113), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(G15));
  AND3_X1   g458(.A1(new_n640), .A2(new_n608), .A3(new_n559), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n499), .A2(new_n467), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n594), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G116), .ZN(G18));
  NAND4_X1  g462(.A1(new_n645), .A2(KEYINPUT100), .A3(new_n468), .A4(new_n601), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n640), .A2(new_n608), .A3(new_n559), .A4(new_n468), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(new_n600), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G119), .ZN(G21));
  AND2_X1   g468(.A1(new_n640), .A2(new_n559), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n530), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n530), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n563), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n655), .A2(new_n626), .A3(new_n646), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G122), .ZN(G24));
  NOR3_X1   g476(.A1(new_n633), .A2(new_n659), .A3(new_n600), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G125), .ZN(G27));
  INV_X1    g479(.A(new_n302), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n297), .A2(new_n299), .A3(new_n666), .ZN(new_n667));
  AOI211_X1 g481(.A(G469), .B(new_n360), .C1(new_n353), .C2(new_n357), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n365), .A2(new_n346), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n347), .A2(new_n355), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(G469), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n364), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT102), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n362), .A2(new_n367), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n566), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT103), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n674), .A2(new_n679), .A3(new_n676), .A4(new_n566), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n667), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n633), .A2(KEYINPUT42), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n553), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n667), .A2(new_n678), .A3(new_n680), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n685));
  NAND2_X1  g499(.A1(KEYINPUT104), .A2(KEYINPUT32), .ZN(new_n686));
  NOR2_X1   g500(.A1(KEYINPUT104), .A2(KEYINPUT32), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n530), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n552), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n687), .B1(new_n530), .B2(new_n686), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n685), .B(new_n561), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n530), .A2(new_n686), .ZN(new_n693));
  INV_X1    g507(.A(new_n687), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n552), .A3(new_n688), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n685), .B1(new_n696), .B2(new_n561), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n684), .A2(new_n698), .A3(new_n633), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n683), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n321), .ZN(G33));
  INV_X1    g516(.A(new_n613), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n681), .A2(KEYINPUT106), .A3(new_n553), .A4(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n667), .A2(new_n678), .A3(new_n553), .A4(new_n680), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n705), .B1(new_n706), .B2(new_n613), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  OR2_X1    g523(.A1(new_n366), .A2(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n366), .A2(KEYINPUT45), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(G469), .A3(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(new_n672), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT46), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT107), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n668), .B1(new_n714), .B2(KEYINPUT107), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n713), .B2(KEYINPUT46), .ZN(new_n718));
  OR3_X1    g532(.A1(new_n713), .A2(new_n717), .A3(KEYINPUT46), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n716), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n720), .A2(new_n566), .A3(new_n616), .ZN(new_n721));
  INV_X1    g535(.A(new_n667), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n582), .A2(new_n414), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT43), .Z(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n564), .A3(new_n601), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n726), .B2(KEYINPUT44), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n721), .B(new_n727), .C1(KEYINPUT44), .C2(new_n726), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G137), .ZN(G39));
  AND2_X1   g543(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n720), .B2(new_n566), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n720), .A2(new_n566), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(KEYINPUT109), .B2(KEYINPUT47), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n732), .B1(new_n734), .B2(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n499), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n736), .A2(new_n608), .A3(new_n633), .A4(new_n722), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n373), .ZN(G42));
  AND2_X1   g552(.A1(new_n724), .A2(new_n461), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n561), .A3(new_n660), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n655), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n667), .A2(new_n663), .A3(new_n678), .A4(new_n680), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n589), .B(new_n612), .C1(new_n591), .C2(new_n592), .ZN(new_n743));
  INV_X1    g557(.A(new_n458), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n600), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n667), .A2(new_n608), .A3(new_n745), .A4(new_n368), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n708), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT112), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n708), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n632), .A2(new_n744), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n583), .B2(new_n632), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n304), .A2(new_n568), .A3(new_n466), .A4(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n602), .A2(new_n554), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT117), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n653), .A2(new_n641), .A3(new_n647), .A4(new_n661), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n701), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n664), .B1(new_n613), .B2(new_n609), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n624), .A2(new_n601), .A3(new_n611), .ZN(new_n763));
  INV_X1    g577(.A(new_n677), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n559), .A2(new_n626), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n636), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT52), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n636), .A2(new_n769), .A3(new_n762), .A4(new_n766), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n768), .A2(KEYINPUT114), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT114), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n753), .A2(KEYINPUT117), .A3(new_n757), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n760), .A2(KEYINPUT53), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n701), .A2(new_n759), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n753), .A2(KEYINPUT113), .A3(new_n778), .A4(new_n757), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n751), .B1(new_n708), .B2(new_n748), .ZN(new_n780));
  AOI211_X1 g594(.A(KEYINPUT112), .B(new_n747), .C1(new_n704), .C2(new_n707), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n778), .B(new_n757), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n768), .A2(new_n770), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n779), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n787), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n775), .B(new_n777), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n773), .A2(new_n784), .A3(new_n779), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n788), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n786), .A2(new_n788), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(KEYINPUT115), .A3(new_n788), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n741), .B(new_n791), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n629), .A2(new_n302), .A3(new_n640), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT119), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n740), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n803), .A2(KEYINPUT120), .A3(KEYINPUT50), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n639), .A2(new_n362), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT110), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n566), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n667), .B(new_n740), .C1(new_n735), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n667), .A2(new_n640), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n809), .A2(new_n625), .A3(new_n499), .A4(new_n462), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n414), .A3(new_n583), .ZN(new_n811));
  INV_X1    g625(.A(new_n809), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n739), .A2(new_n601), .A3(new_n660), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n804), .A2(new_n808), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(KEYINPUT120), .B(KEYINPUT50), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n808), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  OAI22_X1  g634(.A1(new_n814), .A2(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n460), .A2(G953), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n584), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n739), .A2(new_n812), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n698), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT48), .Z(new_n827));
  AND3_X1   g641(.A1(new_n804), .A2(new_n808), .A3(new_n813), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n820), .B1(new_n808), .B2(new_n818), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n811), .A4(new_n816), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n823), .A2(new_n824), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n800), .A2(new_n831), .B1(G952), .B2(G953), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n806), .B(KEYINPUT49), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n303), .A3(new_n625), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n723), .A2(new_n499), .A3(new_n308), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n629), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT111), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n832), .A2(new_n837), .ZN(G75));
  XNOR2_X1  g652(.A(new_n252), .B(new_n277), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT55), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n775), .B1(new_n789), .B2(new_n790), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n360), .A3(new_n294), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n840), .B1(new_n844), .B2(KEYINPUT122), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n846));
  INV_X1    g660(.A(new_n840), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n846), .B(new_n847), .C1(new_n842), .C2(new_n843), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n846), .A3(new_n843), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n381), .A2(G952), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n845), .A2(new_n848), .A3(new_n852), .ZN(G51));
  NAND2_X1  g667(.A1(new_n672), .A2(KEYINPUT57), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n672), .A2(KEYINPUT57), .ZN(new_n855));
  INV_X1    g669(.A(new_n790), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n777), .B1(new_n858), .B2(new_n775), .ZN(new_n859));
  INV_X1    g673(.A(new_n791), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n854), .B(new_n855), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n358), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n841), .A2(new_n360), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(new_n712), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n850), .B1(new_n862), .B2(new_n864), .ZN(G54));
  NAND4_X1  g679(.A1(new_n841), .A2(KEYINPUT58), .A3(G475), .A4(new_n360), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n410), .A2(new_n401), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n866), .A2(KEYINPUT123), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n851), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT123), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G60));
  NAND2_X1  g685(.A1(new_n575), .A2(new_n576), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n791), .B1(new_n798), .B2(new_n799), .ZN(new_n873));
  NAND2_X1  g687(.A1(G478), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT59), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n872), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n841), .A2(new_n776), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n878), .B2(new_n791), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n876), .A2(new_n850), .A3(new_n879), .ZN(G63));
  NAND2_X1  g694(.A1(G217), .A2(G902), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT60), .Z(new_n882));
  NAND2_X1  g696(.A1(new_n841), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n496), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(KEYINPUT124), .A3(new_n851), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n841), .A2(new_n599), .A3(new_n882), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n851), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n850), .B1(new_n883), .B2(new_n884), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n887), .C1(KEYINPUT124), .C2(KEYINPUT61), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(G66));
  AOI21_X1  g707(.A(new_n381), .B1(new_n465), .B2(G224), .ZN(new_n894));
  INV_X1    g708(.A(new_n757), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(new_n759), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n896), .B2(new_n381), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n292), .B(new_n244), .C1(G898), .C2(new_n381), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n897), .B(new_n898), .Z(G69));
  NOR2_X1   g713(.A1(new_n343), .A2(new_n381), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n506), .A2(new_n510), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(new_n408), .Z(new_n903));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n737), .B1(KEYINPUT125), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n630), .A2(new_n636), .A3(new_n762), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(KEYINPUT125), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n906), .B(new_n907), .Z(new_n908));
  NAND4_X1  g722(.A1(new_n618), .A2(new_n553), .A3(new_n667), .A4(new_n755), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n905), .A2(new_n908), .A3(new_n728), .A4(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n901), .B(new_n903), .C1(new_n910), .C2(G953), .ZN(new_n911));
  INV_X1    g725(.A(new_n708), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n737), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n636), .A3(new_n762), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n721), .B(new_n765), .C1(new_n692), .C2(new_n697), .ZN(new_n915));
  INV_X1    g729(.A(new_n701), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n728), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n914), .A2(G953), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n381), .A2(G900), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n900), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n911), .B1(new_n920), .B2(new_n903), .ZN(G72));
  OAI211_X1 g735(.A(new_n795), .B(new_n797), .C1(new_n788), .C2(new_n786), .ZN(new_n922));
  NAND2_X1  g736(.A1(G472), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT63), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n545), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n519), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT126), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT127), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n924), .B1(new_n910), .B2(new_n896), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n850), .B1(new_n931), .B2(new_n621), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n914), .A2(new_n896), .A3(new_n917), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n544), .B1(new_n933), .B2(new_n925), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n518), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n930), .A2(new_n935), .ZN(G57));
endmodule


