

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776;

  XNOR2_X1 U366 ( .A(n453), .B(KEYINPUT19), .ZN(n609) );
  NOR2_X1 U367 ( .A1(n574), .A2(n388), .ZN(n387) );
  AND2_X2 U368 ( .A1(n613), .A2(n555), .ZN(n453) );
  NAND2_X2 U369 ( .A1(n395), .A2(n415), .ZN(n394) );
  AND2_X1 U370 ( .A1(n428), .A2(n439), .ZN(n438) );
  NAND2_X1 U371 ( .A1(n438), .A2(n437), .ZN(n457) );
  BUF_X1 U372 ( .A(n574), .Z(n408) );
  AND2_X1 U373 ( .A1(n434), .A2(n461), .ZN(n433) );
  XNOR2_X1 U374 ( .A(n422), .B(n420), .ZN(n775) );
  NOR2_X1 U375 ( .A1(n603), .A2(KEYINPUT47), .ZN(n604) );
  XNOR2_X1 U376 ( .A(n627), .B(n628), .ZN(n458) );
  NOR2_X1 U377 ( .A1(n560), .A2(n699), .ZN(n462) );
  INV_X1 U378 ( .A(n616), .ZN(n560) );
  AND2_X1 U379 ( .A1(n598), .A2(n597), .ZN(n633) );
  XNOR2_X1 U380 ( .A(n577), .B(n576), .ZN(n639) );
  NAND2_X1 U381 ( .A1(n681), .A2(n680), .ZN(n577) );
  XNOR2_X1 U382 ( .A(n651), .B(n654), .ZN(n655) );
  XNOR2_X1 U383 ( .A(n410), .B(n411), .ZN(n613) );
  INV_X1 U384 ( .A(n701), .ZN(n596) );
  XNOR2_X1 U385 ( .A(n504), .B(n503), .ZN(n567) );
  NOR2_X1 U386 ( .A1(n550), .A2(n480), .ZN(n481) );
  XNOR2_X1 U387 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n484) );
  XNOR2_X1 U388 ( .A(KEYINPUT67), .B(G101), .ZN(n536) );
  AND2_X1 U389 ( .A1(n343), .A2(n344), .ZN(n623) );
  NOR2_X1 U390 ( .A1(n612), .A2(n611), .ZN(n343) );
  AND2_X1 U391 ( .A1(n669), .A2(n622), .ZN(n344) );
  NOR2_X1 U392 ( .A1(n599), .A2(n625), .ZN(n600) );
  NAND2_X1 U393 ( .A1(n457), .A2(n736), .ZN(n345) );
  XNOR2_X1 U394 ( .A(n482), .B(n357), .ZN(n346) );
  NAND2_X1 U395 ( .A1(n457), .A2(n736), .ZN(n456) );
  XNOR2_X1 U396 ( .A(n482), .B(n357), .ZN(n563) );
  XNOR2_X2 U397 ( .A(n456), .B(n459), .ZN(n406) );
  XNOR2_X2 U398 ( .A(n345), .B(n459), .ZN(n407) );
  XNOR2_X2 U399 ( .A(n498), .B(G134), .ZN(n513) );
  NAND2_X1 U400 ( .A1(n349), .A2(n575), .ZN(n383) );
  NAND2_X1 U401 ( .A1(n397), .A2(G953), .ZN(n548) );
  XNOR2_X1 U402 ( .A(n393), .B(n423), .ZN(n392) );
  NAND2_X1 U403 ( .A1(n566), .A2(n567), .ZN(n635) );
  INV_X1 U404 ( .A(KEYINPUT66), .ZN(n427) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n533) );
  OR2_X1 U406 ( .A1(n573), .A2(n572), .ZN(n347) );
  OR2_X1 U407 ( .A1(n560), .A2(n701), .ZN(n573) );
  NAND2_X1 U408 ( .A1(n372), .A2(n371), .ZN(n370) );
  NOR2_X1 U409 ( .A1(n776), .A2(n775), .ZN(n636) );
  NOR2_X1 U410 ( .A1(n591), .A2(n590), .ZN(n413) );
  NOR2_X1 U411 ( .A1(n362), .A2(n425), .ZN(n591) );
  XNOR2_X1 U412 ( .A(G113), .B(KEYINPUT72), .ZN(n467) );
  XNOR2_X1 U413 ( .A(KEYINPUT4), .B(G146), .ZN(n409) );
  XNOR2_X1 U414 ( .A(n361), .B(G143), .ZN(n498) );
  XNOR2_X1 U415 ( .A(G128), .B(KEYINPUT81), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n450), .B(n449), .ZN(n448) );
  XNOR2_X1 U417 ( .A(G116), .B(G107), .ZN(n449) );
  XNOR2_X1 U418 ( .A(n451), .B(G122), .ZN(n450) );
  INV_X1 U419 ( .A(KEYINPUT7), .ZN(n451) );
  XNOR2_X1 U420 ( .A(n447), .B(n446), .ZN(n445) );
  XNOR2_X1 U421 ( .A(KEYINPUT9), .B(KEYINPUT96), .ZN(n447) );
  XNOR2_X1 U422 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n446) );
  XNOR2_X1 U423 ( .A(n634), .B(KEYINPUT39), .ZN(n640) );
  AND2_X1 U424 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U425 ( .A(n554), .B(n455), .ZN(n454) );
  XNOR2_X1 U426 ( .A(n635), .B(KEYINPUT100), .ZN(n677) );
  XNOR2_X1 U427 ( .A(n405), .B(n404), .ZN(n403) );
  AND2_X1 U428 ( .A1(n647), .A2(G953), .ZN(n746) );
  XNOR2_X1 U429 ( .A(n579), .B(n358), .ZN(n382) );
  INV_X1 U430 ( .A(n426), .ZN(n388) );
  AND2_X1 U431 ( .A1(n425), .A2(KEYINPUT66), .ZN(n424) );
  INV_X1 U432 ( .A(n382), .ZN(n379) );
  INV_X1 U433 ( .A(KEYINPUT65), .ZN(n443) );
  INV_X1 U434 ( .A(n547), .ZN(n397) );
  INV_X1 U435 ( .A(G237), .ZN(n473) );
  NAND2_X1 U436 ( .A1(n375), .A2(n374), .ZN(n366) );
  NAND2_X1 U437 ( .A1(n519), .A2(G902), .ZN(n374) );
  INV_X1 U438 ( .A(KEYINPUT48), .ZN(n423) );
  NAND2_X1 U439 ( .A1(n442), .A2(n440), .ZN(n439) );
  NAND2_X1 U440 ( .A1(n643), .A2(n443), .ZN(n442) );
  NAND2_X1 U441 ( .A1(n472), .A2(n441), .ZN(n440) );
  NAND2_X1 U442 ( .A1(n443), .A2(KEYINPUT2), .ZN(n441) );
  XOR2_X1 U443 ( .A(G122), .B(G104), .Z(n491) );
  XNOR2_X1 U444 ( .A(G113), .B(G143), .ZN(n490) );
  INV_X1 U445 ( .A(KEYINPUT69), .ZN(n483) );
  XNOR2_X1 U446 ( .A(n417), .B(n488), .ZN(n493) );
  XNOR2_X1 U447 ( .A(n489), .B(n418), .ZN(n417) );
  INV_X1 U448 ( .A(KEYINPUT95), .ZN(n418) );
  XNOR2_X1 U449 ( .A(n430), .B(KEYINPUT17), .ZN(n429) );
  NAND2_X1 U450 ( .A1(n398), .A2(G224), .ZN(n430) );
  XNOR2_X1 U451 ( .A(n536), .B(KEYINPUT73), .ZN(n389) );
  NAND2_X1 U452 ( .A1(G234), .A2(G237), .ZN(n476) );
  XOR2_X1 U453 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n477) );
  XNOR2_X1 U454 ( .A(n625), .B(n624), .ZN(n376) );
  NAND2_X1 U455 ( .A1(n436), .A2(n460), .ZN(n435) );
  NOR2_X1 U456 ( .A1(n347), .A2(KEYINPUT32), .ZN(n460) );
  OR2_X1 U457 ( .A1(n370), .A2(n368), .ZN(n364) );
  INV_X2 U458 ( .A(G953), .ZN(n398) );
  NAND2_X1 U459 ( .A1(n353), .A2(n416), .ZN(n415) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n755) );
  XNOR2_X1 U461 ( .A(G107), .B(G104), .ZN(n391) );
  XNOR2_X1 U462 ( .A(KEYINPUT80), .B(G110), .ZN(n390) );
  XNOR2_X1 U463 ( .A(KEYINPUT16), .B(G122), .ZN(n469) );
  INV_X1 U464 ( .A(G146), .ZN(n487) );
  XNOR2_X1 U465 ( .A(G119), .B(G137), .ZN(n520) );
  XOR2_X1 U466 ( .A(G110), .B(G128), .Z(n521) );
  INV_X1 U467 ( .A(KEYINPUT64), .ZN(n459) );
  AND2_X1 U468 ( .A1(n454), .A2(n555), .ZN(n614) );
  INV_X1 U469 ( .A(KEYINPUT99), .ZN(n576) );
  NOR2_X1 U470 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U471 ( .A(n605), .B(KEYINPUT6), .ZN(n572) );
  AND2_X1 U472 ( .A1(n396), .A2(G953), .ZN(n479) );
  XNOR2_X1 U473 ( .A(n448), .B(n445), .ZN(n501) );
  XNOR2_X1 U474 ( .A(n378), .B(n377), .ZN(n776) );
  XNOR2_X1 U475 ( .A(n630), .B(KEYINPUT105), .ZN(n377) );
  NOR2_X1 U476 ( .A1(n458), .A2(n629), .ZN(n378) );
  XNOR2_X1 U477 ( .A(n421), .B(KEYINPUT40), .ZN(n420) );
  OR2_X1 U478 ( .A1(n640), .A2(n635), .ZN(n422) );
  INV_X1 U479 ( .A(KEYINPUT104), .ZN(n421) );
  NAND2_X1 U480 ( .A1(n617), .A2(n616), .ZN(n669) );
  INV_X1 U481 ( .A(KEYINPUT60), .ZN(n400) );
  NAND2_X1 U482 ( .A1(n403), .A2(n402), .ZN(n401) );
  INV_X1 U483 ( .A(n746), .ZN(n402) );
  AND2_X1 U484 ( .A1(n382), .A2(n380), .ZN(n695) );
  INV_X1 U485 ( .A(n694), .ZN(n380) );
  AND2_X1 U486 ( .A1(n365), .A2(n363), .ZN(n348) );
  AND2_X1 U487 ( .A1(n574), .A2(KEYINPUT66), .ZN(n349) );
  XOR2_X1 U488 ( .A(n526), .B(n525), .Z(n350) );
  AND2_X1 U489 ( .A1(n369), .A2(n368), .ZN(n351) );
  AND2_X1 U490 ( .A1(n435), .A2(n426), .ZN(n352) );
  XNOR2_X1 U491 ( .A(n755), .B(n389), .ZN(n516) );
  AND2_X1 U492 ( .A1(n362), .A2(n425), .ZN(n353) );
  NOR2_X1 U493 ( .A1(n713), .A2(n458), .ZN(n354) );
  AND2_X1 U494 ( .A1(n642), .A2(n641), .ZN(n355) );
  INV_X1 U495 ( .A(G902), .ZN(n371) );
  INV_X1 U496 ( .A(KEYINPUT1), .ZN(n368) );
  XOR2_X1 U497 ( .A(n570), .B(KEYINPUT35), .Z(n356) );
  XOR2_X1 U498 ( .A(KEYINPUT89), .B(KEYINPUT0), .Z(n357) );
  XNOR2_X1 U499 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n358) );
  NOR2_X1 U500 ( .A1(n376), .A2(n714), .ZN(n717) );
  AND2_X1 U501 ( .A1(n427), .A2(KEYINPUT44), .ZN(n426) );
  XNOR2_X1 U502 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  INV_X1 U503 ( .A(KEYINPUT2), .ZN(n444) );
  AND2_X1 U504 ( .A1(n472), .A2(n443), .ZN(n359) );
  AND2_X1 U505 ( .A1(KEYINPUT65), .A2(n444), .ZN(n360) );
  INV_X1 U506 ( .A(KEYINPUT44), .ZN(n425) );
  XNOR2_X1 U507 ( .A(n362), .B(G122), .ZN(G24) );
  XNOR2_X2 U508 ( .A(n571), .B(n356), .ZN(n362) );
  OR2_X1 U509 ( .A1(n662), .A2(n370), .ZN(n369) );
  INV_X1 U510 ( .A(n366), .ZN(n373) );
  OR2_X1 U511 ( .A1(n662), .A2(n364), .ZN(n363) );
  NAND2_X1 U512 ( .A1(n366), .A2(KEYINPUT1), .ZN(n365) );
  NAND2_X1 U513 ( .A1(n373), .A2(n369), .ZN(n580) );
  NAND2_X2 U514 ( .A1(n348), .A2(n367), .ZN(n616) );
  NAND2_X1 U515 ( .A1(n351), .A2(n373), .ZN(n367) );
  INV_X1 U516 ( .A(n519), .ZN(n372) );
  NAND2_X1 U517 ( .A1(n662), .A2(n519), .ZN(n375) );
  NOR2_X1 U518 ( .A1(n376), .A2(n631), .ZN(n632) );
  NAND2_X1 U519 ( .A1(n376), .A2(n714), .ZN(n716) );
  NAND2_X1 U520 ( .A1(n379), .A2(n682), .ZN(n586) );
  AND2_X1 U521 ( .A1(n382), .A2(n381), .ZN(n696) );
  INV_X1 U522 ( .A(n577), .ZN(n381) );
  NAND2_X1 U523 ( .A1(n384), .A2(n383), .ZN(n414) );
  NAND2_X1 U524 ( .A1(n433), .A2(n435), .ZN(n575) );
  AND2_X1 U525 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U526 ( .A1(n352), .A2(n433), .ZN(n385) );
  NOR2_X1 U527 ( .A1(n387), .A2(n424), .ZN(n386) );
  NAND2_X1 U528 ( .A1(n750), .A2(n766), .ZN(n399) );
  AND2_X2 U529 ( .A1(n392), .A2(n355), .ZN(n766) );
  NAND2_X1 U530 ( .A1(n638), .A2(n637), .ZN(n393) );
  XNOR2_X2 U531 ( .A(n394), .B(KEYINPUT45), .ZN(n750) );
  XNOR2_X1 U532 ( .A(n412), .B(n592), .ZN(n395) );
  NAND2_X1 U533 ( .A1(n398), .A2(G234), .ZN(n499) );
  NAND2_X1 U534 ( .A1(n398), .A2(G227), .ZN(n514) );
  INV_X1 U535 ( .A(G898), .ZN(n396) );
  NAND2_X1 U536 ( .A1(n751), .A2(n398), .ZN(n752) );
  INV_X1 U537 ( .A(n399), .ZN(n731) );
  NAND2_X1 U538 ( .A1(n399), .A2(n360), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n401), .B(n400), .ZN(G60) );
  INV_X1 U540 ( .A(n676), .ZN(n404) );
  NAND2_X1 U541 ( .A1(n406), .A2(G475), .ZN(n405) );
  XNOR2_X2 U542 ( .A(n585), .B(n584), .ZN(n682) );
  XNOR2_X1 U543 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U544 ( .A(n644), .B(KEYINPUT119), .ZN(n645) );
  XNOR2_X1 U545 ( .A(n670), .B(KEYINPUT62), .ZN(n671) );
  NOR2_X1 U546 ( .A1(n714), .A2(n605), .ZN(n593) );
  XNOR2_X1 U547 ( .A(n675), .B(KEYINPUT59), .ZN(n676) );
  NOR2_X1 U548 ( .A1(n650), .A2(n472), .ZN(n410) );
  NAND2_X1 U549 ( .A1(n474), .A2(G210), .ZN(n411) );
  OR2_X2 U550 ( .A1(n546), .A2(n545), .ZN(n574) );
  NAND2_X1 U551 ( .A1(n414), .A2(n413), .ZN(n412) );
  AND2_X1 U552 ( .A1(n408), .A2(n575), .ZN(n416) );
  NAND2_X1 U553 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X2 U554 ( .A(n562), .B(n561), .ZN(n721) );
  BUF_X1 U555 ( .A(n346), .Z(n583) );
  XNOR2_X1 U556 ( .A(n419), .B(n674), .ZN(G57) );
  NOR2_X2 U557 ( .A1(n673), .A2(n746), .ZN(n419) );
  XNOR2_X1 U558 ( .A(n431), .B(n429), .ZN(n464) );
  XNOR2_X1 U559 ( .A(n509), .B(n432), .ZN(n431) );
  XNOR2_X2 U560 ( .A(G125), .B(KEYINPUT18), .ZN(n432) );
  XNOR2_X2 U561 ( .A(G146), .B(KEYINPUT4), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n546), .A2(KEYINPUT32), .ZN(n434) );
  INV_X1 U563 ( .A(n546), .ZN(n436) );
  XNOR2_X2 U564 ( .A(n508), .B(KEYINPUT22), .ZN(n546) );
  NAND2_X1 U565 ( .A1(n731), .A2(n359), .ZN(n437) );
  NOR2_X1 U566 ( .A1(n606), .A2(n677), .ZN(n553) );
  XNOR2_X2 U567 ( .A(n497), .B(n496), .ZN(n566) );
  NAND2_X1 U568 ( .A1(n454), .A2(n453), .ZN(n452) );
  XNOR2_X1 U569 ( .A(n452), .B(n615), .ZN(n617) );
  INV_X1 U570 ( .A(KEYINPUT101), .ZN(n455) );
  NOR2_X1 U571 ( .A1(n458), .A2(n728), .ZN(n729) );
  NAND2_X1 U572 ( .A1(n407), .A2(G472), .ZN(n672) );
  NAND2_X1 U573 ( .A1(n407), .A2(G217), .ZN(n646) );
  NAND2_X1 U574 ( .A1(n407), .A2(G210), .ZN(n656) );
  NAND2_X1 U575 ( .A1(n406), .A2(G469), .ZN(n664) );
  NAND2_X1 U576 ( .A1(n406), .A2(G478), .ZN(n744) );
  NAND2_X1 U577 ( .A1(n347), .A2(KEYINPUT32), .ZN(n461) );
  XNOR2_X1 U578 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U579 ( .A(n718), .B(KEYINPUT85), .ZN(n603) );
  INV_X1 U580 ( .A(n594), .ZN(n595) );
  INV_X1 U581 ( .A(n498), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n465), .B(n516), .ZN(n471) );
  XNOR2_X1 U583 ( .A(G119), .B(G116), .ZN(n466) );
  XNOR2_X1 U584 ( .A(n466), .B(KEYINPUT3), .ZN(n468) );
  XNOR2_X1 U585 ( .A(n468), .B(n467), .ZN(n538) );
  XNOR2_X1 U586 ( .A(n469), .B(KEYINPUT76), .ZN(n470) );
  XNOR2_X1 U587 ( .A(n538), .B(n470), .ZN(n757) );
  XNOR2_X1 U588 ( .A(n471), .B(n757), .ZN(n650) );
  INV_X1 U589 ( .A(n643), .ZN(n472) );
  NAND2_X1 U590 ( .A1(n371), .A2(n473), .ZN(n474) );
  NAND2_X1 U591 ( .A1(n474), .A2(G214), .ZN(n475) );
  XNOR2_X1 U592 ( .A(n475), .B(KEYINPUT90), .ZN(n555) );
  XOR2_X1 U593 ( .A(n477), .B(n476), .Z(n478) );
  NAND2_X1 U594 ( .A1(G952), .A2(n478), .ZN(n727) );
  NOR2_X1 U595 ( .A1(n727), .A2(G953), .ZN(n550) );
  NAND2_X1 U596 ( .A1(n478), .A2(G902), .ZN(n547) );
  XNOR2_X1 U597 ( .A(KEYINPUT91), .B(n479), .ZN(n759) );
  NOR2_X1 U598 ( .A1(n547), .A2(n759), .ZN(n480) );
  NOR2_X2 U599 ( .A1(n609), .A2(n481), .ZN(n482) );
  XNOR2_X1 U600 ( .A(n483), .B(G131), .ZN(n510) );
  INV_X1 U601 ( .A(n484), .ZN(n486) );
  XNOR2_X1 U602 ( .A(G125), .B(G140), .ZN(n485) );
  XNOR2_X1 U603 ( .A(n486), .B(n485), .ZN(n765) );
  XNOR2_X1 U604 ( .A(n765), .B(n487), .ZN(n523) );
  XNOR2_X1 U605 ( .A(n510), .B(n523), .ZN(n495) );
  NAND2_X1 U606 ( .A1(G214), .A2(n533), .ZN(n489) );
  XOR2_X1 U607 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n488) );
  XNOR2_X1 U608 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U609 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U610 ( .A(n495), .B(n494), .ZN(n675) );
  NAND2_X1 U611 ( .A1(n675), .A2(n371), .ZN(n497) );
  XOR2_X1 U612 ( .A(KEYINPUT13), .B(G475), .Z(n496) );
  INV_X1 U613 ( .A(n566), .ZN(n681) );
  XOR2_X1 U614 ( .A(KEYINPUT8), .B(n499), .Z(n524) );
  NAND2_X1 U615 ( .A1(G217), .A2(n524), .ZN(n500) );
  XNOR2_X1 U616 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n513), .B(n502), .ZN(n742) );
  NAND2_X1 U618 ( .A1(n742), .A2(n371), .ZN(n504) );
  INV_X1 U619 ( .A(G478), .ZN(n503) );
  AND2_X1 U620 ( .A1(n681), .A2(n567), .ZN(n626) );
  INV_X1 U621 ( .A(n626), .ZN(n715) );
  NAND2_X1 U622 ( .A1(G234), .A2(n643), .ZN(n505) );
  XNOR2_X1 U623 ( .A(KEYINPUT20), .B(n505), .ZN(n528) );
  AND2_X1 U624 ( .A1(n528), .A2(G221), .ZN(n506) );
  XNOR2_X1 U625 ( .A(n506), .B(KEYINPUT21), .ZN(n702) );
  INV_X1 U626 ( .A(n702), .ZN(n552) );
  NOR2_X1 U627 ( .A1(n715), .A2(n552), .ZN(n507) );
  NAND2_X1 U628 ( .A1(n563), .A2(n507), .ZN(n508) );
  XNOR2_X1 U629 ( .A(n409), .B(G137), .ZN(n511) );
  XNOR2_X1 U630 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X2 U631 ( .A(n513), .B(n512), .ZN(n764) );
  XNOR2_X1 U632 ( .A(n514), .B(G140), .ZN(n515) );
  XNOR2_X1 U633 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U634 ( .A(n517), .B(n764), .ZN(n662) );
  INV_X1 U635 ( .A(KEYINPUT71), .ZN(n518) );
  XNOR2_X1 U636 ( .A(n518), .B(G469), .ZN(n519) );
  XNOR2_X1 U637 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U638 ( .A(n523), .B(n522), .ZN(n527) );
  XOR2_X1 U639 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n526) );
  NAND2_X1 U640 ( .A1(G221), .A2(n524), .ZN(n525) );
  XNOR2_X1 U641 ( .A(n527), .B(n350), .ZN(n644) );
  NAND2_X1 U642 ( .A1(n644), .A2(n371), .ZN(n532) );
  XOR2_X1 U643 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n530) );
  NAND2_X1 U644 ( .A1(n528), .A2(G217), .ZN(n529) );
  XNOR2_X1 U645 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X2 U646 ( .A(n532), .B(n531), .ZN(n701) );
  OR2_X1 U647 ( .A1(n616), .A2(n596), .ZN(n542) );
  NAND2_X1 U648 ( .A1(G210), .A2(n533), .ZN(n534) );
  XNOR2_X1 U649 ( .A(n534), .B(KEYINPUT5), .ZN(n535) );
  XNOR2_X1 U650 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U651 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U652 ( .A(n764), .B(n539), .ZN(n670) );
  OR2_X2 U653 ( .A1(n670), .A2(G902), .ZN(n541) );
  INV_X1 U654 ( .A(G472), .ZN(n540) );
  XNOR2_X2 U655 ( .A(n541), .B(n540), .ZN(n605) );
  OR2_X1 U656 ( .A1(n542), .A2(n572), .ZN(n543) );
  OR2_X1 U657 ( .A1(n546), .A2(n543), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n588), .B(G101), .ZN(G3) );
  INV_X1 U659 ( .A(n605), .ZN(n704) );
  NOR2_X1 U660 ( .A1(n701), .A2(n704), .ZN(n544) );
  NAND2_X1 U661 ( .A1(n560), .A2(n544), .ZN(n545) );
  XNOR2_X1 U662 ( .A(n408), .B(G110), .ZN(G12) );
  NOR2_X1 U663 ( .A1(n548), .A2(G900), .ZN(n549) );
  NOR2_X1 U664 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U665 ( .A1(n552), .A2(n551), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n596), .A2(n594), .ZN(n606) );
  AND2_X1 U667 ( .A1(n553), .A2(n572), .ZN(n554) );
  INV_X1 U668 ( .A(n555), .ZN(n714) );
  XNOR2_X1 U669 ( .A(n614), .B(KEYINPUT102), .ZN(n556) );
  AND2_X1 U670 ( .A1(n556), .A2(n560), .ZN(n558) );
  INV_X1 U671 ( .A(KEYINPUT43), .ZN(n557) );
  XNOR2_X1 U672 ( .A(n558), .B(n557), .ZN(n559) );
  INV_X1 U673 ( .A(n613), .ZN(n625) );
  NAND2_X1 U674 ( .A1(n559), .A2(n625), .ZN(n642) );
  XNOR2_X1 U675 ( .A(n642), .B(G140), .ZN(G42) );
  NAND2_X1 U676 ( .A1(n701), .A2(n702), .ZN(n699) );
  NAND2_X1 U677 ( .A1(n462), .A2(n572), .ZN(n562) );
  XNOR2_X1 U678 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n561) );
  NAND2_X1 U679 ( .A1(n721), .A2(n346), .ZN(n565) );
  XNOR2_X1 U680 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n564) );
  XNOR2_X1 U681 ( .A(n565), .B(n564), .ZN(n569) );
  INV_X1 U682 ( .A(n567), .ZN(n680) );
  NAND2_X1 U683 ( .A1(n566), .A2(n680), .ZN(n602) );
  INV_X1 U684 ( .A(n602), .ZN(n568) );
  INV_X1 U685 ( .A(KEYINPUT87), .ZN(n570) );
  XNOR2_X1 U686 ( .A(n575), .B(G119), .ZN(G21) );
  NAND2_X1 U687 ( .A1(n635), .A2(n639), .ZN(n718) );
  INV_X1 U688 ( .A(n603), .ZN(n587) );
  NOR2_X1 U689 ( .A1(n699), .A2(n605), .ZN(n578) );
  AND2_X1 U690 ( .A1(n616), .A2(n578), .ZN(n708) );
  NAND2_X1 U691 ( .A1(n583), .A2(n708), .ZN(n579) );
  INV_X1 U692 ( .A(n580), .ZN(n631) );
  OR2_X1 U693 ( .A1(n699), .A2(n631), .ZN(n581) );
  NOR2_X1 U694 ( .A1(n581), .A2(n704), .ZN(n582) );
  NAND2_X1 U695 ( .A1(n583), .A2(n582), .ZN(n585) );
  INV_X1 U696 ( .A(KEYINPUT93), .ZN(n584) );
  NAND2_X1 U697 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U698 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U699 ( .A(KEYINPUT88), .ZN(n592) );
  XNOR2_X1 U700 ( .A(n593), .B(KEYINPUT30), .ZN(n598) );
  NAND2_X1 U701 ( .A1(n633), .A2(n580), .ZN(n599) );
  XNOR2_X1 U702 ( .A(n600), .B(KEYINPUT103), .ZN(n601) );
  NOR2_X1 U703 ( .A1(n602), .A2(n601), .ZN(n689) );
  XNOR2_X1 U704 ( .A(n689), .B(KEYINPUT86), .ZN(n612) );
  XNOR2_X1 U705 ( .A(n604), .B(KEYINPUT77), .ZN(n610) );
  NOR2_X1 U706 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U707 ( .A(n607), .B(KEYINPUT28), .ZN(n608) );
  NAND2_X1 U708 ( .A1(n608), .A2(n580), .ZN(n629) );
  OR2_X1 U709 ( .A1(n629), .A2(n609), .ZN(n691) );
  NOR2_X1 U710 ( .A1(n610), .A2(n691), .ZN(n611) );
  XOR2_X1 U711 ( .A(KEYINPUT106), .B(KEYINPUT36), .Z(n615) );
  INV_X1 U712 ( .A(n718), .ZN(n618) );
  NAND2_X1 U713 ( .A1(n618), .A2(KEYINPUT47), .ZN(n619) );
  XNOR2_X1 U714 ( .A(n619), .B(KEYINPUT84), .ZN(n621) );
  NAND2_X1 U715 ( .A1(n691), .A2(KEYINPUT47), .ZN(n620) );
  AND2_X1 U716 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U717 ( .A(n623), .B(KEYINPUT70), .ZN(n638) );
  INV_X1 U718 ( .A(KEYINPUT42), .ZN(n630) );
  INV_X1 U719 ( .A(KEYINPUT41), .ZN(n628) );
  XNOR2_X1 U720 ( .A(KEYINPUT38), .B(KEYINPUT79), .ZN(n624) );
  NAND2_X1 U721 ( .A1(n626), .A2(n717), .ZN(n627) );
  XNOR2_X1 U722 ( .A(n636), .B(KEYINPUT46), .ZN(n637) );
  NOR2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n697) );
  INV_X1 U724 ( .A(n697), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n731), .A2(KEYINPUT2), .ZN(n736) );
  XNOR2_X1 U726 ( .A(n646), .B(n645), .ZN(n648) );
  INV_X1 U727 ( .A(G952), .ZN(n647) );
  NOR2_X2 U728 ( .A1(n648), .A2(n746), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT120), .ZN(G66) );
  BUF_X1 U730 ( .A(n650), .Z(n651) );
  XOR2_X1 U731 ( .A(KEYINPUT55), .B(KEYINPUT82), .Z(n653) );
  XNOR2_X1 U732 ( .A(KEYINPUT114), .B(KEYINPUT54), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  NOR2_X2 U735 ( .A1(n657), .A2(n746), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n658), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U737 ( .A(KEYINPUT116), .B(KEYINPUT57), .ZN(n660) );
  XNOR2_X1 U738 ( .A(KEYINPUT58), .B(KEYINPUT115), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n665) );
  NOR2_X2 U741 ( .A1(n665), .A2(n746), .ZN(n667) );
  INV_X1 U742 ( .A(KEYINPUT117), .ZN(n666) );
  XNOR2_X1 U743 ( .A(n667), .B(n666), .ZN(G54) );
  XOR2_X1 U744 ( .A(G125), .B(KEYINPUT37), .Z(n668) );
  XNOR2_X1 U745 ( .A(n669), .B(n668), .ZN(G27) );
  INV_X1 U746 ( .A(KEYINPUT63), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n672), .B(n671), .ZN(n673) );
  BUF_X1 U748 ( .A(n677), .Z(n694) );
  NOR2_X1 U749 ( .A1(n694), .A2(n682), .ZN(n679) );
  XNOR2_X1 U750 ( .A(G104), .B(KEYINPUT107), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n679), .B(n678), .ZN(G6) );
  NOR2_X1 U752 ( .A1(n577), .A2(n682), .ZN(n684) );
  XNOR2_X1 U753 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n683) );
  XNOR2_X1 U754 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U755 ( .A(G107), .B(n685), .ZN(G9) );
  NOR2_X1 U756 ( .A1(n691), .A2(n577), .ZN(n687) );
  XNOR2_X1 U757 ( .A(KEYINPUT29), .B(KEYINPUT108), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U759 ( .A(G128), .B(n688), .ZN(G30) );
  XNOR2_X1 U760 ( .A(n689), .B(G143), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(KEYINPUT109), .ZN(G45) );
  NOR2_X1 U762 ( .A1(n694), .A2(n691), .ZN(n692) );
  XOR2_X1 U763 ( .A(KEYINPUT110), .B(n692), .Z(n693) );
  XNOR2_X1 U764 ( .A(G146), .B(n693), .ZN(G48) );
  XOR2_X1 U765 ( .A(G113), .B(n695), .Z(G15) );
  XOR2_X1 U766 ( .A(G116), .B(n696), .Z(G18) );
  XOR2_X1 U767 ( .A(G134), .B(n697), .Z(G36) );
  XNOR2_X1 U768 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT51), .ZN(n712) );
  NAND2_X1 U770 ( .A1(n560), .A2(n699), .ZN(n700) );
  XNOR2_X1 U771 ( .A(n700), .B(KEYINPUT50), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U773 ( .A(KEYINPUT49), .B(n703), .Z(n705) );
  NOR2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n710) );
  INV_X1 U776 ( .A(n708), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U778 ( .A(n712), .B(n711), .Z(n713) );
  NAND2_X1 U779 ( .A1(n716), .A2(n626), .ZN(n720) );
  NAND2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  AND2_X1 U781 ( .A1(n720), .A2(n719), .ZN(n722) );
  INV_X1 U782 ( .A(n721), .ZN(n728) );
  NOR2_X1 U783 ( .A1(n722), .A2(n728), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n354), .A2(n723), .ZN(n724) );
  XOR2_X1 U785 ( .A(n724), .B(KEYINPUT113), .Z(n725) );
  XNOR2_X1 U786 ( .A(KEYINPUT52), .B(n725), .ZN(n726) );
  NOR2_X1 U787 ( .A1(n727), .A2(n726), .ZN(n730) );
  NOR2_X1 U788 ( .A1(n730), .A2(n729), .ZN(n739) );
  NOR2_X1 U789 ( .A1(n731), .A2(KEYINPUT83), .ZN(n732) );
  OR2_X1 U790 ( .A1(n732), .A2(KEYINPUT2), .ZN(n735) );
  INV_X1 U791 ( .A(KEYINPUT83), .ZN(n733) );
  NAND2_X1 U792 ( .A1(n733), .A2(KEYINPUT2), .ZN(n734) );
  NAND2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U795 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U796 ( .A1(n740), .A2(G953), .ZN(n741) );
  XNOR2_X1 U797 ( .A(n741), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U798 ( .A(KEYINPUT118), .B(n742), .Z(n743) );
  XNOR2_X1 U799 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U800 ( .A1(n746), .A2(n745), .ZN(G63) );
  XOR2_X1 U801 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n748) );
  NAND2_X1 U802 ( .A1(G224), .A2(G953), .ZN(n747) );
  XNOR2_X1 U803 ( .A(n748), .B(n747), .ZN(n749) );
  NAND2_X1 U804 ( .A1(n749), .A2(G898), .ZN(n754) );
  BUF_X1 U805 ( .A(n750), .Z(n751) );
  XNOR2_X1 U806 ( .A(n752), .B(KEYINPUT122), .ZN(n753) );
  NAND2_X1 U807 ( .A1(n754), .A2(n753), .ZN(n762) );
  XNOR2_X1 U808 ( .A(n755), .B(KEYINPUT123), .ZN(n756) );
  XNOR2_X1 U809 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n758), .B(G101), .ZN(n760) );
  NAND2_X1 U811 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U812 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U813 ( .A(KEYINPUT124), .B(n763), .Z(G69) );
  XOR2_X1 U814 ( .A(n765), .B(n764), .Z(n769) );
  XNOR2_X1 U815 ( .A(n766), .B(n769), .ZN(n767) );
  NOR2_X1 U816 ( .A1(G953), .A2(n767), .ZN(n768) );
  XNOR2_X1 U817 ( .A(n768), .B(KEYINPUT125), .ZN(n774) );
  XNOR2_X1 U818 ( .A(n769), .B(G227), .ZN(n770) );
  NAND2_X1 U819 ( .A1(n770), .A2(G900), .ZN(n771) );
  XNOR2_X1 U820 ( .A(KEYINPUT126), .B(n771), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n772), .A2(G953), .ZN(n773) );
  NAND2_X1 U822 ( .A1(n774), .A2(n773), .ZN(G72) );
  XOR2_X1 U823 ( .A(n775), .B(G131), .Z(G33) );
  XOR2_X1 U824 ( .A(G137), .B(n776), .Z(G39) );
endmodule

