//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  OAI211_X1 g003(.A(new_n188), .B(G146), .C1(new_n189), .C2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(KEYINPUT68), .A3(new_n192), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n188), .A2(G146), .ZN(new_n202));
  AND4_X1   g016(.A1(new_n197), .A2(new_n199), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n195), .B(new_n196), .C1(new_n200), .C2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G131), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(G137), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n211), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT0), .B(G128), .C1(new_n198), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n201), .A2(new_n202), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n219), .A2(KEYINPUT64), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n212), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G116), .B(G119), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n230), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n216), .A2(new_n227), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n235), .B2(new_n237), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n216), .A2(new_n227), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n233), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n235), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT28), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(G902), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n216), .A2(new_n227), .A3(KEYINPUT30), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n212), .A2(new_n215), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n190), .A2(KEYINPUT68), .A3(new_n192), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT68), .B1(new_n190), .B2(new_n192), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n198), .A2(new_n197), .A3(new_n199), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n256), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n225), .A2(new_n212), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n218), .A2(new_n222), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT66), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n223), .A2(new_n268), .A3(new_n226), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n264), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n233), .B(new_n255), .C1(new_n270), .C2(KEYINPUT30), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n235), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n251), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n235), .B1(new_n270), .B2(new_n234), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n240), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n252), .B(new_n273), .C1(new_n276), .C2(new_n251), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n187), .B1(new_n254), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n235), .A3(new_n250), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT31), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n271), .A2(new_n282), .A3(new_n235), .A4(new_n250), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n266), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n268), .B1(new_n223), .B2(new_n226), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n216), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n233), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n237), .B1(new_n288), .B2(new_n235), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n235), .A2(new_n237), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n251), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n276), .A2(KEYINPUT70), .A3(new_n251), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n284), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n298), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n281), .A2(new_n283), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT70), .B1(new_n276), .B2(new_n251), .ZN(new_n304));
  AOI211_X1 g118(.A(new_n295), .B(new_n250), .C1(new_n240), .C2(new_n275), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n302), .B1(new_n306), .B2(new_n299), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n279), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT71), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT32), .B1(new_n298), .B2(new_n300), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n302), .A3(new_n299), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n279), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(G234), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(G140), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT73), .B(G140), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(new_n320), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n319), .B(G125), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(KEYINPUT16), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(G125), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n191), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G110), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n189), .A2(G119), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n335), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n333), .A2(G128), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n338), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n342), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n320), .A2(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n329), .A2(new_n348), .A3(new_n191), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n332), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n328), .A2(new_n331), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G146), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n328), .A2(new_n191), .A3(new_n331), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n344), .A2(new_n345), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(G110), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n351), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G221), .A3(G234), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n360), .B(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT75), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n354), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n358), .B1(new_n365), .B2(new_n332), .ZN(new_n366));
  INV_X1    g180(.A(new_n351), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n369));
  INV_X1    g183(.A(new_n363), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n367), .A3(new_n363), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n359), .A2(new_n375), .A3(new_n363), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n377), .A3(new_n317), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n364), .A2(new_n371), .B1(new_n374), .B2(new_n376), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT25), .B1(new_n381), .B2(new_n317), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n318), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n318), .A2(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n315), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n318), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n378), .A2(new_n379), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n381), .A2(KEYINPUT25), .A3(new_n317), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n385), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(KEYINPUT77), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G214), .B1(G237), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n230), .A2(KEYINPUT5), .ZN(new_n396));
  INV_X1    g210(.A(G116), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n397), .A2(KEYINPUT5), .A3(G119), .ZN(new_n398));
  INV_X1    g212(.A(G113), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n396), .A2(new_n400), .B1(new_n229), .B2(new_n230), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G107), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G101), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(G107), .ZN(new_n409));
  OAI22_X1  g223(.A1(new_n402), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n412));
  INV_X1    g226(.A(G107), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G104), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G101), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n411), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n412), .B1(new_n411), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n401), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n411), .A2(KEYINPUT4), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n408), .B1(new_n421), .B2(KEYINPUT79), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n407), .A2(new_n423), .A3(new_n409), .A4(new_n410), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n414), .B1(new_n426), .B2(new_n404), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n410), .A2(new_n409), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT79), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n424), .A3(G101), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n233), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n419), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n419), .B(new_n434), .C1(new_n425), .C2(new_n432), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n204), .A2(new_n320), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n223), .A2(G125), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n361), .A2(G224), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT86), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n433), .A2(new_n445), .A3(new_n435), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n438), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(KEYINPUT7), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(G125), .B1(new_n259), .B2(new_n263), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n266), .A2(new_n320), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n439), .A2(new_n440), .A3(new_n448), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n431), .A2(new_n233), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n422), .A2(new_n424), .ZN(new_n456));
  INV_X1    g270(.A(new_n420), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n411), .A2(new_n416), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT81), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n411), .A2(new_n412), .A3(new_n416), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n455), .A2(new_n458), .B1(new_n462), .B2(new_n401), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n454), .B1(new_n463), .B2(new_n434), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n434), .B(KEYINPUT8), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n411), .A2(new_n416), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n396), .A2(KEYINPUT87), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n230), .A2(new_n468), .A3(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n400), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n470), .A3(new_n232), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n471), .A2(KEYINPUT88), .B1(new_n401), .B2(new_n466), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n471), .A2(KEYINPUT88), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n464), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n447), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n447), .A2(new_n475), .A3(new_n477), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n395), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n429), .A2(G101), .A3(new_n424), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n223), .B(new_n431), .C1(new_n482), .C2(new_n420), .ZN(new_n483));
  OAI211_X1 g297(.A(KEYINPUT10), .B(new_n204), .C1(new_n417), .C2(new_n418), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT10), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n193), .B1(new_n261), .B2(new_n262), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n459), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT83), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n483), .A2(new_n484), .A3(new_n490), .A4(new_n487), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n226), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n483), .A2(new_n484), .A3(new_n265), .A4(new_n487), .ZN(new_n493));
  XNOR2_X1  g307(.A(G110), .B(G140), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n361), .A2(G227), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n466), .A2(new_n204), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n459), .A2(new_n486), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n226), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT12), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n459), .A2(new_n263), .A3(new_n259), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n459), .B2(new_n486), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n508), .A2(KEYINPUT82), .A3(new_n503), .A4(new_n226), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n509), .A3(new_n493), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n492), .A2(new_n499), .B1(new_n510), .B2(new_n496), .ZN(new_n511));
  OAI21_X1  g325(.A(G469), .B1(new_n511), .B2(G902), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(G469), .C1(new_n511), .C2(G902), .ZN(new_n515));
  INV_X1    g329(.A(G469), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n506), .A2(new_n517), .A3(new_n509), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n506), .B2(new_n509), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n518), .A2(new_n519), .A3(new_n498), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n497), .B1(new_n492), .B2(new_n493), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n516), .B(new_n317), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT9), .B(G234), .ZN(new_n524));
  OAI21_X1  g338(.A(G221), .B1(new_n524), .B2(G902), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n349), .A2(KEYINPUT90), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n323), .A2(new_n327), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(new_n191), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n323), .A2(new_n327), .A3(new_n529), .A4(G146), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(KEYINPUT18), .B2(G131), .ZN(new_n532));
  INV_X1    g346(.A(G237), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n361), .A3(G214), .ZN(new_n534));
  NOR2_X1   g348(.A1(KEYINPUT89), .A2(G143), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(KEYINPUT89), .A2(G143), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n537), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(G214), .B2(new_n246), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n532), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(G214), .B(new_n246), .C1(new_n539), .C2(new_n535), .ZN(new_n542));
  INV_X1    g356(.A(new_n532), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n537), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n531), .A2(KEYINPUT18), .A3(G131), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n528), .A2(new_n530), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n205), .B1(new_n542), .B2(new_n544), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n205), .A3(new_n544), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(KEYINPUT94), .A3(KEYINPUT17), .ZN(new_n554));
  INV_X1    g368(.A(new_n205), .ZN(new_n555));
  OAI211_X1 g369(.A(KEYINPUT17), .B(new_n555), .C1(new_n538), .C2(new_n540), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n548), .B1(new_n355), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G113), .B(G122), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G104), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n560), .B1(KEYINPUT95), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(KEYINPUT95), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n548), .B(new_n565), .C1(new_n355), .C2(new_n559), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n317), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G475), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT20), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT92), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n527), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n323), .A2(new_n327), .A3(KEYINPUT92), .A4(KEYINPUT19), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g389(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n576));
  AND4_X1   g390(.A1(new_n329), .A2(new_n575), .A3(new_n348), .A4(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n191), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n332), .B1(new_n550), .B2(new_n552), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n548), .A2(new_n562), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n563), .A2(new_n560), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(G475), .A2(G902), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n569), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n560), .A2(new_n563), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n582), .ZN(new_n587));
  AND4_X1   g401(.A1(new_n569), .A2(new_n586), .A3(new_n587), .A4(new_n584), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n568), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n524), .A2(new_n316), .A3(G953), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  INV_X1    g409(.A(G122), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(KEYINPUT96), .A2(G122), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n397), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n596), .A2(G116), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n188), .A2(G128), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n188), .A2(G128), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n207), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n604), .ZN(new_n606));
  OAI21_X1  g420(.A(G134), .B1(new_n606), .B2(new_n602), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n601), .A2(new_n413), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n598), .ZN(new_n609));
  NOR2_X1   g423(.A1(KEYINPUT96), .A2(G122), .ZN(new_n610));
  OAI21_X1  g424(.A(G116), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n397), .A2(G122), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(KEYINPUT14), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT14), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n600), .A2(KEYINPUT98), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(KEYINPUT14), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n611), .A2(new_n614), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G107), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G107), .B1(new_n599), .B2(new_n600), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n611), .A2(new_n413), .A3(new_n613), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT13), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT97), .B1(new_n604), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n626), .A2(new_n188), .A3(KEYINPUT13), .A4(G128), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n604), .A2(new_n624), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n625), .A2(new_n627), .A3(new_n628), .A4(new_n603), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G134), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n623), .A2(new_n630), .A3(new_n605), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n594), .B1(new_n620), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n605), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n621), .B2(new_n622), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n635), .A2(new_n630), .B1(new_n608), .B2(new_n619), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n594), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n593), .B1(new_n638), .B2(new_n317), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n620), .A2(new_n631), .A3(new_n594), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n593), .B(new_n317), .C1(new_n640), .C2(new_n632), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n592), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n591), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(G234), .A2(G237), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(G952), .A3(new_n361), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n317), .B1(G234), .B2(G237), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(G953), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT21), .B(G898), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n589), .A2(new_n645), .A3(new_n653), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n481), .A2(new_n523), .A3(new_n525), .A4(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n309), .A2(new_n314), .A3(new_n393), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G101), .ZN(G3));
  NOR2_X1   g471(.A1(new_n298), .A2(new_n300), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n523), .A2(new_n525), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n393), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT33), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n640), .B2(new_n632), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n632), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT101), .B1(new_n636), .B2(new_n594), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT33), .A4(new_n637), .ZN(new_n673));
  OAI211_X1 g487(.A(KEYINPUT100), .B(new_n666), .C1(new_n640), .C2(new_n632), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n590), .A2(G902), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n669), .A2(new_n673), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n638), .A2(new_n317), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(G478), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n589), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n653), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n481), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n665), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT34), .B(G104), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G6));
  NAND3_X1  g500(.A1(new_n586), .A2(new_n587), .A3(new_n584), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT20), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n586), .A2(new_n587), .A3(new_n569), .A4(new_n584), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n689), .A2(KEYINPUT103), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n643), .A2(new_n644), .B1(G475), .B2(new_n567), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n481), .A2(new_n692), .A3(new_n682), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT104), .Z(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n665), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT35), .B(G107), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G9));
  INV_X1    g513(.A(new_n660), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n370), .A2(KEYINPUT36), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n368), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n384), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n481), .B1(new_n390), .B2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n700), .A2(new_n705), .A3(new_n658), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n523), .A2(new_n525), .A3(new_n654), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT37), .B(G110), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G12));
  NOR2_X1   g524(.A1(new_n361), .A2(G900), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n649), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(KEYINPUT105), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n647), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n693), .A2(new_n691), .A3(new_n690), .A4(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n663), .A2(new_n705), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n309), .A3(new_n314), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XNOR2_X1  g533(.A(new_n715), .B(KEYINPUT39), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n664), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n723));
  INV_X1    g537(.A(new_n272), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n251), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n317), .B1(new_n243), .B2(new_n250), .ZN(new_n726));
  OAI21_X1  g540(.A(G472), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n312), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n479), .A2(new_n480), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT38), .Z(new_n730));
  NAND2_X1  g544(.A1(new_n383), .A2(new_n703), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n589), .A2(new_n394), .A3(new_n645), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n722), .A2(new_n723), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  AOI22_X1  g549(.A1(new_n688), .A2(new_n689), .B1(G475), .B2(new_n567), .ZN(new_n736));
  INV_X1    g550(.A(new_n680), .ZN(new_n737));
  INV_X1    g551(.A(new_n715), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n739), .B(new_n481), .C1(new_n390), .C2(new_n704), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n663), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n309), .A2(new_n314), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G146), .ZN(G48));
  AOI21_X1  g557(.A(new_n313), .B1(new_n312), .B2(new_n279), .ZN(new_n744));
  AOI211_X1 g558(.A(KEYINPUT71), .B(new_n278), .C1(new_n310), .C2(new_n311), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n383), .A2(new_n385), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT77), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n390), .A2(new_n391), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n315), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n744), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n520), .A2(new_n521), .ZN(new_n753));
  OAI21_X1  g567(.A(G469), .B1(new_n753), .B2(G902), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n525), .A3(new_n522), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n683), .A2(new_n681), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT41), .B(G113), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G15));
  NAND2_X1  g574(.A1(new_n756), .A2(new_n695), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G116), .ZN(G18));
  NAND2_X1  g576(.A1(new_n731), .A2(new_n654), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n754), .A2(new_n481), .A3(new_n525), .A4(new_n522), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n309), .A2(new_n765), .A3(new_n314), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  OAI21_X1  g581(.A(new_n251), .B1(new_n245), .B2(KEYINPUT106), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n240), .A2(KEYINPUT106), .A3(new_n244), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n303), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n299), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n748), .A2(new_n660), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n481), .A2(new_n589), .A3(new_n682), .A4(new_n645), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n755), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G122), .ZN(G24));
  NAND3_X1  g590(.A1(new_n731), .A2(new_n660), .A3(new_n771), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n589), .A2(new_n680), .A3(new_n715), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n589), .A2(new_n680), .A3(KEYINPUT107), .A4(new_n715), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n777), .A2(new_n782), .A3(new_n764), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n320), .ZN(G27));
  NAND3_X1  g598(.A1(new_n479), .A2(new_n394), .A3(new_n480), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT108), .ZN(new_n786));
  INV_X1    g600(.A(new_n525), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n522), .B2(new_n512), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n479), .A2(new_n789), .A3(new_n394), .A4(new_n480), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n782), .A3(KEYINPUT42), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n309), .A3(new_n314), .A4(new_n393), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n786), .A2(new_n788), .A3(new_n790), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n780), .A2(new_n781), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n308), .A2(new_n794), .A3(new_n795), .A4(new_n748), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT42), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(G131), .Z(G33));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n692), .A2(new_n800), .A3(new_n693), .A4(new_n715), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n716), .A2(KEYINPUT109), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n791), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n309), .A2(new_n804), .A3(new_n314), .A4(new_n393), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NAND2_X1  g620(.A1(new_n511), .A2(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT110), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n511), .A2(new_n809), .A3(KEYINPUT45), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(G469), .B1(new_n511), .B2(KEYINPUT45), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n516), .A2(new_n317), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(KEYINPUT46), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT46), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n812), .B1(new_n808), .B2(new_n810), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n818), .B1(new_n819), .B2(new_n815), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n820), .A3(new_n522), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n720), .A2(new_n525), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n823), .B(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n736), .A2(new_n680), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT43), .B1(new_n828), .B2(KEYINPUT113), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n661), .A3(KEYINPUT44), .A4(new_n731), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n786), .A2(new_n790), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n661), .A3(new_n731), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT44), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n827), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G137), .ZN(G39));
  NOR2_X1   g652(.A1(new_n744), .A2(new_n745), .ZN(new_n839));
  INV_X1    g653(.A(new_n833), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n750), .A2(new_n739), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n821), .A2(new_n525), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT47), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT47), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n821), .A2(new_n845), .A3(new_n525), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  NOR3_X1   g662(.A1(new_n746), .A2(new_n395), .A3(new_n787), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT114), .ZN(new_n850));
  INV_X1    g664(.A(new_n728), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n754), .A2(new_n522), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT49), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n730), .A2(new_n736), .A3(new_n680), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n850), .A2(new_n851), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT115), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n706), .A2(new_n707), .B1(new_n772), .B2(new_n774), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n736), .A2(new_n645), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n681), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n683), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n662), .A2(new_n393), .A3(new_n664), .A4(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n656), .A2(new_n857), .A3(new_n766), .A4(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n793), .A2(new_n797), .A3(new_n805), .ZN(new_n863));
  INV_X1    g677(.A(new_n755), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n751), .B(new_n864), .C1(new_n695), .C2(new_n757), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n568), .A2(new_n715), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n645), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n525), .A2(new_n523), .A3(new_n692), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n309), .A2(new_n314), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n795), .A2(new_n660), .A3(new_n771), .A4(new_n788), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n390), .A2(new_n704), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n833), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n862), .A2(new_n863), .A3(new_n865), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n777), .ZN(new_n876));
  INV_X1    g690(.A(new_n764), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n795), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n718), .A2(new_n742), .A3(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n481), .A2(new_n788), .A3(new_n589), .A4(new_n645), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n872), .A2(KEYINPUT116), .A3(new_n715), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT116), .B1(new_n872), .B2(new_n715), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n880), .B(new_n728), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n879), .A2(KEYINPUT117), .A3(KEYINPUT52), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n783), .B1(new_n839), .B2(new_n717), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n742), .A4(new_n883), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n718), .A2(new_n742), .A3(new_n878), .A4(new_n883), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n884), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n887), .B(KEYINPUT52), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n862), .A2(new_n863), .A3(new_n865), .A4(new_n874), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n894), .A2(new_n895), .A3(new_n893), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n875), .A2(new_n884), .A3(new_n891), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n893), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT51), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n833), .A2(new_n755), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n904), .A2(new_n648), .A3(new_n831), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n876), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n851), .A2(new_n393), .A3(new_n648), .A4(new_n904), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n736), .A2(new_n737), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n772), .A2(new_n648), .A3(new_n831), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n730), .A2(new_n864), .A3(new_n395), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(KEYINPUT50), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT50), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  OAI221_X1 g726(.A(new_n906), .B1(new_n907), .B2(new_n908), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n840), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n844), .A2(new_n846), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n852), .A2(new_n787), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n903), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(KEYINPUT118), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(KEYINPUT118), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n361), .A2(G952), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n909), .B2(new_n877), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT48), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n746), .B1(new_n312), .B2(new_n279), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n905), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n905), .B2(new_n924), .ZN(new_n926));
  OAI221_X1 g740(.A(new_n922), .B1(new_n681), .B2(new_n907), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n913), .A2(new_n917), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(KEYINPUT51), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n919), .A2(new_n920), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n902), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(G952), .A2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n856), .B1(new_n931), .B2(new_n932), .ZN(G75));
  AOI21_X1  g747(.A(new_n317), .B1(new_n892), .B2(new_n896), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G210), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n438), .A2(new_n446), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n444), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n935), .B2(new_n936), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n361), .A2(G952), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(G51));
  INV_X1    g757(.A(new_n898), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n897), .B1(new_n892), .B2(new_n896), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n815), .B(KEYINPUT119), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT57), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n946), .A2(new_n948), .B1(new_n521), .B2(new_n520), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n814), .B(KEYINPUT120), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n934), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n934), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n942), .B1(new_n949), .B2(new_n954), .ZN(G54));
  INV_X1    g769(.A(new_n942), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n957));
  INV_X1    g771(.A(new_n583), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n957), .A2(KEYINPUT122), .A3(new_n958), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G60));
  NAND3_X1  g778(.A1(new_n669), .A2(new_n673), .A3(new_n674), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT59), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n902), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n956), .B1(new_n946), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n891), .A2(new_n884), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n793), .A2(new_n797), .A3(new_n805), .ZN(new_n977));
  INV_X1    g791(.A(new_n873), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n869), .B2(new_n870), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n980), .A2(KEYINPUT53), .A3(new_n862), .A4(new_n865), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n886), .A2(new_n889), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT53), .B1(new_n875), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n975), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n381), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n942), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n974), .B1(new_n892), .B2(new_n896), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n702), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n987), .A2(KEYINPUT123), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n956), .B1(new_n989), .B2(new_n381), .ZN(new_n994));
  INV_X1    g808(.A(new_n702), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n995), .B(new_n974), .C1(new_n892), .C2(new_n896), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n992), .B(new_n993), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n991), .A2(new_n997), .ZN(G66));
  INV_X1    g812(.A(G224), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n652), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n862), .A2(new_n865), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n937), .B1(G898), .B2(new_n361), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT124), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G69));
  OAI21_X1  g820(.A(new_n255), .B1(new_n270), .B2(KEYINPUT30), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n574), .A2(new_n578), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n977), .B(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n481), .A2(new_n589), .A3(new_n645), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n836), .A2(new_n832), .B1(new_n924), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n847), .B(new_n879), .C1(new_n826), .C2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n361), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n711), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1016), .A2(KEYINPUT126), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(KEYINPUT126), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1009), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n361), .B1(G227), .B2(G900), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1009), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n734), .A2(new_n879), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT62), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  OR4_X1    g841(.A1(new_n752), .A2(new_n721), .A3(new_n833), .A4(new_n859), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1027), .A2(new_n837), .A3(new_n847), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n361), .A3(new_n1022), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1020), .A2(new_n1024), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1024), .B1(new_n1020), .B2(new_n1030), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1031), .A2(new_n1032), .ZN(G72));
  NAND2_X1  g847(.A1(G472), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT63), .Z(new_n1035));
  OAI21_X1  g849(.A(new_n1035), .B1(new_n1029), .B2(new_n1001), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n725), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n1011), .A2(new_n1015), .A3(new_n1001), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1035), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n724), .B(new_n251), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1037), .A2(new_n956), .A3(new_n1040), .ZN(new_n1041));
  AOI211_X1 g855(.A(new_n1039), .B(new_n901), .C1(new_n280), .C2(new_n273), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1041), .A2(new_n1042), .ZN(G57));
endmodule


