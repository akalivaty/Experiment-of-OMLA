//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT67), .ZN(G160));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(new_n458), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  MUX2_X1   g051(.A(G100), .B(G112), .S(G2105), .Z(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  OAI211_X1 g055(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g057(.A(G138), .B(new_n458), .C1(new_n470), .C2(new_n471), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n461), .A2(new_n485), .A3(G138), .A4(new_n458), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n458), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n489), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n489), .A2(new_n490), .A3(new_n493), .A4(KEYINPUT69), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n487), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(G543), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT5), .B(G543), .Z(new_n510));
  NOR2_X1   g085(.A1(new_n505), .A2(new_n506), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n501), .B(KEYINPUT70), .C1(new_n506), .C2(new_n505), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n508), .B1(new_n514), .B2(G88), .ZN(G166));
  AND2_X1   g090(.A1(new_n501), .A2(G63), .ZN(new_n516));
  AND3_X1   g091(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n507), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT71), .B(G51), .Z(new_n520));
  INV_X1    g095(.A(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n514), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  NAND2_X1  g102(.A1(new_n514), .A2(G90), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n510), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G651), .B1(new_n519), .B2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND3_X1  g109(.A1(new_n512), .A2(G81), .A3(new_n513), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n519), .A2(G43), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n510), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT72), .B1(new_n541), .B2(G651), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n501), .A2(G56), .ZN(new_n544));
  AOI211_X1 g119(.A(new_n543), .B(new_n503), .C1(new_n544), .C2(new_n539), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n537), .B(new_n538), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n536), .B(new_n535), .C1(new_n542), .C2(new_n545), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n519), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n514), .A2(G91), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n501), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT74), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(G299));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND2_X1  g139(.A1(new_n514), .A2(G87), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n501), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n519), .B2(G49), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n514), .A2(G86), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n510), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n519), .B2(G48), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n569), .A2(new_n573), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n503), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n519), .A2(G47), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT77), .B(G85), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n514), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n501), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G54), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n503), .B1(new_n591), .B2(new_n507), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT78), .Z(new_n593));
  NAND3_X1  g168(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n512), .A2(new_n513), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n589), .B1(new_n600), .B2(new_n588), .ZN(G284));
  AOI21_X1  g176(.A(new_n589), .B1(new_n600), .B2(new_n588), .ZN(G321));
  MUX2_X1   g177(.A(G286), .B(G299), .S(new_n588), .Z(G297));
  MUX2_X1   g178(.A(G286), .B(G299), .S(new_n588), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n600), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND3_X1  g181(.A1(new_n600), .A2(new_n605), .A3(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n549), .A2(new_n588), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT11), .Z(G282));
  INV_X1    g185(.A(new_n609), .ZN(G323));
  NAND2_X1  g186(.A1(new_n473), .A2(G2104), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT79), .B(G2100), .Z(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  MUX2_X1   g192(.A(G99), .B(G111), .S(G2105), .Z(new_n618));
  AOI22_X1  g193(.A1(new_n475), .A2(G123), .B1(G2104), .B2(new_n618), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n473), .A2(KEYINPUT80), .A3(G135), .ZN(new_n620));
  AOI21_X1  g195(.A(KEYINPUT80), .B1(new_n473), .B2(G135), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT81), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n628), .B2(new_n630), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n632), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT82), .Z(new_n640));
  INV_X1    g215(.A(G14), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT18), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n649), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(KEYINPUT17), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(KEYINPUT17), .A3(new_n648), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n648), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n655), .B1(new_n646), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n651), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  INV_X1    g246(.A(new_n666), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G29), .A2(G32), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n458), .A2(G105), .A3(G2104), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT94), .Z(new_n687));
  INV_X1    g262(.A(G141), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n462), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n475), .A2(G129), .ZN(new_n690));
  NAND3_X1  g265(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT26), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n685), .B1(new_n696), .B2(G29), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT27), .B(G1996), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G27), .A2(G29), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G164), .B2(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G2078), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(G160), .A2(G29), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  AND2_X1   g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  NOR2_X1   g282(.A1(KEYINPUT24), .A2(G34), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n705), .A2(G2084), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(G2084), .B1(new_n705), .B2(new_n709), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G2078), .B2(new_n702), .ZN(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  OR2_X1    g288(.A1(G29), .A2(G35), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n479), .B2(new_n706), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT29), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n697), .A2(new_n699), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n704), .A2(new_n710), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n706), .A2(G33), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n459), .A2(G103), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G139), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n462), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n458), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n719), .B1(new_n727), .B2(new_n706), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2072), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G21), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G286), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n729), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n730), .A2(G5), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G301), .B2(G16), .ZN(new_n738));
  INV_X1    g313(.A(G1961), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n716), .A2(new_n713), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n738), .A2(new_n739), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT30), .B(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n706), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n622), .B2(new_n706), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n743), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G299), .A2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n730), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G1956), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n736), .A2(new_n742), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n718), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n706), .A2(G26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n473), .A2(G140), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n475), .A2(G128), .ZN(new_n761));
  MUX2_X1   g336(.A(G104), .B(G116), .S(G2105), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2104), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n706), .ZN(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n600), .B2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n769), .B1(G1348), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(G1348), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n730), .A2(G19), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n546), .A2(new_n548), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1341), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n774), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n757), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n774), .B2(new_n779), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT97), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n784), .A2(new_n785), .A3(new_n780), .A4(new_n757), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G6), .A2(G16), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  OAI211_X1 g365(.A(new_n789), .B(new_n790), .C1(G305), .C2(new_n730), .ZN(new_n791));
  INV_X1    g366(.A(new_n790), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n730), .B1(new_n576), .B2(new_n578), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n788), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n730), .A2(G23), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G288), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT89), .B1(new_n800), .B2(G16), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n800), .A2(KEYINPUT89), .A3(G16), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n801), .B(new_n802), .C1(G166), .C2(new_n730), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1971), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n807));
  NOR2_X1   g382(.A1(G25), .A2(G29), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n473), .A2(G131), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n475), .A2(G119), .ZN(new_n810));
  OAI21_X1  g385(.A(KEYINPUT87), .B1(G95), .B2(G2105), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR3_X1   g387(.A1(KEYINPUT87), .A2(G95), .A3(G2105), .ZN(new_n813));
  OAI221_X1 g388(.A(G2104), .B1(G107), .B2(new_n458), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n809), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n808), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XOR2_X1   g392(.A(new_n816), .B(new_n817), .Z(new_n818));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n819));
  NAND2_X1  g394(.A1(G290), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n583), .A2(KEYINPUT88), .A3(new_n584), .A4(new_n586), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n730), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G1986), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n730), .A2(G24), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n823), .B1(new_n822), .B2(new_n825), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n818), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n795), .A2(new_n829), .A3(new_n805), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT90), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n828), .B2(new_n830), .ZN(new_n833));
  OAI211_X1 g408(.A(KEYINPUT91), .B(new_n807), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n828), .A2(new_n830), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT90), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT91), .B1(new_n839), .B2(new_n807), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n787), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n835), .A2(new_n840), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(G311));
  OR2_X1    g418(.A1(new_n835), .A2(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n835), .A2(new_n840), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(KEYINPUT98), .A3(new_n845), .A4(new_n787), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n841), .B2(new_n842), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(G150));
  AOI22_X1  g424(.A1(new_n514), .A2(G93), .B1(G55), .B2(new_n519), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n510), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n503), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n593), .A2(new_n599), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n605), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n549), .A2(new_n857), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n547), .A2(new_n850), .A3(new_n856), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n862), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n869), .B(new_n870), .C1(new_n867), .C2(new_n866), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n859), .B1(new_n871), .B2(new_n872), .ZN(G145));
  XOR2_X1   g448(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n874));
  MUX2_X1   g449(.A(G106), .B(G118), .S(G2105), .Z(new_n875));
  AOI22_X1  g450(.A1(new_n475), .A2(G130), .B1(G2104), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n462), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n613), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n694), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n764), .B(KEYINPUT92), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G164), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n766), .A2(new_n499), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n727), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n883), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT101), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n694), .A3(new_n886), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n696), .A2(new_n883), .A3(new_n884), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n696), .B1(new_n883), .B2(new_n884), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n727), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n815), .B(KEYINPUT102), .Z(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n894), .B2(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n880), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n894), .A2(new_n897), .ZN(new_n903));
  INV_X1    g478(.A(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n879), .A3(new_n899), .ZN(new_n906));
  XNOR2_X1  g481(.A(G160), .B(new_n479), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n622), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n908), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n900), .A2(new_n901), .A3(new_n880), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n879), .B1(new_n905), .B2(new_n899), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT103), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(new_n912), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  AOI211_X1 g493(.A(new_n874), .B(new_n911), .C1(new_n916), .C2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n874), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(new_n911), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n919), .A2(new_n923), .ZN(G395));
  NOR2_X1   g499(.A1(new_n857), .A2(G868), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n600), .A2(KEYINPUT105), .A3(G299), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT105), .B1(new_n600), .B2(G299), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n600), .A2(G299), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT41), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n926), .A2(new_n931), .A3(new_n927), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n600), .A2(new_n605), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n865), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n929), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(G305), .B(G303), .ZN(new_n943));
  XNOR2_X1  g518(.A(G290), .B(G288), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n942), .B(new_n946), .Z(new_n947));
  AOI21_X1  g522(.A(new_n925), .B1(new_n947), .B2(G868), .ZN(G295));
  AOI21_X1  g523(.A(new_n925), .B1(new_n947), .B2(G868), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g525(.A1(G171), .A2(KEYINPUT107), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(G286), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  AOI21_X1  g528(.A(G168), .B1(new_n953), .B2(G301), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(new_n865), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n865), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n929), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n930), .B(new_n932), .C1(new_n957), .C2(new_n956), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n945), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n910), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n945), .B1(new_n959), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n960), .ZN(new_n965));
  INV_X1    g540(.A(new_n945), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n910), .A4(new_n961), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n968), .B2(KEYINPUT108), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n964), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n964), .B2(new_n969), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n950), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n964), .A2(new_n969), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n970), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n964), .A2(new_n969), .A3(new_n971), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(G397));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n499), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n467), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n473), .A2(G137), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n984), .A2(G40), .A3(new_n460), .A4(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n882), .A2(G2067), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n766), .A2(new_n768), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n987), .B1(new_n991), .B2(new_n881), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n987), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n996), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n992), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n696), .A2(new_n994), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n990), .B(new_n1000), .C1(new_n994), .C2(new_n694), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n815), .A2(new_n817), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n989), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n987), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(KEYINPUT48), .A3(new_n987), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT48), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1005), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(new_n1008), .B2(new_n996), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n815), .B(new_n817), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1006), .B(new_n1009), .C1(new_n1011), .C2(new_n996), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n999), .A2(new_n1004), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1384), .B1(new_n487), .B2(new_n498), .ZN(new_n1014));
  INV_X1    g589(.A(G40), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n464), .A2(new_n467), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G8), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n577), .B(G1981), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT49), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(G8), .A3(new_n1017), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  INV_X1    g597(.A(G288), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n577), .A2(G1981), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1018), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1016), .B1(new_n1014), .B2(KEYINPUT45), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n982), .B(G1384), .C1(new_n487), .C2(new_n498), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(G1971), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(KEYINPUT110), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1016), .B1(new_n1014), .B2(new_n1033), .ZN(new_n1034));
  AOI211_X1 g609(.A(KEYINPUT50), .B(G1384), .C1(new_n487), .C2(new_n498), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1031), .A2(KEYINPUT110), .B1(new_n713), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1027), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G303), .A2(G8), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT55), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1018), .B1(G1976), .B2(new_n1023), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(new_n1045), .C1(G1976), .C2(new_n1023), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1021), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1026), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1042), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1014), .A2(new_n1033), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT111), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n986), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1035), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1031), .B1(new_n1056), .B2(G2090), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1041), .B1(new_n1057), .B2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT113), .B1(new_n1036), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1034), .A2(new_n1035), .A3(new_n1062), .A4(G2084), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1014), .A2(KEYINPUT45), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n983), .A2(new_n1065), .A3(new_n1016), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(KEYINPUT112), .A3(new_n733), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n733), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1027), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G168), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT63), .B1(new_n1059), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(KEYINPUT63), .C1(new_n1041), .C2(new_n1038), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n1050), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1049), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1053), .A2(new_n1060), .A3(new_n1051), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1062), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1036), .A2(KEYINPUT113), .A3(new_n1060), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1079), .A2(new_n1083), .A3(KEYINPUT117), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G168), .A2(new_n1027), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n986), .B1(new_n981), .B2(new_n982), .ZN(new_n1092));
  INV_X1    g667(.A(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(KEYINPUT53), .A3(new_n1093), .A4(new_n1065), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n739), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(KEYINPUT122), .A3(new_n1095), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1066), .B2(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT117), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1064), .A2(new_n1085), .A3(new_n1071), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1027), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1088), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT119), .B1(new_n1087), .B2(new_n1027), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1110), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1072), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1088), .A2(KEYINPUT51), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1118), .A2(KEYINPUT120), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT120), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1091), .B(new_n1109), .C1(new_n1117), .C2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1107), .A2(KEYINPUT62), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1056), .A2(new_n754), .B1(new_n1030), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n557), .B2(KEYINPUT114), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(G299), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(KEYINPUT116), .A2(KEYINPUT61), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1017), .A2(G2067), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1053), .A2(new_n1051), .ZN(new_n1132));
  INV_X1    g707(.A(G1348), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n860), .A2(KEYINPUT60), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1130), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1092), .A2(new_n994), .A3(new_n1065), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1017), .A2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n777), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n549), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1136), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1134), .A2(new_n860), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1036), .A2(G1348), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n600), .B1(new_n1147), .B2(new_n1131), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1145), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1129), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1131), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1128), .A2(new_n1126), .B1(new_n1154), .B2(new_n600), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n860), .A4(new_n1153), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT115), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(KEYINPUT116), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(KEYINPUT116), .B2(new_n1160), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1157), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1151), .B(new_n1155), .C1(new_n1156), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1150), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1100), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1030), .B2(new_n1093), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT126), .B1(new_n1096), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1101), .A2(new_n1170), .A3(new_n1095), .A4(new_n1094), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1166), .B1(new_n1172), .B2(G171), .ZN(new_n1173));
  AOI211_X1 g748(.A(KEYINPUT127), .B(G301), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1098), .A2(G301), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT125), .Z(new_n1178));
  AOI21_X1  g753(.A(new_n1165), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1101), .A2(new_n1095), .A3(new_n1094), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1105), .B(new_n1106), .C1(G171), .C2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1124), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1110), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1114), .B(G8), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1089), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1185), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1090), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1123), .B1(new_n1184), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1078), .B1(new_n1192), .B2(new_n1059), .ZN(new_n1193));
  XNOR2_X1  g768(.A(G290), .B(new_n823), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n996), .B1(new_n1011), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1013), .B1(new_n1193), .B2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g771(.A1(new_n921), .A2(new_n922), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n643), .A2(G319), .ZN(new_n1199));
  NOR3_X1   g773(.A1(new_n1199), .A2(G227), .A3(G229), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1198), .A2(new_n975), .A3(new_n1200), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


