//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n227), .B(new_n230), .ZN(G358));
  XOR2_X1   g0031(.A(G107), .B(G116), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G87), .B(G97), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G351));
  AND2_X1   g0040(.A1(G33), .A2(G41), .ZN(new_n241));
  OAI21_X1  g0041(.A(KEYINPUT66), .B1(new_n241), .B2(new_n211), .ZN(new_n242));
  INV_X1    g0042(.A(G1), .ZN(new_n243));
  OAI21_X1  g0043(.A(new_n243), .B1(G41), .B2(G45), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT66), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n246), .A2(new_n247), .A3(G1), .A4(G13), .ZN(new_n248));
  NAND4_X1  g0048(.A1(new_n242), .A2(new_n245), .A3(G274), .A4(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(G223), .B1(new_n259), .B2(G77), .ZN(new_n260));
  INV_X1    g0060(.A(G222), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(new_n255), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n241), .A2(new_n211), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n250), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n242), .A2(new_n248), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT67), .B1(new_n267), .B2(new_n245), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT67), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n242), .A2(new_n269), .A3(new_n244), .A4(new_n248), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G226), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G50), .ZN(new_n276));
  INV_X1    g0076(.A(G58), .ZN(new_n277));
  INV_X1    g0077(.A(G68), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n279), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT69), .B1(new_n253), .B2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n212), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n211), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n291), .A3(new_n211), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n276), .B1(new_n243), .B2(G20), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n290), .A2(new_n297), .A3(new_n292), .A4(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n295), .A2(new_n212), .A3(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n276), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n299), .B2(new_n302), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n294), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n266), .A2(new_n306), .A3(new_n272), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n275), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  XOR2_X1   g0109(.A(new_n305), .B(KEYINPUT9), .Z(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n273), .A2(G200), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(KEYINPUT73), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n313), .B1(new_n316), .B2(new_n273), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n311), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n314), .B1(new_n310), .B2(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n309), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n256), .A2(G238), .B1(new_n259), .B2(G107), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n259), .A2(G1698), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(G232), .ZN(new_n325));
  INV_X1    g0125(.A(G232), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n263), .A2(KEYINPUT71), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n322), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n265), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n250), .B1(new_n271), .B2(G244), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(new_n306), .ZN(new_n331));
  INV_X1    g0131(.A(new_n289), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT72), .B1(new_n332), .B2(new_n297), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n301), .A2(new_n289), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n243), .A2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G77), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n301), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n286), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT15), .B(G87), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n285), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n289), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n339), .A2(new_n341), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n329), .A2(new_n330), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n331), .B(new_n347), .C1(new_n348), .C2(G169), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n339), .A2(new_n341), .A3(new_n346), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n329), .A2(new_n330), .A3(G190), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(new_n351), .C1(new_n348), .C2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n321), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n301), .A2(new_n278), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n278), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n285), .B2(new_n340), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT11), .B1(new_n358), .B2(new_n293), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n337), .A2(G68), .A3(new_n338), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n271), .A2(G238), .ZN(new_n366));
  OAI211_X1 g0166(.A(G232), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n367));
  OAI211_X1 g0167(.A(G226), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n250), .B1(new_n265), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT13), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G238), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n268), .B2(new_n270), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n370), .A2(new_n265), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n249), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT13), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n373), .A2(new_n378), .A3(G190), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n365), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n352), .B1(new_n373), .B2(new_n378), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT75), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n372), .B1(new_n366), .B2(new_n371), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n375), .A2(new_n377), .A3(KEYINPUT13), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n383), .B(G169), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n373), .A2(new_n378), .A3(G179), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT74), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n274), .B1(new_n373), .B2(new_n378), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n383), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n390), .B2(new_n389), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n387), .B(new_n388), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n382), .B1(new_n394), .B2(new_n364), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n242), .A2(G232), .A3(new_n244), .A4(new_n248), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n249), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT78), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT78), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n249), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT77), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(KEYINPUT77), .A2(G33), .A3(G87), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(G223), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(G179), .B1(new_n409), .B2(new_n265), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n399), .A2(new_n401), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n265), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n404), .A2(new_n405), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n256), .B2(G226), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n412), .B1(new_n414), .B2(new_n407), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n274), .B1(new_n415), .B2(new_n398), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n293), .A2(new_n301), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n286), .B1(new_n243), .B2(G20), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n418), .A2(new_n419), .B1(new_n301), .B2(new_n286), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n277), .A2(new_n278), .ZN(new_n421));
  NOR2_X1   g0221(.A1(G58), .A2(G68), .ZN(new_n422));
  OAI21_X1  g0222(.A(G20), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n280), .A2(G159), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n257), .A2(new_n258), .A3(new_n427), .A4(G20), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT76), .B1(new_n257), .B2(new_n258), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n254), .A2(new_n430), .A3(new_n255), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n431), .A3(new_n212), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n428), .B1(new_n432), .B2(new_n427), .ZN(new_n433));
  OAI211_X1 g0233(.A(KEYINPUT16), .B(new_n426), .C1(new_n433), .C2(new_n278), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT16), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n254), .A2(new_n212), .A3(new_n255), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n427), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n278), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n439), .B2(new_n425), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n434), .A2(new_n289), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n417), .B1(new_n420), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  INV_X1    g0244(.A(new_n420), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT7), .B1(new_n259), .B2(new_n212), .ZN(new_n446));
  OAI21_X1  g0246(.A(G68), .B1(new_n446), .B2(new_n428), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n426), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n332), .B1(new_n448), .B2(new_n435), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n445), .B1(new_n449), .B2(new_n434), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n444), .B1(new_n450), .B2(new_n417), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT79), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n443), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n434), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n440), .A2(new_n289), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n420), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n417), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(KEYINPUT79), .A3(new_n444), .ZN(new_n459));
  AND2_X1   g0259(.A1(KEYINPUT80), .A2(G190), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT80), .A2(G190), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n409), .B2(new_n265), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n399), .A2(new_n401), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n352), .B1(new_n415), .B2(new_n398), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n441), .A2(new_n466), .A3(new_n420), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(KEYINPUT17), .A3(new_n466), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n469), .A2(KEYINPUT81), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT81), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n453), .B(new_n459), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n354), .A2(new_n396), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n297), .A2(G97), .ZN(new_n475));
  OAI21_X1  g0275(.A(G107), .B1(new_n446), .B2(new_n428), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT6), .ZN(new_n477));
  AND2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n202), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n475), .B1(new_n484), .B2(new_n289), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n243), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n290), .A2(new_n297), .A3(new_n292), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT82), .B1(new_n492), .B2(G41), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  INV_X1    g0294(.A(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT5), .ZN(new_n496));
  INV_X1    g0296(.A(G45), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n492), .A2(G41), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n493), .A2(new_n496), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(G257), .A3(new_n242), .A4(new_n248), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n242), .A2(G274), .A3(new_n248), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n500), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G244), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n256), .A2(G250), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n265), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n504), .A2(G179), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n274), .B1(new_n504), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n491), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI211_X1 g0315(.A(new_n489), .B(new_n475), .C1(new_n484), .C2(new_n289), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n511), .A2(new_n265), .ZN(new_n517));
  OAI21_X1  g0317(.A(G200), .B1(new_n517), .B2(new_n503), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n504), .A2(G190), .A3(new_n512), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT25), .ZN(new_n522));
  AOI21_X1  g0322(.A(G107), .B1(new_n522), .B2(KEYINPUT91), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n301), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n487), .A2(new_n480), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(G20), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT89), .B1(new_n212), .B2(G107), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT23), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT89), .B(new_n534), .C1(new_n212), .C2(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n212), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n537), .A2(KEYINPUT22), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(KEYINPUT22), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(KEYINPUT24), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n537), .B(KEYINPUT22), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n536), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n289), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT90), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n540), .A2(KEYINPUT24), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n542), .A3(new_n536), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n289), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n529), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G250), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n554), .C1(new_n253), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n265), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n242), .A2(G274), .A3(new_n248), .ZN(new_n558));
  AND4_X1   g0358(.A1(new_n496), .A2(new_n493), .A3(new_n498), .A4(new_n499), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n500), .A2(G264), .A3(new_n242), .A4(new_n248), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n352), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT93), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(new_n561), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(KEYINPUT92), .A3(new_n316), .A4(new_n560), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT92), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n562), .B2(G190), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(KEYINPUT93), .A3(new_n352), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n565), .A2(new_n568), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n521), .B1(new_n552), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n262), .A2(new_n212), .A3(G68), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT85), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n285), .B2(new_n488), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n212), .B1(new_n369), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(G87), .B2(new_n203), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n262), .A2(KEYINPUT85), .A3(new_n212), .A4(G68), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n576), .A2(new_n578), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n289), .B1(new_n301), .B2(new_n344), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  OR3_X1    g0384(.A1(new_n487), .A2(new_n584), .A3(new_n344), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n487), .B2(new_n344), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT87), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n583), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n592));
  OAI211_X1 g0392(.A(G238), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n530), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n265), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT83), .B1(new_n497), .B2(G1), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT83), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n243), .A3(G45), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n598), .A3(G250), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT84), .B1(new_n267), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n596), .A2(new_n598), .A3(G250), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n242), .A4(new_n248), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n242), .A2(G274), .A3(new_n248), .A4(new_n498), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n595), .A2(new_n600), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n605), .A2(G179), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n274), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n589), .A2(new_n591), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G87), .ZN(new_n609));
  OR3_X1    g0409(.A1(new_n487), .A2(KEYINPUT88), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT88), .B1(new_n487), .B2(new_n609), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n583), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n605), .A2(new_n316), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n605), .A2(G200), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  OAI211_X1 g0419(.A(G264), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n620));
  OAI211_X1 g0420(.A(G257), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n254), .A2(G303), .A3(new_n255), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n265), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n500), .A2(G270), .A3(new_n242), .A4(new_n248), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n560), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G169), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n486), .A2(G116), .ZN(new_n628));
  INV_X1    g0428(.A(new_n335), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n334), .B1(new_n301), .B2(new_n289), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G116), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n296), .A2(G20), .A3(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n288), .A2(new_n211), .B1(G20), .B2(new_n632), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n510), .B(new_n212), .C1(G33), .C2(new_n488), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT20), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n619), .B1(new_n627), .B2(new_n639), .ZN(new_n640));
  OAI221_X1 g0440(.A(new_n633), .B1(new_n637), .B2(new_n636), .C1(new_n336), .C2(new_n628), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(KEYINPUT21), .A3(new_n626), .A4(G169), .ZN(new_n642));
  AND4_X1   g0442(.A1(G179), .A2(new_n560), .A3(new_n624), .A4(new_n625), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n626), .A2(G200), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n560), .A2(new_n624), .A3(new_n462), .A4(new_n625), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n639), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n640), .A2(new_n642), .A3(new_n644), .A4(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n550), .B1(new_n549), .B2(new_n289), .ZN(new_n649));
  AOI211_X1 g0449(.A(KEYINPUT90), .B(new_n332), .C1(new_n547), .C2(new_n548), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n528), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n562), .A2(G179), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n274), .B2(new_n562), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n648), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n474), .A2(new_n573), .A3(new_n618), .A4(new_n654), .ZN(G372));
  AND2_X1   g0455(.A1(new_n443), .A2(new_n451), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n382), .ZN(new_n658));
  INV_X1    g0458(.A(new_n349), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n394), .A2(new_n364), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n472), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n469), .A2(KEYINPUT81), .A3(new_n470), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n657), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n319), .A2(new_n320), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n309), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n474), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n504), .A2(G179), .A3(new_n512), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n503), .B1(new_n265), .B2(new_n511), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n274), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT97), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n669), .B(new_n673), .C1(new_n670), .C2(new_n274), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n672), .A2(new_n491), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n594), .A2(KEYINPUT94), .A3(new_n265), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT94), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n595), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n588), .B(new_n606), .C1(new_n681), .C2(G169), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT95), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n680), .A2(new_n678), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n683), .B(G200), .C1(new_n684), .C2(new_n677), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT95), .B1(new_n681), .B2(new_n352), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n615), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n675), .A2(new_n676), .A3(new_n682), .A4(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n515), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n608), .A2(new_n689), .A3(new_n617), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n691), .A3(new_n682), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n640), .A2(new_n644), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n642), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n651), .B2(new_n653), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n546), .A2(new_n551), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n572), .A3(new_n528), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n515), .A2(new_n520), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n682), .A4(new_n687), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n695), .B1(new_n699), .B2(KEYINPUT96), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n687), .A2(new_n682), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT96), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n573), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n692), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n667), .B1(new_n668), .B2(new_n704), .ZN(G369));
  NAND2_X1  g0505(.A1(new_n651), .A2(new_n653), .ZN(new_n706));
  INV_X1    g0506(.A(new_n296), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n707), .A2(KEYINPUT27), .A3(G20), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT27), .B1(new_n707), .B2(G20), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G213), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G343), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n712), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n697), .B1(new_n552), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n713), .B1(new_n706), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n714), .A2(new_n639), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n694), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n648), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g0520(.A(KEYINPUT98), .B(G330), .Z(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n694), .A2(new_n714), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT99), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n713), .B1(new_n728), .B2(new_n716), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n729), .ZN(G399));
  INV_X1    g0530(.A(new_n206), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(G1), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n209), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n573), .A2(new_n618), .A3(new_n654), .A4(new_n714), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n605), .A2(new_n566), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n670), .A3(new_n643), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(KEYINPUT100), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n742), .B1(new_n741), .B2(KEYINPUT100), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n562), .A2(new_n626), .A3(new_n306), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n681), .A2(new_n745), .A3(new_n670), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n739), .B1(new_n747), .B2(new_n714), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n741), .A2(KEYINPUT100), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  INV_X1    g0550(.A(new_n746), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n741), .A2(KEYINPUT100), .A3(new_n742), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n738), .A2(new_n748), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n721), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  OAI211_X1 g0559(.A(KEYINPUT101), .B(new_n759), .C1(new_n704), .C2(new_n712), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n695), .A2(new_n699), .B1(KEYINPUT26), .B2(new_n690), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n687), .A2(new_n682), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n672), .A2(new_n491), .A3(new_n674), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT26), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n682), .ZN(new_n765));
  OAI211_X1 g0565(.A(KEYINPUT29), .B(new_n714), .C1(new_n761), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT101), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n706), .A2(new_n642), .A3(new_n693), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n703), .A3(new_n770), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n688), .A2(new_n682), .A3(new_n691), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n712), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n768), .B1(new_n773), .B2(KEYINPUT29), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n758), .B1(new_n767), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n737), .B1(new_n777), .B2(G1), .ZN(G364));
  INV_X1    g0578(.A(new_n723), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n295), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n243), .B1(new_n780), .B2(G45), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OR3_X1    g0582(.A1(new_n732), .A2(new_n782), .A3(KEYINPUT102), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT102), .B1(new_n732), .B2(new_n782), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n722), .B2(new_n720), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n211), .B1(G20), .B2(new_n274), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n212), .A2(new_n306), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n792), .A2(new_n352), .A3(G190), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n212), .A2(G179), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(new_n316), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n793), .A2(G68), .B1(G107), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n462), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n798), .A2(new_n352), .A3(new_n792), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n800), .B2(new_n276), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n791), .A2(new_n316), .A3(new_n352), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n802), .A2(KEYINPUT104), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(KEYINPUT104), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n801), .B1(G77), .B2(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n798), .A2(G200), .A3(new_n792), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n262), .B1(new_n809), .B2(new_n277), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G179), .A2(G200), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n212), .B1(new_n811), .B2(G190), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n488), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n794), .A2(G190), .A3(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n609), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n810), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n811), .A2(G20), .A3(new_n316), .ZN(new_n817));
  INV_X1    g0617(.A(G159), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT32), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n807), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n259), .B1(new_n814), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n802), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n823), .B(new_n825), .C1(new_n799), .C2(G326), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  INV_X1    g0627(.A(G329), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n795), .A2(new_n827), .B1(new_n828), .B2(new_n817), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT105), .Z(new_n830));
  INV_X1    g0630(.A(new_n812), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G294), .ZN(new_n832));
  XNOR2_X1  g0632(.A(KEYINPUT33), .B(G317), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n808), .A2(G322), .B1(new_n793), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n826), .A2(new_n830), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n790), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(G13), .A2(G33), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(G20), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n789), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n429), .A2(new_n431), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n731), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n497), .B2(new_n210), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n239), .B2(new_n497), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n262), .A2(new_n206), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT103), .Z(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G355), .B1(new_n632), .B2(new_n731), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n841), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n836), .A2(new_n850), .A3(new_n785), .ZN(new_n851));
  INV_X1    g0651(.A(new_n839), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n720), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n788), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NAND2_X1  g0655(.A1(new_n771), .A2(new_n772), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n347), .A2(new_n712), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n349), .A2(new_n353), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT107), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n349), .A2(new_n353), .A3(new_n860), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n856), .A2(new_n714), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n659), .A2(new_n712), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n859), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n773), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n786), .B1(new_n866), .B2(new_n758), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n758), .B2(new_n866), .ZN(new_n868));
  AOI22_X1  g0668(.A1(G137), .A2(new_n799), .B1(new_n808), .B2(G143), .ZN(new_n869));
  INV_X1    g0669(.A(G150), .ZN(new_n870));
  INV_X1    g0670(.A(new_n793), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .C1(new_n818), .C2(new_n805), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT34), .ZN(new_n873));
  INV_X1    g0673(.A(new_n842), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n796), .A2(G68), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n875), .B1(new_n276), .B2(new_n814), .C1(new_n277), .C2(new_n812), .ZN(new_n876));
  INV_X1    g0676(.A(new_n817), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n874), .B(new_n876), .C1(G132), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n871), .A2(KEYINPUT106), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n871), .A2(KEYINPUT106), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n883), .A2(G283), .B1(G116), .B2(new_n806), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n262), .B(new_n813), .C1(G311), .C2(new_n877), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n795), .A2(new_n609), .ZN(new_n886));
  INV_X1    g0686(.A(new_n814), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(G107), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(G294), .A2(new_n808), .B1(new_n799), .B2(G303), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n884), .A2(new_n885), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n790), .B1(new_n879), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n789), .A2(new_n837), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n785), .B(new_n891), .C1(new_n340), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n838), .B2(new_n865), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n868), .A2(new_n894), .ZN(G384));
  OR2_X1    g0695(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(G116), .A3(new_n213), .A4(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  OAI211_X1 g0699(.A(new_n210), .B(G77), .C1(new_n277), .C2(new_n278), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n276), .A2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n243), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n426), .B1(new_n433), .B2(new_n278), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n435), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n293), .A3(new_n434), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n906), .A2(new_n420), .B1(new_n417), .B2(new_n710), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n441), .A2(new_n466), .A3(new_n420), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n710), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n456), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n458), .A2(new_n911), .A3(new_n912), .A4(new_n467), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n906), .A2(new_n420), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n910), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n473), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n920), .B(new_n914), .C1(new_n473), .C2(new_n917), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT39), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n394), .A2(new_n364), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n712), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n908), .A2(new_n442), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT109), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n450), .B2(new_n710), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n927), .A2(new_n911), .B1(KEYINPUT37), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n458), .A2(new_n911), .A3(new_n467), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n710), .B1(new_n441), .B2(new_n420), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT37), .B1(new_n932), .B2(KEYINPUT109), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n469), .A2(new_n470), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n932), .B1(new_n656), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n926), .B1(new_n921), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n923), .A2(new_n925), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n365), .A2(new_n714), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n394), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT108), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n394), .A2(KEYINPUT108), .A3(new_n941), .ZN(new_n945));
  INV_X1    g0745(.A(new_n941), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n944), .A2(new_n945), .B1(new_n395), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n349), .A2(new_n712), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n947), .B1(new_n863), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n453), .A2(new_n459), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n916), .B1(new_n663), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n920), .B1(new_n952), .B2(new_n914), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n918), .A2(KEYINPUT38), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n656), .A2(new_n710), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n940), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n774), .A2(new_n760), .A3(new_n474), .A4(new_n766), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(new_n667), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n958), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n755), .A2(new_n865), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT110), .B1(new_n947), .B2(new_n962), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n859), .A2(new_n864), .A3(new_n861), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n746), .B1(new_n749), .B2(KEYINPUT30), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n739), .B(new_n714), .C1(new_n965), .C2(new_n752), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT31), .B1(new_n753), .B2(new_n712), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n964), .B1(new_n968), .B2(new_n738), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n924), .A2(new_n658), .A3(new_n946), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT108), .B1(new_n394), .B2(new_n941), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n394), .A2(KEYINPUT108), .A3(new_n941), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT40), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT110), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n969), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n963), .A2(new_n976), .A3(new_n955), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n969), .A2(new_n973), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n938), .B1(KEYINPUT38), .B2(new_n918), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT40), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n668), .A2(new_n756), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n721), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n961), .A2(new_n984), .B1(new_n243), .B2(new_n780), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n961), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n903), .B1(new_n985), .B2(new_n986), .ZN(G367));
  OAI221_X1 g0787(.A(new_n840), .B1(new_n206), .B2(new_n344), .C1(new_n844), .C2(new_n230), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(new_n786), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n613), .A2(new_n712), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n701), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n682), .B2(new_n990), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n809), .A2(new_n870), .B1(new_n278), .B2(new_n812), .ZN(new_n993));
  INV_X1    g0793(.A(G143), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n800), .A2(new_n994), .B1(new_n340), .B2(new_n795), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n259), .B1(new_n877), .B2(G137), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n277), .B2(new_n814), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n993), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n276), .B2(new_n805), .C1(new_n818), .C2(new_n882), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n795), .A2(new_n488), .B1(new_n812), .B2(new_n480), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n822), .A2(new_n809), .B1(new_n800), .B2(new_n824), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G283), .C2(new_n806), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n555), .B2(new_n882), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n842), .B1(G317), .B2(new_n877), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n887), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT46), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n814), .B2(new_n632), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n999), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT47), .Z(new_n1010));
  OAI221_X1 g0810(.A(new_n989), .B1(new_n852), .B2(new_n992), .C1(new_n1010), .C2(new_n790), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n675), .A2(new_n712), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n698), .B1(new_n516), .B2(new_n714), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n729), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT44), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n729), .A2(new_n1018), .A3(new_n1014), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n729), .B2(new_n1014), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n725), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1017), .A2(new_n725), .A3(new_n1021), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n728), .B(new_n716), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT113), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n723), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n723), .B(new_n1027), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n777), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n732), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n782), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n728), .A2(new_n716), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1014), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n1037), .A2(KEYINPUT42), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT42), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1014), .B(KEYINPUT111), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n706), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n689), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1039), .B(new_n1040), .C1(new_n1043), .C2(new_n712), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n724), .A2(new_n1041), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT112), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1050), .A2(new_n1051), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1051), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n1054), .A3(new_n1049), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1011), .B1(new_n1036), .B2(new_n1056), .ZN(G387));
  NAND2_X1  g0857(.A1(new_n777), .A2(new_n1031), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1032), .A2(new_n776), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n732), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n799), .A2(G159), .B1(G97), .B2(new_n796), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n808), .A2(G50), .B1(G77), .B2(new_n887), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n802), .A2(new_n278), .B1(new_n812), .B2(new_n344), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n342), .B2(new_n793), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n874), .B1(G150), .B2(new_n877), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n842), .B1(G326), .B2(new_n877), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G317), .A2(new_n808), .B1(new_n799), .B2(G322), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n822), .B2(new_n805), .C1(new_n882), .C2(new_n824), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n887), .A2(G294), .B1(new_n831), .B2(G283), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1067), .B1(new_n632), .B2(new_n795), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1066), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n789), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n734), .B(new_n497), .C1(new_n278), .C2(new_n340), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(KEYINPUT114), .ZN(new_n1082));
  OR3_X1    g0882(.A1(new_n286), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT50), .B1(new_n286), .B2(G50), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT114), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1084), .C1(new_n1080), .C2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n843), .B1(new_n1082), .B2(new_n1086), .C1(new_n227), .C2(new_n497), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n848), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1087), .B1(G107), .B2(new_n206), .C1(new_n734), .C2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n785), .B1(new_n1089), .B2(new_n840), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1079), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n717), .B2(new_n839), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1031), .B2(new_n782), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1060), .A2(new_n1093), .ZN(G393));
  INV_X1    g0894(.A(new_n1024), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n1022), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n782), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n235), .A2(new_n844), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n841), .B1(G97), .B2(new_n731), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n785), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G311), .A2(new_n808), .B1(new_n799), .B2(G317), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  AOI21_X1  g0903(.A(new_n262), .B1(new_n877), .B2(G322), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n480), .B2(new_n795), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n802), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1106), .A2(G294), .B1(new_n831), .B2(G116), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n827), .B2(new_n814), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1105), .B(new_n1108), .C1(new_n883), .C2(G303), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G150), .A2(new_n799), .B1(new_n808), .B2(G159), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT51), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n874), .A2(new_n886), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n831), .A2(G77), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n814), .A2(new_n278), .B1(new_n994), .B2(new_n817), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1112), .B(new_n1113), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n805), .B2(new_n286), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n883), .B2(G50), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1103), .A2(new_n1109), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1101), .B1(new_n790), .B2(new_n1121), .C1(new_n1041), .C2(new_n852), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1025), .A2(new_n1058), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n732), .B1(new_n1025), .B2(new_n1058), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1097), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(G390));
  NOR2_X1   g0925(.A1(new_n979), .A2(new_n925), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n714), .B(new_n862), .C1(new_n761), .C2(new_n765), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n949), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n973), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n756), .A2(new_n721), .A3(new_n964), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n973), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n863), .A2(new_n949), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n925), .B1(new_n1133), .B2(new_n973), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n935), .A2(new_n937), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n920), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n954), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(KEYINPUT39), .B2(new_n922), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1130), .B(new_n1132), .C1(new_n1134), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n925), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n948), .B1(new_n773), .B2(new_n862), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n947), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n939), .B1(new_n955), .B2(new_n926), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1142), .A2(new_n1143), .B1(new_n1129), .B2(new_n1126), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n969), .A2(new_n973), .A3(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n837), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n892), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n786), .B1(new_n342), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n883), .A2(G137), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  NAND2_X1  g0952(.A1(new_n806), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n808), .A2(G132), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n799), .A2(G128), .B1(G50), .B2(new_n796), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OR3_X1    g0956(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT53), .B1(new_n814), .B2(new_n870), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n259), .B1(new_n877), .B2(G125), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n831), .A2(G159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G116), .A2(new_n808), .B1(new_n799), .B2(G283), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n262), .B(new_n815), .C1(G294), .C2(new_n877), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n875), .A3(new_n1113), .A4(new_n1163), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n882), .A2(new_n480), .B1(new_n805), .B2(new_n488), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n1156), .A2(new_n1161), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1150), .B1(new_n1166), .B2(new_n789), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT117), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1147), .A2(new_n782), .B1(new_n1148), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n474), .A2(G330), .A3(new_n755), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n959), .A2(new_n667), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1128), .B1(new_n1131), .B2(new_n973), .ZN(new_n1173));
  INV_X1    g0973(.A(G330), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n947), .B1(new_n962), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1145), .B1(new_n1131), .B2(new_n973), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1133), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1172), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n733), .B1(new_n1146), .B2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1175), .A2(new_n1173), .B1(new_n1177), .B2(new_n1133), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n1171), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n1139), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1181), .A2(KEYINPUT116), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT116), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1169), .B1(new_n1185), .B2(new_n1186), .ZN(G378));
  NAND2_X1  g0987(.A1(new_n981), .A2(G330), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n305), .A2(new_n910), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n321), .A2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n309), .B(new_n1190), .C1(new_n319), .C2(new_n320), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1189), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n321), .A2(new_n1191), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1189), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1196), .A2(new_n1193), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1188), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n940), .A2(new_n956), .A3(new_n957), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1199), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n981), .A2(G330), .A3(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n981), .B2(G330), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1174), .B(new_n1199), .C1(new_n977), .C2(new_n980), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n958), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1207), .A3(KEYINPUT120), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT120), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1200), .A2(new_n1201), .A3(new_n1209), .A4(new_n1203), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1172), .B1(new_n1146), .B2(new_n1182), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT57), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n733), .B1(new_n1215), .B2(new_n1211), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1208), .A2(new_n782), .A3(new_n1210), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n785), .B1(new_n276), .B2(new_n892), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n814), .A2(new_n340), .B1(new_n827), .B2(new_n817), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n874), .A2(new_n495), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G58), .C2(new_n796), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT118), .Z(new_n1223));
  AOI22_X1  g1023(.A1(new_n799), .A2(G116), .B1(G68), .B2(new_n831), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT119), .Z(new_n1225));
  OAI22_X1  g1025(.A1(new_n809), .A2(new_n480), .B1(new_n344), .B2(new_n802), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G97), .B2(new_n793), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT58), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n799), .A2(G125), .B1(G137), .B2(new_n1106), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n808), .A2(G128), .B1(G132), .B2(new_n793), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n887), .A2(new_n1152), .B1(new_n831), .B2(G150), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n877), .C2(G124), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n818), .B2(new_n795), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1235), .B2(KEYINPUT59), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G50), .B1(new_n253), .B2(new_n495), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1236), .A2(new_n1239), .B1(new_n1221), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1230), .A2(new_n1231), .A3(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1219), .B1(new_n790), .B2(new_n1242), .C1(new_n1202), .C2(new_n838), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1218), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1217), .A2(new_n1244), .ZN(G375));
  NAND2_X1  g1045(.A1(new_n1182), .A2(new_n1171), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1180), .A2(new_n1035), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1179), .A2(new_n782), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n947), .A2(new_n837), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT121), .Z(new_n1250));
  AOI21_X1  g1050(.A(new_n785), .B1(new_n278), .B2(new_n892), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n883), .A2(G116), .B1(G107), .B2(new_n806), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n809), .A2(new_n827), .B1(new_n344), .B2(new_n812), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n800), .A2(new_n555), .B1(new_n488), .B2(new_n814), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n259), .B1(new_n817), .B2(new_n822), .C1(new_n795), .C2(new_n340), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n883), .A2(new_n1152), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n808), .A2(G137), .B1(G159), .B2(new_n887), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n799), .A2(G132), .B1(G58), .B2(new_n796), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1106), .A2(G150), .B1(new_n831), .B2(G50), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n874), .B1(G128), .B2(new_n877), .ZN(new_n1261));
  AND4_X1   g1061(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1252), .A2(new_n1256), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1250), .B(new_n1251), .C1(new_n790), .C2(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1248), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1247), .A2(new_n1265), .ZN(G381));
  NAND2_X1  g1066(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1267), .A2(new_n1169), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1217), .A2(new_n1244), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1060), .A2(new_n854), .A3(new_n1093), .ZN(new_n1270));
  OR3_X1    g1070(.A1(G390), .A2(G384), .A3(new_n1270), .ZN(new_n1271));
  OR4_X1    g1071(.A1(G387), .A2(new_n1269), .A3(G381), .A4(new_n1271), .ZN(G407));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G343), .C2(new_n1269), .ZN(G409));
  INV_X1    g1073(.A(G390), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G387), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n776), .B1(new_n1096), .B2(new_n1031), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n781), .B1(new_n1276), .B2(new_n1034), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1056), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT124), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1279), .A2(new_n1280), .A3(G390), .A4(new_n1011), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1270), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT123), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1282), .A2(KEYINPUT123), .A3(new_n1270), .ZN(new_n1286));
  AND4_X1   g1086(.A1(new_n1275), .A2(new_n1281), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1279), .A2(new_n1011), .A3(G390), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT124), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(G387), .A2(new_n1274), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1291), .A2(new_n1292), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1275), .A2(new_n1288), .A3(KEYINPUT125), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  INV_X1    g1097(.A(G213), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1298), .A2(G343), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1217), .A2(G378), .A3(new_n1244), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n782), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1243), .B(new_n1302), .C1(new_n1212), .C2(new_n1034), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1268), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1299), .B1(new_n1300), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1246), .B1(new_n1183), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1182), .A2(new_n1171), .A3(KEYINPUT60), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n732), .A3(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(G384), .A3(new_n1265), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1309), .B2(new_n1265), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G2897), .B(new_n1299), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1299), .A2(G2897), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1310), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1297), .B1(new_n1305), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT126), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1320), .B(new_n1297), .C1(new_n1305), .C2(new_n1317), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1305), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT122), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1305), .A2(KEYINPUT122), .A3(new_n1322), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT62), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1296), .B1(new_n1325), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1323), .A2(new_n1331), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1332), .A2(new_n1296), .A3(new_n1318), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1327), .A2(new_n1331), .A3(new_n1328), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1330), .A2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(new_n1314), .A2(new_n1310), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(KEYINPUT127), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1296), .A2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1300), .B1(KEYINPUT127), .B2(new_n1337), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1341), .B1(G375), .B2(new_n1268), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1290), .A2(new_n1295), .A3(new_n1338), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1340), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1342), .B1(new_n1340), .B2(new_n1343), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(G402));
endmodule


