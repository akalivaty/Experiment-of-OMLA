//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(new_n207));
  XOR2_X1   g0007(.A(KEYINPUT67), .B(G244), .Z(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(new_n202), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n207), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n207), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT0), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n227), .A2(G50), .A3(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n216), .B(new_n219), .C1(new_n222), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  AND2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  OAI21_X1  g0051(.A(KEYINPUT68), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(G223), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1698), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n261), .A2(G222), .B1(new_n250), .B2(G77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT69), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n256), .A2(new_n265), .A3(new_n262), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n271), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(G226), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n220), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n221), .A2(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT70), .B1(new_n223), .B2(KEYINPUT8), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(KEYINPUT70), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT71), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT71), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n286), .B(new_n282), .C1(new_n283), .C2(KEYINPUT70), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n281), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n221), .A2(new_n258), .A3(KEYINPUT72), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT72), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G20), .B2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G150), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n293), .A2(new_n294), .B1(new_n221), .B2(new_n201), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n280), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT73), .ZN(new_n298));
  INV_X1    g0098(.A(new_n297), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n280), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n297), .A2(KEYINPUT73), .A3(new_n220), .A4(new_n279), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n270), .A2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  MUX2_X1   g0103(.A(new_n297), .B(new_n303), .S(G50), .Z(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n278), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n276), .A2(G169), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT75), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n296), .A2(new_n310), .A3(new_n304), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n296), .B2(new_n304), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT9), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n305), .A2(KEYINPUT75), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT9), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n296), .A2(new_n310), .A3(new_n304), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n268), .B2(new_n275), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(G190), .B2(new_n276), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n318), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n309), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n299), .A2(new_n280), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G68), .A3(new_n302), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n280), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n292), .A2(G50), .ZN(new_n331));
  INV_X1    g0131(.A(new_n281), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(G77), .B1(G20), .B2(new_n224), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT11), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n299), .A2(new_n224), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT12), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(KEYINPUT11), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n329), .A2(new_n335), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n261), .A2(G226), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n267), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n272), .B1(G238), .B2(new_n274), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n346), .B1(new_n345), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g0149(.A(G200), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT13), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(G190), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n340), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G169), .B1(new_n348), .B2(new_n349), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n352), .A2(G179), .A3(new_n353), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(G169), .C1(new_n348), .C2(new_n349), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n355), .B1(new_n361), .B2(new_n339), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n250), .B2(new_n221), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n260), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n292), .A2(G159), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G58), .A2(G68), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n225), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G20), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT77), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n289), .B2(new_n291), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n221), .B1(new_n225), .B2(new_n368), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n366), .B(KEYINPUT16), .C1(new_n371), .C2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n259), .A2(new_n221), .A3(new_n260), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n224), .B1(new_n381), .B2(new_n364), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n367), .A2(new_n370), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n377), .A2(new_n280), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n303), .B1(new_n285), .B2(new_n287), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n285), .A2(new_n287), .A3(new_n299), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  AND2_X1   g0190(.A1(G1), .A2(G13), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G41), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(G226), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n253), .A2(KEYINPUT78), .A3(G226), .A4(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(G223), .B(new_n251), .C1(new_n248), .C2(new_n249), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n393), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n272), .ZN(new_n405));
  INV_X1    g0205(.A(new_n274), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n235), .ZN(new_n407));
  OAI21_X1  g0207(.A(G169), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n272), .B1(G232), .B2(new_n274), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n396), .B2(new_n397), .ZN(new_n411));
  OAI211_X1 g0211(.A(G179), .B(new_n409), .C1(new_n411), .C2(new_n393), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n389), .A2(new_n390), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n390), .B1(new_n389), .B2(new_n413), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(G190), .B(new_n409), .C1(new_n411), .C2(new_n393), .ZN(new_n417));
  OAI21_X1  g0217(.A(G200), .B1(new_n404), .B2(new_n407), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n385), .A2(new_n388), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n420), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n252), .A2(G238), .A3(new_n255), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n261), .A2(G232), .B1(new_n250), .B2(G107), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n393), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n405), .B1(new_n406), .B2(new_n208), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n277), .ZN(new_n429));
  INV_X1    g0229(.A(G169), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n426), .B2(new_n427), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n293), .A2(new_n283), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT15), .B(G87), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n433), .A2(new_n281), .B1(new_n221), .B2(new_n202), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n280), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n202), .B1(new_n270), .B2(G20), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n326), .A2(new_n436), .B1(new_n202), .B2(new_n299), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n429), .A2(new_n431), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n438), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n428), .B2(new_n320), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n442), .A2(KEYINPUT74), .B1(G190), .B2(new_n428), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n362), .A2(new_n416), .A3(new_n423), .A4(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT81), .B1(new_n325), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n318), .A2(new_n322), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT10), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n308), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n446), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G303), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n259), .A2(new_n457), .A3(new_n260), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G264), .A2(G1698), .ZN(new_n459));
  INV_X1    g0259(.A(G257), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G1698), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n458), .B(new_n267), .C1(new_n250), .C2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n269), .B1(new_n391), .B2(new_n392), .ZN(new_n463));
  INV_X1    g0263(.A(G41), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n463), .A2(new_n465), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n465), .A3(new_n469), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G270), .A3(new_n393), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n462), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n473), .A2(G169), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n270), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n297), .A2(new_n475), .A3(new_n220), .A4(new_n279), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G116), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n299), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n279), .A2(new_n220), .B1(G20), .B2(new_n479), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n221), .C1(G33), .C2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n481), .A2(KEYINPUT20), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT20), .B1(new_n481), .B2(new_n484), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n478), .B(new_n480), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT21), .B1(new_n474), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G190), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n473), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n480), .B1(new_n476), .B2(new_n479), .ZN(new_n492));
  INV_X1    g0292(.A(new_n486), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n481), .A2(KEYINPUT20), .A3(new_n484), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n473), .A2(G200), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(KEYINPUT21), .A2(G169), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n485), .A2(new_n486), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n473), .B(new_n498), .C1(new_n499), .C2(new_n492), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT85), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n473), .A2(new_n277), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n500), .A2(new_n501), .B1(new_n487), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n487), .A2(KEYINPUT85), .A3(new_n473), .A4(new_n498), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT86), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n473), .A2(new_n498), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n501), .B1(new_n506), .B2(new_n495), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n487), .ZN(new_n508));
  AND4_X1   g0308(.A1(KEYINPUT86), .A2(new_n507), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n489), .B(new_n497), .C1(new_n505), .C2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G257), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n511));
  OAI211_X1 g0311(.A(G250), .B(new_n251), .C1(new_n248), .C2(new_n249), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n267), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n471), .A2(G264), .A3(new_n393), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(new_n470), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT90), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n471), .A2(KEYINPUT90), .A3(G264), .A4(new_n393), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n515), .A2(new_n520), .A3(new_n470), .A4(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n518), .A2(G169), .B1(new_n523), .B2(G179), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT23), .B1(new_n221), .B2(G107), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  INV_X1    g0326(.A(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(G20), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT88), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT88), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n525), .A2(new_n528), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n221), .B(G87), .C1(new_n248), .C2(new_n249), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n253), .A2(new_n537), .A3(new_n221), .A4(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g0339(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n534), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n280), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT89), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT89), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n280), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n527), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT25), .B1(new_n299), .B2(new_n527), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n527), .B2(new_n476), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n524), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n517), .A2(new_n490), .B1(new_n522), .B2(new_n320), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n547), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n297), .A2(G97), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n477), .B2(G97), .ZN(new_n558));
  OAI21_X1  g0358(.A(G107), .B1(new_n363), .B2(new_n365), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n202), .B1(new_n289), .B2(new_n291), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  AND2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n527), .A2(KEYINPUT6), .A3(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n560), .B1(new_n566), .B2(G20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT82), .B1(new_n568), .B2(new_n280), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT82), .ZN(new_n570));
  AOI211_X1 g0370(.A(new_n570), .B(new_n330), .C1(new_n559), .C2(new_n567), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n558), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n471), .A2(G257), .A3(new_n393), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n470), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT84), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n251), .A2(G244), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n259), .B2(new_n260), .ZN(new_n577));
  XNOR2_X1  g0377(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G250), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n259), .B2(new_n260), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n577), .A2(KEYINPUT4), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(new_n251), .C1(new_n248), .C2(new_n249), .ZN(new_n584));
  XOR2_X1   g0384(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT84), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n579), .A2(new_n582), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  AOI211_X1 g0387(.A(G179), .B(new_n574), .C1(new_n587), .C2(new_n267), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n267), .ZN(new_n590));
  INV_X1    g0390(.A(new_n574), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n430), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n572), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n527), .A2(KEYINPUT6), .A3(G97), .ZN(new_n595));
  XNOR2_X1  g0395(.A(G97), .B(G107), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n561), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n597), .A2(new_n221), .B1(new_n293), .B2(new_n202), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n527), .B1(new_n381), .B2(new_n364), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n280), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n570), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n568), .A2(KEYINPUT82), .A3(new_n280), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n574), .B1(new_n587), .B2(new_n267), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  AOI211_X1 g0405(.A(G190), .B(new_n574), .C1(new_n587), .C2(new_n267), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n603), .B(new_n558), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n253), .A2(new_n221), .A3(G68), .ZN(new_n608));
  INV_X1    g0408(.A(G87), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n483), .A3(new_n527), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n343), .A2(new_n221), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT19), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n281), .B2(new_n483), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n608), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n280), .B1(new_n299), .B2(new_n433), .ZN(new_n616));
  INV_X1    g0416(.A(new_n433), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n477), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n270), .A2(new_n269), .A3(G45), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n580), .B1(new_n466), .B2(G1), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n393), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(G238), .A2(G1698), .ZN(new_n623));
  INV_X1    g0423(.A(G244), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n624), .B2(G1698), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n625), .A2(new_n253), .B1(G33), .B2(G116), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n626), .B2(new_n393), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n430), .ZN(new_n628));
  INV_X1    g0428(.A(new_n622), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(G1698), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(G238), .B2(G1698), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n631), .A2(new_n250), .B1(new_n258), .B2(new_n479), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n632), .B2(new_n267), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n277), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n619), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(G190), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n627), .A2(G200), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n477), .A2(G87), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n616), .A4(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n556), .A2(new_n594), .A3(new_n607), .A4(new_n640), .ZN(new_n641));
  NOR4_X1   g0441(.A1(new_n456), .A2(new_n510), .A3(new_n553), .A4(new_n641), .ZN(G372));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n361), .A2(new_n339), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n340), .A2(new_n350), .A3(new_n354), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n440), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n423), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n416), .B1(new_n449), .B2(new_n450), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n643), .B1(new_n649), .B2(new_n308), .ZN(new_n650));
  INV_X1    g0450(.A(new_n423), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n644), .B2(new_n646), .ZN(new_n652));
  INV_X1    g0452(.A(new_n416), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n652), .A2(new_n653), .B1(new_n324), .B2(new_n323), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(KEYINPUT91), .A3(new_n309), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n594), .A2(new_n607), .A3(new_n640), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n507), .A2(new_n504), .A3(new_n508), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n488), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n551), .B1(new_n544), .B2(new_n546), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n524), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(new_n661), .A3(new_n556), .ZN(new_n662));
  INV_X1    g0462(.A(new_n635), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n635), .A2(new_n639), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n594), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n588), .B1(new_n430), .B2(new_n592), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n572), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n663), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n656), .B1(new_n456), .B2(new_n671), .ZN(G369));
  NAND3_X1  g0472(.A1(new_n270), .A2(new_n221), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n495), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n658), .B2(new_n488), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n510), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n534), .A2(new_n539), .ZN(new_n685));
  INV_X1    g0485(.A(new_n540), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n545), .B1(new_n689), .B2(new_n280), .ZN(new_n690));
  INV_X1    g0490(.A(new_n546), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n552), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n524), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n556), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n660), .A2(new_n679), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n695), .A2(new_n696), .B1(new_n694), .B2(new_n679), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n684), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n695), .A2(new_n696), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT86), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n658), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n503), .A2(KEYINPUT86), .A3(new_n504), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n488), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n678), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n699), .A2(new_n704), .B1(new_n553), .B2(new_n679), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n217), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n610), .A2(G116), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT92), .Z(new_n710));
  NOR3_X1   g0510(.A1(new_n708), .A2(new_n710), .A3(new_n270), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n230), .B2(new_n708), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT28), .Z(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n520), .A2(new_n521), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n502), .A2(new_n715), .A3(new_n515), .A4(new_n633), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n716), .B2(new_n592), .ZN(new_n717));
  AND4_X1   g0517(.A1(new_n515), .A2(new_n633), .A3(new_n520), .A4(new_n521), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n502), .A4(new_n604), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n473), .A2(new_n277), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n627), .A2(KEYINPUT93), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n722), .B(new_n622), .C1(new_n626), .C2(new_n393), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n592), .A3(new_n522), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n717), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n726), .B2(new_n678), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n497), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n488), .B(new_n731), .C1(new_n701), .C2(new_n702), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n678), .B1(new_n692), .B2(new_n693), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(new_n657), .A4(new_n556), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n594), .A2(new_n607), .A3(new_n640), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n551), .B(new_n554), .C1(new_n544), .C2(new_n546), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(KEYINPUT94), .A3(new_n732), .A4(new_n733), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n730), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G330), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n678), .B1(new_n662), .B2(new_n669), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n489), .B1(new_n505), .B2(new_n509), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT95), .B1(new_n747), .B2(new_n553), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT95), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n694), .A2(new_n703), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(new_n739), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n678), .B1(new_n751), .B2(new_n669), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n746), .B1(new_n752), .B2(new_n745), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n743), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n713), .B1(new_n754), .B2(G1), .ZN(G364));
  AND2_X1   g0555(.A1(new_n221), .A2(G13), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n270), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n708), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n684), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n682), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n707), .A2(new_n250), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G355), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G116), .B2(new_n217), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n707), .A2(new_n253), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G45), .B2(new_n229), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n766), .A2(KEYINPUT96), .B1(G45), .B2(new_n243), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n220), .B1(G20), .B2(new_n430), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n759), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n221), .A2(G179), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G190), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n253), .B1(new_n780), .B2(G329), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n490), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n277), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n781), .B1(new_n457), .B2(new_n782), .C1(new_n783), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  NAND2_X1  g0589(.A1(G20), .A2(G179), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT97), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n778), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n784), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n789), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n777), .A2(new_n490), .A3(G200), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT99), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n788), .B(new_n797), .C1(G283), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n793), .A2(G200), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT98), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT98), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(new_n490), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT33), .B(G317), .Z(new_n808));
  NAND2_X1  g0608(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n490), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G326), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n803), .B1(new_n807), .B2(new_n808), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n787), .A2(new_n483), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n782), .A2(new_n609), .ZN(new_n815));
  OR3_X1    g0615(.A1(new_n814), .A2(new_n250), .A3(new_n815), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n223), .A2(new_n795), .B1(new_n794), .B2(new_n202), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n780), .A2(G159), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT32), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n801), .A2(new_n527), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n816), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G50), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n224), .B2(new_n807), .C1(new_n811), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n776), .B1(new_n824), .B2(new_n773), .ZN(new_n825));
  INV_X1    g0625(.A(new_n772), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n682), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n761), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NOR2_X1   g0629(.A1(new_n439), .A2(new_n678), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n443), .A2(new_n444), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n441), .B2(new_n679), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n832), .B2(new_n439), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(new_n744), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(new_n743), .ZN(new_n836));
  INV_X1    g0636(.A(new_n759), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n743), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n773), .A2(new_n770), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n837), .B1(new_n202), .B2(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n250), .B1(new_n779), .B2(new_n789), .C1(new_n787), .C2(new_n483), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n479), .A2(new_n794), .B1(new_n795), .B2(new_n783), .ZN(new_n843));
  INV_X1    g0643(.A(new_n782), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n842), .B(new_n843), .C1(G107), .C2(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n609), .B2(new_n801), .C1(new_n811), .C2(new_n457), .ZN(new_n846));
  INV_X1    g0646(.A(new_n807), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(G283), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n795), .ZN(new_n849));
  INV_X1    g0649(.A(new_n794), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n849), .B1(new_n850), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n294), .B2(new_n807), .C1(new_n811), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT34), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n782), .A2(new_n822), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n253), .B1(new_n779), .B2(new_n856), .C1(new_n787), .C2(new_n223), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n855), .B(new_n857), .C1(G68), .C2(new_n802), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n848), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n773), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n841), .B1(new_n771), .B2(new_n833), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n839), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  AOI21_X1  g0663(.A(new_n830), .B1(new_n744), .B2(new_n833), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n415), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n389), .A2(new_n390), .A3(new_n413), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n419), .A2(new_n422), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n285), .A2(new_n287), .A3(new_n299), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n285), .A2(new_n287), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n303), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n367), .A2(KEYINPUT77), .A3(new_n370), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n375), .B1(new_n373), .B2(new_n374), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n381), .A2(new_n364), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n874), .A2(new_n875), .B1(new_n876), .B2(G68), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n330), .B1(new_n877), .B2(KEYINPUT16), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n366), .B1(new_n371), .B2(new_n376), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n378), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n873), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n676), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n870), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n419), .B1(new_n881), .B2(new_n676), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n878), .A2(new_n880), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n886), .A2(new_n388), .B1(new_n408), .B2(new_n412), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n389), .A2(new_n413), .ZN(new_n889));
  INV_X1    g0689(.A(new_n676), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n389), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n889), .A2(new_n891), .A3(new_n892), .A4(new_n419), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n883), .A2(new_n884), .A3(new_n894), .A4(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n888), .A2(new_n893), .ZN(new_n897));
  INV_X1    g0697(.A(new_n882), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n416), .B2(new_n423), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n894), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(KEYINPUT100), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n339), .A2(new_n678), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n362), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n361), .A2(new_n339), .A3(new_n678), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n865), .A2(new_n895), .A3(new_n902), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n653), .A2(new_n676), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n361), .A2(new_n339), .A3(new_n679), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n889), .A2(new_n891), .A3(new_n419), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(new_n892), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n891), .B1(new_n416), .B2(new_n423), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n896), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n901), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n909), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n455), .A2(new_n753), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n656), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT102), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n729), .B1(new_n727), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n726), .A2(KEYINPUT102), .A3(KEYINPUT31), .A4(new_n678), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n736), .B2(new_n740), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n906), .A2(new_n833), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT103), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n925), .A2(new_n926), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n679), .B1(new_n660), .B2(new_n524), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n932), .A2(new_n737), .A3(new_n738), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT94), .B1(new_n933), .B2(new_n732), .ZN(new_n934));
  NOR4_X1   g0734(.A1(new_n641), .A2(new_n932), .A3(new_n510), .A4(new_n735), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT103), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n906), .A2(new_n833), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n916), .B2(new_n901), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n930), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n936), .A2(new_n902), .A3(new_n938), .A4(new_n895), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n455), .A2(new_n936), .ZN(new_n947));
  OAI21_X1  g0747(.A(G330), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n946), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n923), .A2(new_n949), .B1(new_n270), .B2(new_n756), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n923), .B2(new_n949), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(G116), .A4(new_n222), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT36), .Z(new_n955));
  NAND3_X1  g0755(.A1(new_n230), .A2(G77), .A3(new_n368), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n822), .A2(G68), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n270), .B(G13), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n951), .A2(new_n955), .A3(new_n958), .ZN(G367));
  NAND2_X1  g0759(.A1(new_n699), .A2(new_n704), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n697), .B2(new_n704), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(new_n683), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n754), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n572), .A2(new_n678), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n594), .A2(new_n607), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n667), .A2(new_n572), .A3(new_n678), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n705), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT45), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n705), .A2(new_n969), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(KEYINPUT44), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT104), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n972), .A2(KEYINPUT44), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n977), .A2(new_n973), .A3(new_n974), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT105), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n698), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n965), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n971), .A3(new_n975), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT105), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(new_n698), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n754), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n708), .B(KEYINPUT41), .Z(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n758), .B1(new_n989), .B2(KEYINPUT106), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT106), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n991), .A3(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n699), .A2(new_n704), .A3(new_n969), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n594), .B1(new_n694), .B2(new_n967), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n994), .A2(KEYINPUT42), .B1(new_n679), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(KEYINPUT42), .B2(new_n994), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n616), .A2(new_n638), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n678), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n640), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n635), .A2(new_n1000), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n997), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n998), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n698), .B1(new_n967), .B2(new_n968), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n993), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1004), .A2(new_n772), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n765), .A2(new_n239), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n775), .B1(new_n707), .B2(new_n617), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n837), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n810), .A2(G143), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n787), .A2(new_n224), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n250), .B1(new_n780), .B2(G137), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n223), .C2(new_n782), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G150), .B2(new_n849), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1016), .B(new_n1021), .C1(new_n202), .C2(new_n801), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n807), .A2(new_n372), .B1(new_n822), .B2(new_n794), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(KEYINPUT108), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT108), .B2(new_n1023), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n782), .A2(new_n479), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT46), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n802), .A2(G97), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n850), .A2(G283), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n786), .A2(G107), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT107), .B(G317), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n253), .B1(new_n780), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1027), .B(new_n1033), .C1(G303), .C2(new_n849), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n783), .B2(new_n807), .C1(new_n789), .C2(new_n811), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1025), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT47), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n860), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1012), .B(new_n1015), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1011), .A2(new_n1041), .ZN(G387));
  OAI21_X1  g0842(.A(new_n250), .B1(new_n779), .B2(new_n812), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G303), .A2(new_n850), .B1(new_n849), .B2(new_n1031), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n789), .B2(new_n807), .C1(new_n811), .C2(new_n796), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G294), .A2(new_n844), .B1(new_n786), .B2(G283), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT49), .Z(new_n1051));
  AOI211_X1 g0851(.A(new_n1043), .B(new_n1051), .C1(G116), .C2(new_n802), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n807), .A2(new_n872), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n253), .B1(new_n779), .B2(new_n294), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n787), .A2(new_n433), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G77), .C2(new_n844), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G50), .A2(new_n849), .B1(new_n850), .B2(G68), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n1028), .A3(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1053), .B(new_n1058), .C1(G159), .C2(new_n810), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n773), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n765), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n236), .B2(G45), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n710), .B2(new_n762), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n283), .A2(G50), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT50), .Z(new_n1065));
  OAI21_X1  g0865(.A(new_n466), .B1(new_n224), .B2(new_n202), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1065), .A2(new_n710), .A3(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1063), .A2(new_n1067), .B1(G107), .B2(new_n217), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n837), .B1(new_n1068), .B2(new_n774), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1060), .B(new_n1069), .C1(new_n697), .C2(new_n826), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n963), .A2(new_n758), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT109), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n708), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n965), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(KEYINPUT110), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n754), .B2(new_n963), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1074), .A2(KEYINPUT110), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1070), .B(new_n1072), .C1(new_n1076), .C2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n982), .A2(new_n980), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n976), .A2(new_n698), .A3(new_n978), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1080), .A3(new_n758), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1061), .A2(new_n246), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n774), .B1(new_n217), .B2(new_n483), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n759), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n250), .B1(new_n779), .B2(new_n796), .C1(new_n787), .C2(new_n479), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n794), .A2(new_n783), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n844), .A2(G283), .ZN(new_n1087));
  NOR4_X1   g0887(.A1(new_n820), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n810), .A2(G317), .B1(G311), .B2(new_n849), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT52), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1088), .B1(new_n457), .B2(new_n807), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1093), .A2(KEYINPUT112), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n810), .A2(G150), .B1(G159), .B2(new_n849), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  NOR2_X1   g0896(.A1(new_n801), .A2(new_n609), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n787), .A2(new_n202), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n250), .B(new_n1098), .C1(G143), .C2(new_n780), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n224), .B2(new_n782), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n794), .A2(new_n283), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n847), .B2(G50), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1097), .B(new_n1100), .C1(new_n1102), .C2(KEYINPUT111), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1096), .B(new_n1103), .C1(KEYINPUT111), .C2(new_n1102), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1093), .A2(KEYINPUT112), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1094), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1084), .B1(new_n1106), .B2(new_n773), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n826), .B2(new_n969), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1081), .A2(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT113), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(KEYINPUT113), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n981), .A2(new_n985), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1073), .B1(new_n1114), .B2(new_n964), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(G390));
  NAND3_X1  g0918(.A1(new_n936), .A2(G330), .A3(new_n938), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n906), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n910), .B1(new_n864), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n912), .A3(new_n918), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n911), .B1(new_n916), .B2(new_n901), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n832), .A2(new_n439), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n830), .B1(new_n752), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n1120), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1119), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n730), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n934), .B2(new_n935), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1131), .A2(G330), .A3(new_n833), .A4(new_n906), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1127), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n736), .A2(new_n740), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n742), .B1(new_n1134), .B2(new_n931), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n455), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n921), .A2(new_n1136), .A3(new_n656), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT114), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1131), .A2(G330), .A3(new_n833), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1140), .A2(new_n1120), .B1(new_n1135), .B2(new_n938), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1141), .B2(new_n864), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n741), .A2(new_n742), .A3(new_n834), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1119), .B1(new_n1143), .B2(new_n906), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(KEYINPUT114), .A3(new_n865), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1132), .A2(new_n1125), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n906), .B1(new_n1135), .B2(new_n833), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1138), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT115), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1151), .B2(new_n1133), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1149), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1128), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1122), .A2(new_n1126), .A3(new_n1132), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1154), .A2(new_n1158), .A3(KEYINPUT115), .A4(new_n1138), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n708), .B1(new_n1133), .B2(new_n1151), .C1(new_n1153), .C2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n912), .A2(new_n770), .A3(new_n918), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n872), .A2(new_n840), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n801), .A2(new_n224), .B1(new_n783), .B2(new_n779), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n810), .A2(G283), .B1(KEYINPUT117), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(KEYINPUT117), .B2(new_n1163), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1098), .A2(new_n253), .A3(new_n815), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G97), .A2(new_n850), .B1(new_n849), .B2(G116), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n807), .C2(new_n527), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT116), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n253), .B1(new_n801), .B2(new_n822), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n847), .A2(G137), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1172));
  INV_X1    g0972(.A(G125), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n787), .A2(new_n372), .B1(new_n1173), .B2(new_n779), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT54), .B(G143), .Z(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n850), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT53), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n782), .A2(new_n294), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n795), .A2(new_n856), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1180));
  INV_X1    g0980(.A(G128), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1176), .B(new_n1180), .C1(new_n811), .C2(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1165), .A2(new_n1168), .B1(new_n1172), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n837), .B(new_n1162), .C1(new_n1183), .C2(new_n773), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1133), .A2(new_n758), .B1(new_n1161), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1160), .A2(new_n1185), .ZN(G378));
  INV_X1    g0986(.A(new_n840), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n759), .B1(G50), .B2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1189));
  OR2_X1    g0989(.A1(new_n451), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n451), .A2(new_n1189), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n676), .B1(new_n314), .B2(new_n316), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1190), .A2(new_n1193), .A3(new_n1191), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n771), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1018), .B1(new_n795), .B2(new_n527), .C1(new_n433), .C2(new_n794), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n802), .A2(G58), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n253), .A2(G41), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G283), .B2(new_n780), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1200), .B(new_n1203), .C1(new_n202), .C2(new_n782), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT118), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT118), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n483), .C2(new_n807), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1199), .B(new_n1208), .C1(G116), .C2(new_n810), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT58), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n844), .A2(new_n1175), .B1(new_n786), .B2(G150), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n794), .B2(new_n852), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G128), .B2(new_n849), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n856), .B2(new_n807), .C1(new_n811), .C2(new_n1173), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n802), .A2(G159), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1209), .A2(KEYINPUT58), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1202), .B(new_n822), .C1(G33), .C2(G41), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1210), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1188), .B(new_n1198), .C1(new_n773), .C2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1137), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n942), .A2(new_n945), .A3(G330), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1197), .A2(new_n942), .A3(G330), .A4(new_n945), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n920), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1227), .A2(new_n1228), .A3(new_n920), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(KEYINPUT121), .A3(new_n1232), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n1229), .A2(new_n1230), .A3(KEYINPUT121), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1224), .A2(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n708), .A2(KEYINPUT57), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1223), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1141), .A2(new_n1139), .A3(new_n864), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT114), .B1(new_n1144), .B2(new_n865), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1150), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1133), .A3(new_n1137), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT115), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1151), .A2(new_n1152), .A3(new_n1133), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1138), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1073), .A2(KEYINPUT57), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n757), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT120), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1231), .A2(KEYINPUT119), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1232), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n920), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT119), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT120), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1251), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1248), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1238), .A2(new_n1258), .ZN(G375));
  AOI22_X1  g1059(.A1(new_n847), .A2(G116), .B1(G107), .B2(new_n850), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n783), .B2(new_n811), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT122), .Z(new_n1262));
  NOR2_X1   g1062(.A1(new_n801), .A2(new_n202), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1055), .B1(new_n849), .B2(G283), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT123), .Z(new_n1265));
  OAI221_X1 g1065(.A(new_n250), .B1(new_n779), .B2(new_n457), .C1(new_n483), .C2(new_n782), .ZN(new_n1266));
  NOR4_X1   g1066(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1267), .A2(KEYINPUT124), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n810), .A2(G132), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n253), .B1(new_n779), .B2(new_n1181), .C1(new_n787), .C2(new_n822), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n852), .A2(new_n795), .B1(new_n794), .B2(new_n294), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(G159), .C2(new_n844), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n847), .A2(new_n1175), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1272), .A3(new_n1273), .A4(new_n1200), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1267), .B2(KEYINPUT124), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n773), .B1(new_n1268), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n837), .B1(new_n224), .B2(new_n840), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(new_n771), .C2(new_n906), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1241), .B2(new_n758), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n988), .B1(new_n1154), .B2(new_n1138), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1149), .B(new_n1137), .C1(new_n1142), .C2(new_n1145), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1280), .B1(new_n1281), .B2(new_n1282), .ZN(G381));
  NAND3_X1  g1083(.A1(new_n1011), .A2(new_n1041), .A3(new_n1117), .ZN(new_n1284));
  OR2_X1    g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1284), .A2(G384), .A3(G381), .A4(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(G375), .A2(G378), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(G407));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1286), .B2(new_n677), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(G213), .ZN(G409));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  OAI21_X1  g1091(.A(KEYINPUT60), .B1(new_n1282), .B2(KEYINPUT125), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT60), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1293), .B(new_n1294), .C1(new_n1241), .C2(new_n1137), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1151), .A2(new_n1073), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1280), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n862), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(G384), .A3(new_n1280), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n677), .A2(G213), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1238), .A2(new_n1258), .A3(G378), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1249), .B1(new_n1231), .B2(KEYINPUT119), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1252), .A2(new_n1253), .A3(KEYINPUT120), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1232), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1250), .A2(new_n1254), .A3(new_n1251), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1307), .A2(new_n1224), .A3(new_n988), .A4(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1223), .B1(new_n1235), .B2(new_n758), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1160), .A2(new_n1185), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n1301), .B(new_n1303), .C1(new_n1304), .C2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1291), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1297), .A2(G384), .A3(new_n1280), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1297), .B2(new_n1280), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT126), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1299), .A2(new_n1320), .A3(new_n1300), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1303), .A2(G2897), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1304), .A2(new_n1313), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1302), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1301), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1326), .A2(new_n1329), .A3(new_n1302), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1316), .A2(new_n1328), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1009), .B1(new_n990), .B2(new_n992), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1041), .ZN(new_n1334));
  OAI21_X1  g1134(.A(G390), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(G393), .B(G396), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1284), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1284), .B2(new_n1335), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1332), .A2(new_n1340), .ZN(new_n1341));
  OR2_X1    g1141(.A1(new_n1314), .A2(KEYINPUT63), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1314), .A2(KEYINPUT63), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1339), .A2(new_n1342), .A3(new_n1343), .A4(new_n1328), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1341), .A2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1312), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1304), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1347), .B(new_n1301), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1348), .B(new_n1339), .ZN(G402));
endmodule


