

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U324 ( .A(G22GAT), .B(G141GAT), .Z(n291) );
  XOR2_X1 U325 ( .A(n390), .B(n347), .Z(n292) );
  XNOR2_X1 U326 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n409) );
  XNOR2_X1 U327 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U328 ( .A(n360), .B(n359), .ZN(n361) );
  INV_X1 U329 ( .A(G190GAT), .ZN(n452) );
  XNOR2_X1 U330 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n294) );
  XNOR2_X1 U333 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U335 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n296) );
  XNOR2_X1 U336 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U338 ( .A(n298), .B(n297), .Z(n300) );
  XOR2_X1 U339 ( .A(G50GAT), .B(G162GAT), .Z(n412) );
  XOR2_X1 U340 ( .A(G134GAT), .B(KEYINPUT77), .Z(n312) );
  XNOR2_X1 U341 ( .A(n412), .B(n312), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U343 ( .A(G99GAT), .B(G85GAT), .Z(n363) );
  XOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .Z(n333) );
  XOR2_X1 U345 ( .A(n363), .B(n333), .Z(n302) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U348 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U349 ( .A(KEYINPUT68), .B(KEYINPUT7), .Z(n306) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G29GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U352 ( .A(KEYINPUT8), .B(n307), .Z(n362) );
  XNOR2_X1 U353 ( .A(n362), .B(G92GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n551) );
  XOR2_X1 U355 ( .A(G120GAT), .B(KEYINPUT83), .Z(n311) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n431) );
  XOR2_X1 U358 ( .A(n312), .B(n431), .Z(n314) );
  NAND2_X1 U359 ( .A1(G225GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U361 ( .A(n315), .B(KEYINPUT6), .Z(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT2), .B(KEYINPUT92), .Z(n317) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n425) );
  XNOR2_X1 U365 ( .A(n425), .B(KEYINPUT94), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G162GAT), .Z(n321) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(G148GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U370 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U371 ( .A(G57GAT), .B(KEYINPUT93), .Z(n325) );
  XNOR2_X1 U372 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n327) );
  XNOR2_X1 U375 ( .A(G127GAT), .B(G155GAT), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n540) );
  XNOR2_X1 U379 ( .A(G8GAT), .B(G183GAT), .ZN(n332) );
  XNOR2_X1 U380 ( .A(n332), .B(G211GAT), .ZN(n380) );
  XOR2_X1 U381 ( .A(KEYINPUT95), .B(n333), .Z(n335) );
  NAND2_X1 U382 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n338) );
  XOR2_X1 U384 ( .A(G64GAT), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n374) );
  XOR2_X1 U387 ( .A(n338), .B(n374), .Z(n344) );
  XOR2_X1 U388 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n340) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n436) );
  XOR2_X1 U391 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n342) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n413) );
  XNOR2_X1 U394 ( .A(n436), .B(n413), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n380), .B(n345), .ZN(n513) );
  XOR2_X1 U397 ( .A(G1GAT), .B(KEYINPUT69), .Z(n390) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(G50GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n291), .B(n346), .ZN(n347) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n292), .B(n348), .ZN(n360) );
  XOR2_X1 U402 ( .A(G15GAT), .B(G113GAT), .Z(n350) );
  XNOR2_X1 U403 ( .A(G169GAT), .B(G197GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U405 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n352) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U408 ( .A(n354), .B(n353), .Z(n358) );
  XOR2_X1 U409 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n356) );
  XNOR2_X1 U410 ( .A(KEYINPUT70), .B(KEYINPUT64), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n567) );
  XNOR2_X1 U413 ( .A(G120GAT), .B(n363), .ZN(n364) );
  XNOR2_X1 U414 ( .A(n364), .B(KEYINPUT73), .ZN(n378) );
  XOR2_X1 U415 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n366) );
  XNOR2_X1 U416 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n366), .B(n365), .ZN(n371) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(G78GAT), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n367), .B(G148GAT), .ZN(n424) );
  XNOR2_X1 U420 ( .A(n424), .B(KEYINPUT31), .ZN(n369) );
  AND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U423 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U424 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n373) );
  XNOR2_X1 U425 ( .A(G71GAT), .B(G57GAT), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n379) );
  XNOR2_X1 U427 ( .A(n374), .B(n379), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n378), .B(n377), .ZN(n399) );
  INV_X1 U430 ( .A(n399), .ZN(n572) );
  XNOR2_X1 U431 ( .A(n380), .B(n379), .ZN(n394) );
  XOR2_X1 U432 ( .A(G22GAT), .B(G155GAT), .Z(n417) );
  XOR2_X1 U433 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XOR2_X1 U434 ( .A(n417), .B(n432), .Z(n382) );
  NAND2_X1 U435 ( .A1(G231GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U437 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n384) );
  XNOR2_X1 U438 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(n386), .B(n385), .Z(n392) );
  XOR2_X1 U441 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n388) );
  XNOR2_X1 U442 ( .A(G78GAT), .B(G64GAT), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n575) );
  XNOR2_X1 U447 ( .A(KEYINPUT36), .B(n551), .ZN(n579) );
  NOR2_X1 U448 ( .A1(n575), .A2(n579), .ZN(n395) );
  XOR2_X1 U449 ( .A(KEYINPUT45), .B(n395), .Z(n396) );
  NOR2_X1 U450 ( .A1(n399), .A2(n396), .ZN(n397) );
  NAND2_X1 U451 ( .A1(n567), .A2(n397), .ZN(n407) );
  INV_X1 U452 ( .A(KEYINPUT41), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n498) );
  INV_X1 U454 ( .A(n567), .ZN(n543) );
  NAND2_X1 U455 ( .A1(n498), .A2(n543), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n400), .B(KEYINPUT46), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n575), .B(KEYINPUT110), .ZN(n563) );
  NAND2_X1 U458 ( .A1(n401), .A2(n563), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n402), .B(KEYINPUT111), .ZN(n403) );
  NAND2_X1 U460 ( .A1(n403), .A2(n551), .ZN(n405) );
  XOR2_X1 U461 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  NAND2_X1 U463 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n408), .B(KEYINPUT48), .ZN(n539) );
  NAND2_X1 U465 ( .A1(n513), .A2(n539), .ZN(n410) );
  NOR2_X1 U466 ( .A1(n540), .A2(n411), .ZN(n566) );
  XOR2_X1 U467 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U470 ( .A(n416), .B(KEYINPUT90), .Z(n419) );
  XNOR2_X1 U471 ( .A(n417), .B(KEYINPUT24), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U473 ( .A(G204GAT), .B(G211GAT), .Z(n421) );
  XNOR2_X1 U474 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U476 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n463) );
  NAND2_X1 U479 ( .A1(n566), .A2(n463), .ZN(n429) );
  XOR2_X1 U480 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n430), .B(KEYINPUT121), .ZN(n451) );
  XOR2_X1 U483 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U484 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U486 ( .A(n435), .B(G71GAT), .Z(n438) );
  XNOR2_X1 U487 ( .A(n436), .B(G176GAT), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U489 ( .A(G134GAT), .B(G190GAT), .Z(n440) );
  XNOR2_X1 U490 ( .A(G43GAT), .B(G99GAT), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U492 ( .A(n442), .B(n441), .Z(n450) );
  XOR2_X1 U493 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n444) );
  XNOR2_X1 U494 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U496 ( .A(G183GAT), .B(KEYINPUT86), .Z(n446) );
  XNOR2_X1 U497 ( .A(KEYINPUT87), .B(KEYINPUT20), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n522) );
  NAND2_X1 U501 ( .A1(n451), .A2(n522), .ZN(n562) );
  NOR2_X1 U502 ( .A1(n551), .A2(n562), .ZN(n455) );
  XNOR2_X1 U503 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n453) );
  XOR2_X1 U504 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n473) );
  NOR2_X1 U505 ( .A1(n567), .A2(n399), .ZN(n485) );
  XOR2_X1 U506 ( .A(KEYINPUT27), .B(n513), .Z(n464) );
  INV_X1 U507 ( .A(n464), .ZN(n457) );
  NOR2_X1 U508 ( .A1(n463), .A2(n522), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n456), .B(KEYINPUT26), .ZN(n565) );
  NAND2_X1 U510 ( .A1(n457), .A2(n565), .ZN(n542) );
  NAND2_X1 U511 ( .A1(n513), .A2(n522), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n458), .A2(n463), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  XOR2_X1 U514 ( .A(KEYINPUT96), .B(n460), .Z(n461) );
  AND2_X1 U515 ( .A1(n542), .A2(n461), .ZN(n462) );
  NOR2_X1 U516 ( .A1(n540), .A2(n462), .ZN(n467) );
  XOR2_X1 U517 ( .A(n463), .B(KEYINPUT28), .Z(n518) );
  NOR2_X1 U518 ( .A1(n518), .A2(n464), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n540), .A2(n465), .ZN(n524) );
  NOR2_X1 U520 ( .A1(n522), .A2(n524), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n482) );
  INV_X1 U522 ( .A(n575), .ZN(n548) );
  NAND2_X1 U523 ( .A1(n548), .A2(n551), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT82), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT16), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n482), .A2(n470), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT97), .B(n471), .Z(n499) );
  AND2_X1 U528 ( .A1(n485), .A2(n499), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n479), .A2(n540), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U531 ( .A(G1GAT), .B(n474), .Z(G1324GAT) );
  NAND2_X1 U532 ( .A1(n513), .A2(n479), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U535 ( .A1(n479), .A2(n522), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U537 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NAND2_X1 U538 ( .A1(n479), .A2(n518), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT100), .ZN(n481) );
  XNOR2_X1 U540 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  NOR2_X1 U541 ( .A1(n579), .A2(n482), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n575), .A2(n483), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n484), .ZN(n511) );
  NAND2_X1 U544 ( .A1(n485), .A2(n511), .ZN(n488) );
  XNOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n496) );
  NAND2_X1 U548 ( .A1(n540), .A2(n496), .ZN(n490) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n513), .A2(n496), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n493) );
  NAND2_X1 U555 ( .A1(n496), .A2(n522), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U558 ( .A1(n496), .A2(n518), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n501) );
  INV_X1 U561 ( .A(n498), .ZN(n558) );
  NOR2_X1 U562 ( .A1(n543), .A2(n558), .ZN(n510) );
  AND2_X1 U563 ( .A1(n499), .A2(n510), .ZN(n505) );
  NAND2_X1 U564 ( .A1(n505), .A2(n540), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n513), .A2(n505), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n505), .A2(n522), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U572 ( .A1(n505), .A2(n518), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT106), .Z(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  AND2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n540), .A2(n519), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n513), .A2(n519), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U582 ( .A1(n519), .A2(n522), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n517), .ZN(G1338GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(KEYINPUT44), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NAND2_X1 U588 ( .A1(n522), .A2(n539), .ZN(n523) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U590 ( .A(KEYINPUT113), .B(n525), .Z(n531) );
  NAND2_X1 U591 ( .A1(n531), .A2(n543), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U594 ( .A1(n531), .A2(n498), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n530) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n533) );
  INV_X1 U599 ( .A(n531), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n563), .A2(n534), .ZN(n532) );
  XOR2_X1 U601 ( .A(n533), .B(n532), .Z(G1342GAT) );
  NOR2_X1 U602 ( .A1(n534), .A2(n551), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n536) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT117), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n543), .A2(n553), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U612 ( .A1(n553), .A2(n498), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT118), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n553), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  XOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT119), .Z(n555) );
  INV_X1 U619 ( .A(n551), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U622 ( .A1(n567), .A2(n562), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  NOR2_X1 U625 ( .A1(n562), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n561), .ZN(G1349GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U630 ( .A(G183GAT), .B(n564), .Z(G1350GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n578) );
  NOR2_X1 U632 ( .A1(n567), .A2(n578), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n578), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(n576), .Z(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

