

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n650), .A2(n649), .ZN(n652) );
  NOR2_X1 U556 ( .A1(n550), .A2(n549), .ZN(G160) );
  XOR2_X1 U557 ( .A(G543), .B(KEYINPUT0), .Z(n521) );
  AND2_X1 U558 ( .A1(n745), .A2(n744), .ZN(n522) );
  AND2_X1 U559 ( .A1(n748), .A2(n747), .ZN(n523) );
  INV_X1 U560 ( .A(KEYINPUT27), .ZN(n653) );
  XNOR2_X1 U561 ( .A(n653), .B(KEYINPUT95), .ZN(n654) );
  XNOR2_X1 U562 ( .A(n655), .B(n654), .ZN(n657) );
  INV_X1 U563 ( .A(KEYINPUT31), .ZN(n651) );
  AND2_X1 U564 ( .A1(n643), .A2(n744), .ZN(n722) );
  NOR2_X1 U565 ( .A1(n746), .A2(n522), .ZN(n747) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n545) );
  NOR2_X1 U567 ( .A1(G651), .A2(n571), .ZN(n805) );
  INV_X1 U568 ( .A(KEYINPUT78), .ZN(n538) );
  NOR2_X1 U569 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U570 ( .A(n752), .B(KEYINPUT104), .ZN(n753) );
  XNOR2_X1 U571 ( .A(n538), .B(KEYINPUT8), .ZN(n539) );
  XNOR2_X1 U572 ( .A(G168), .B(n539), .ZN(G286) );
  NOR2_X1 U573 ( .A1(n558), .A2(n557), .ZN(G164) );
  INV_X1 U574 ( .A(G651), .ZN(n528) );
  NOR2_X1 U575 ( .A1(G543), .A2(n528), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n524), .Z(n798) );
  NAND2_X1 U577 ( .A1(G63), .A2(n798), .ZN(n526) );
  XNOR2_X1 U578 ( .A(KEYINPUT66), .B(n521), .ZN(n571) );
  NAND2_X1 U579 ( .A1(G51), .A2(n805), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U581 ( .A(KEYINPUT6), .B(n527), .ZN(n535) );
  NOR2_X2 U582 ( .A1(n571), .A2(n528), .ZN(n797) );
  NAND2_X1 U583 ( .A1(n797), .A2(G76), .ZN(n529) );
  XNOR2_X1 U584 ( .A(n529), .B(KEYINPUT76), .ZN(n532) );
  NOR2_X1 U585 ( .A1(G543), .A2(G651), .ZN(n801) );
  NAND2_X1 U586 ( .A1(n801), .A2(G89), .ZN(n530) );
  XNOR2_X1 U587 ( .A(KEYINPUT4), .B(n530), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U589 ( .A(n533), .B(KEYINPUT5), .Z(n534) );
  XOR2_X1 U590 ( .A(KEYINPUT7), .B(n536), .Z(n537) );
  XOR2_X1 U591 ( .A(KEYINPUT77), .B(n537), .Z(G168) );
  INV_X1 U592 ( .A(G2105), .ZN(n546) );
  INV_X1 U593 ( .A(G2104), .ZN(n540) );
  NOR2_X1 U594 ( .A1(n546), .A2(n540), .ZN(n896) );
  NAND2_X1 U595 ( .A1(n896), .A2(G113), .ZN(n544) );
  NOR2_X1 U596 ( .A1(n540), .A2(G2105), .ZN(n541) );
  XNOR2_X2 U597 ( .A(n541), .B(KEYINPUT64), .ZN(n892) );
  NAND2_X1 U598 ( .A1(n892), .A2(G101), .ZN(n542) );
  XOR2_X1 U599 ( .A(KEYINPUT23), .B(n542), .Z(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n550) );
  XOR2_X2 U601 ( .A(KEYINPUT17), .B(n545), .Z(n891) );
  NAND2_X1 U602 ( .A1(G137), .A2(n891), .ZN(n548) );
  NOR2_X1 U603 ( .A1(G2104), .A2(n546), .ZN(n895) );
  NAND2_X1 U604 ( .A1(G125), .A2(n895), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n891), .A2(G138), .ZN(n551) );
  XNOR2_X1 U607 ( .A(KEYINPUT91), .B(n551), .ZN(n558) );
  NAND2_X1 U608 ( .A1(n892), .A2(G102), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(KEYINPUT90), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G114), .A2(n896), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G126), .A2(n895), .ZN(n553) );
  AND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G85), .A2(n801), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n559), .B(KEYINPUT65), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G60), .A2(n798), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G47), .A2(n805), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U619 ( .A(KEYINPUT67), .B(n562), .Z(n563) );
  NOR2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n797), .A2(G72), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(G290) );
  NAND2_X1 U623 ( .A1(G49), .A2(n805), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G74), .A2(G651), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U626 ( .A1(n798), .A2(n569), .ZN(n570) );
  XOR2_X1 U627 ( .A(KEYINPUT85), .B(n570), .Z(n573) );
  NAND2_X1 U628 ( .A1(G87), .A2(n571), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n573), .A2(n572), .ZN(G288) );
  NAND2_X1 U630 ( .A1(G73), .A2(n797), .ZN(n574) );
  XNOR2_X1 U631 ( .A(n574), .B(KEYINPUT2), .ZN(n581) );
  NAND2_X1 U632 ( .A1(G61), .A2(n798), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G48), .A2(n805), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n801), .A2(G86), .ZN(n577) );
  XOR2_X1 U636 ( .A(KEYINPUT86), .B(n577), .Z(n578) );
  NOR2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U639 ( .A1(G64), .A2(n798), .ZN(n582) );
  XOR2_X1 U640 ( .A(KEYINPUT68), .B(n582), .Z(n589) );
  NAND2_X1 U641 ( .A1(G90), .A2(n801), .ZN(n584) );
  NAND2_X1 U642 ( .A1(G77), .A2(n797), .ZN(n583) );
  NAND2_X1 U643 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U644 ( .A(n585), .B(KEYINPUT9), .ZN(n587) );
  NAND2_X1 U645 ( .A1(G52), .A2(n805), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U647 ( .A1(n589), .A2(n588), .ZN(G171) );
  NAND2_X1 U648 ( .A1(G88), .A2(n801), .ZN(n591) );
  NAND2_X1 U649 ( .A1(G75), .A2(n797), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U651 ( .A1(n805), .A2(G50), .ZN(n593) );
  NAND2_X1 U652 ( .A1(n798), .A2(G62), .ZN(n592) );
  NAND2_X1 U653 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U654 ( .A1(n595), .A2(n594), .ZN(G166) );
  INV_X1 U655 ( .A(G166), .ZN(G303) );
  NOR2_X1 U656 ( .A1(G164), .A2(G1384), .ZN(n639) );
  NAND2_X1 U657 ( .A1(G160), .A2(G40), .ZN(n637) );
  NOR2_X1 U658 ( .A1(n639), .A2(n637), .ZN(n634) );
  NAND2_X1 U659 ( .A1(G117), .A2(n896), .ZN(n597) );
  NAND2_X1 U660 ( .A1(G129), .A2(n895), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G105), .A2(n892), .ZN(n598) );
  XOR2_X1 U663 ( .A(KEYINPUT38), .B(n598), .Z(n599) );
  NOR2_X1 U664 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U665 ( .A(n601), .B(KEYINPUT92), .ZN(n603) );
  NAND2_X1 U666 ( .A1(G141), .A2(n891), .ZN(n602) );
  NAND2_X1 U667 ( .A1(n603), .A2(n602), .ZN(n906) );
  NOR2_X1 U668 ( .A1(G1996), .A2(n906), .ZN(n922) );
  AND2_X1 U669 ( .A1(n906), .A2(G1996), .ZN(n611) );
  NAND2_X1 U670 ( .A1(G107), .A2(n896), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G119), .A2(n895), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U673 ( .A1(G131), .A2(n891), .ZN(n607) );
  NAND2_X1 U674 ( .A1(G95), .A2(n892), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n608) );
  OR2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n883) );
  AND2_X1 U677 ( .A1(n883), .A2(G1991), .ZN(n610) );
  NOR2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n925) );
  INV_X1 U679 ( .A(n634), .ZN(n612) );
  NOR2_X1 U680 ( .A1(n925), .A2(n612), .ZN(n632) );
  NOR2_X1 U681 ( .A1(G1986), .A2(G290), .ZN(n613) );
  NOR2_X1 U682 ( .A1(G1991), .A2(n883), .ZN(n934) );
  NOR2_X1 U683 ( .A1(n613), .A2(n934), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n614), .B(KEYINPUT102), .ZN(n615) );
  NOR2_X1 U685 ( .A1(n632), .A2(n615), .ZN(n616) );
  NOR2_X1 U686 ( .A1(n922), .A2(n616), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(KEYINPUT39), .ZN(n627) );
  NAND2_X1 U688 ( .A1(G116), .A2(n896), .ZN(n619) );
  NAND2_X1 U689 ( .A1(G128), .A2(n895), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT35), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G140), .A2(n891), .ZN(n622) );
  NAND2_X1 U693 ( .A1(G104), .A2(n892), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U695 ( .A(KEYINPUT34), .B(n623), .Z(n624) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U697 ( .A(n626), .B(KEYINPUT36), .Z(n887) );
  XNOR2_X1 U698 ( .A(G2067), .B(KEYINPUT37), .ZN(n628) );
  OR2_X1 U699 ( .A1(n887), .A2(n628), .ZN(n937) );
  NAND2_X1 U700 ( .A1(n627), .A2(n937), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n887), .A2(n628), .ZN(n935) );
  NAND2_X1 U702 ( .A1(n629), .A2(n935), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n634), .A2(n630), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n631), .B(KEYINPUT103), .ZN(n751) );
  INV_X1 U705 ( .A(n632), .ZN(n636) );
  XOR2_X1 U706 ( .A(G1986), .B(G290), .Z(n987) );
  NAND2_X1 U707 ( .A1(n987), .A2(n937), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n749) );
  NOR2_X1 U710 ( .A1(G1976), .A2(G288), .ZN(n729) );
  AND2_X1 U711 ( .A1(n729), .A2(KEYINPUT33), .ZN(n641) );
  INV_X1 U712 ( .A(n637), .ZN(n638) );
  NAND2_X2 U713 ( .A1(n639), .A2(n638), .ZN(n710) );
  NAND2_X1 U714 ( .A1(n710), .A2(G8), .ZN(n640) );
  XNOR2_X2 U715 ( .A(n640), .B(KEYINPUT93), .ZN(n744) );
  NAND2_X1 U716 ( .A1(n641), .A2(n744), .ZN(n736) );
  XOR2_X1 U717 ( .A(G1981), .B(KEYINPUT101), .Z(n642) );
  XNOR2_X1 U718 ( .A(G305), .B(n642), .ZN(n974) );
  INV_X1 U719 ( .A(n744), .ZN(n732) );
  INV_X1 U720 ( .A(G1966), .ZN(n643) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n710), .ZN(n719) );
  NOR2_X1 U722 ( .A1(n722), .A2(n719), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G8), .A2(n644), .ZN(n645) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n645), .ZN(n646) );
  NOR2_X1 U725 ( .A1(G168), .A2(n646), .ZN(n650) );
  INV_X1 U726 ( .A(G1961), .ZN(n996) );
  NAND2_X1 U727 ( .A1(n710), .A2(n996), .ZN(n648) );
  INV_X1 U728 ( .A(n710), .ZN(n676) );
  XNOR2_X1 U729 ( .A(G2078), .B(KEYINPUT25), .ZN(n952) );
  NAND2_X1 U730 ( .A1(n676), .A2(n952), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n705) );
  NOR2_X1 U732 ( .A1(G171), .A2(n705), .ZN(n649) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(n709) );
  NAND2_X1 U734 ( .A1(G2072), .A2(n676), .ZN(n655) );
  AND2_X1 U735 ( .A1(n710), .A2(G1956), .ZN(n656) );
  NOR2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n666) );
  NAND2_X1 U737 ( .A1(G65), .A2(n798), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G53), .A2(n805), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U740 ( .A1(G91), .A2(n801), .ZN(n661) );
  NAND2_X1 U741 ( .A1(G78), .A2(n797), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U743 ( .A1(n663), .A2(n662), .ZN(n920) );
  NOR2_X1 U744 ( .A1(n666), .A2(n920), .ZN(n665) );
  XOR2_X1 U745 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n664) );
  XNOR2_X1 U746 ( .A(n665), .B(n664), .ZN(n702) );
  NAND2_X1 U747 ( .A1(n666), .A2(n920), .ZN(n700) );
  NAND2_X1 U748 ( .A1(G79), .A2(n797), .ZN(n668) );
  NAND2_X1 U749 ( .A1(G54), .A2(n805), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n668), .A2(n667), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G92), .A2(n801), .ZN(n670) );
  NAND2_X1 U752 ( .A1(G66), .A2(n798), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U754 ( .A(n671), .B(KEYINPUT73), .Z(n672) );
  NOR2_X1 U755 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U756 ( .A(KEYINPUT15), .B(n674), .ZN(n675) );
  XNOR2_X1 U757 ( .A(KEYINPUT74), .B(n675), .ZN(n978) );
  NAND2_X1 U758 ( .A1(G1348), .A2(n710), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n676), .A2(G2067), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n678), .A2(n677), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n978), .A2(n696), .ZN(n680) );
  NAND2_X1 U762 ( .A1(G1341), .A2(n710), .ZN(n679) );
  NAND2_X1 U763 ( .A1(n680), .A2(n679), .ZN(n695) );
  NAND2_X1 U764 ( .A1(G43), .A2(n805), .ZN(n691) );
  NAND2_X1 U765 ( .A1(n798), .A2(G56), .ZN(n681) );
  XNOR2_X1 U766 ( .A(KEYINPUT14), .B(n681), .ZN(n688) );
  NAND2_X1 U767 ( .A1(G81), .A2(n801), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n682), .B(KEYINPUT12), .ZN(n683) );
  XNOR2_X1 U769 ( .A(n683), .B(KEYINPUT70), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G68), .A2(n797), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U772 ( .A(KEYINPUT13), .B(n686), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U774 ( .A(KEYINPUT71), .B(n689), .ZN(n690) );
  NAND2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n779) );
  INV_X1 U776 ( .A(n779), .ZN(n972) );
  XNOR2_X1 U777 ( .A(G1996), .B(KEYINPUT97), .ZN(n951) );
  NOR2_X1 U778 ( .A1(n710), .A2(n951), .ZN(n692) );
  XOR2_X1 U779 ( .A(KEYINPUT26), .B(n692), .Z(n693) );
  NAND2_X1 U780 ( .A1(n972), .A2(n693), .ZN(n694) );
  NOR2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n698) );
  NOR2_X1 U782 ( .A1(n978), .A2(n696), .ZN(n697) );
  NOR2_X1 U783 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U784 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U785 ( .A1(n702), .A2(n701), .ZN(n704) );
  XOR2_X1 U786 ( .A(KEYINPUT98), .B(KEYINPUT29), .Z(n703) );
  XNOR2_X1 U787 ( .A(n704), .B(n703), .ZN(n707) );
  NAND2_X1 U788 ( .A1(n705), .A2(G171), .ZN(n706) );
  NAND2_X1 U789 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U790 ( .A1(n709), .A2(n708), .ZN(n720) );
  NAND2_X1 U791 ( .A1(n720), .A2(G286), .ZN(n716) );
  NOR2_X1 U792 ( .A1(G1971), .A2(n732), .ZN(n712) );
  NOR2_X1 U793 ( .A1(G2090), .A2(n710), .ZN(n711) );
  NOR2_X1 U794 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U795 ( .A1(n713), .A2(G303), .ZN(n714) );
  XOR2_X1 U796 ( .A(KEYINPUT99), .B(n714), .Z(n715) );
  NAND2_X1 U797 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U798 ( .A1(n717), .A2(G8), .ZN(n718) );
  XNOR2_X1 U799 ( .A(n718), .B(KEYINPUT32), .ZN(n726) );
  NAND2_X1 U800 ( .A1(G8), .A2(n719), .ZN(n724) );
  INV_X1 U801 ( .A(n720), .ZN(n721) );
  NOR2_X1 U802 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U803 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U804 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U805 ( .A(n727), .B(KEYINPUT100), .ZN(n737) );
  NOR2_X1 U806 ( .A1(G1971), .A2(G303), .ZN(n728) );
  NOR2_X1 U807 ( .A1(n729), .A2(n728), .ZN(n988) );
  NAND2_X1 U808 ( .A1(n737), .A2(n988), .ZN(n730) );
  NAND2_X1 U809 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NAND2_X1 U810 ( .A1(n730), .A2(n982), .ZN(n731) );
  NOR2_X1 U811 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U812 ( .A1(KEYINPUT33), .A2(n733), .ZN(n734) );
  NOR2_X1 U813 ( .A1(n974), .A2(n734), .ZN(n735) );
  NAND2_X1 U814 ( .A1(n736), .A2(n735), .ZN(n748) );
  INV_X1 U815 ( .A(n737), .ZN(n740) );
  NAND2_X1 U816 ( .A1(G166), .A2(G8), .ZN(n738) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U818 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U819 ( .A1(n744), .A2(n741), .ZN(n746) );
  NOR2_X1 U820 ( .A1(G1981), .A2(G305), .ZN(n742) );
  XNOR2_X1 U821 ( .A(n742), .B(KEYINPUT94), .ZN(n743) );
  XNOR2_X1 U822 ( .A(n743), .B(KEYINPUT24), .ZN(n745) );
  NOR2_X1 U823 ( .A1(n749), .A2(n523), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n754) );
  INV_X1 U825 ( .A(KEYINPUT40), .ZN(n752) );
  XNOR2_X1 U826 ( .A(n754), .B(n753), .ZN(G329) );
  XOR2_X1 U827 ( .A(G2435), .B(G2454), .Z(n756) );
  XNOR2_X1 U828 ( .A(G2430), .B(G2438), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n756), .B(n755), .ZN(n763) );
  XOR2_X1 U830 ( .A(G2446), .B(KEYINPUT105), .Z(n758) );
  XNOR2_X1 U831 ( .A(G2451), .B(G2443), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n758), .B(n757), .ZN(n759) );
  XOR2_X1 U833 ( .A(n759), .B(G2427), .Z(n761) );
  XNOR2_X1 U834 ( .A(G1348), .B(G1341), .ZN(n760) );
  XNOR2_X1 U835 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U836 ( .A(n763), .B(n762), .ZN(n764) );
  AND2_X1 U837 ( .A1(n764), .A2(G14), .ZN(G401) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  INV_X1 U840 ( .A(G132), .ZN(G219) );
  INV_X1 U841 ( .A(G82), .ZN(G220) );
  XOR2_X1 U842 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n766) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U844 ( .A(n766), .B(n765), .ZN(G223) );
  INV_X1 U845 ( .A(G223), .ZN(n835) );
  NAND2_X1 U846 ( .A1(n835), .A2(G567), .ZN(n767) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  NAND2_X1 U848 ( .A1(G860), .A2(n972), .ZN(n768) );
  XNOR2_X1 U849 ( .A(n768), .B(KEYINPUT72), .ZN(G153) );
  INV_X1 U850 ( .A(G171), .ZN(G301) );
  INV_X1 U851 ( .A(n978), .ZN(n792) );
  NOR2_X1 U852 ( .A1(G868), .A2(n792), .ZN(n769) );
  XNOR2_X1 U853 ( .A(n769), .B(KEYINPUT75), .ZN(n771) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n771), .A2(n770), .ZN(G284) );
  INV_X1 U856 ( .A(G868), .ZN(n818) );
  NAND2_X1 U857 ( .A1(n920), .A2(n818), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT79), .ZN(n774) );
  NOR2_X1 U859 ( .A1(G286), .A2(n818), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(G297) );
  INV_X1 U861 ( .A(G860), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n775), .A2(G559), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n776), .A2(n792), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U865 ( .A1(G868), .A2(n792), .ZN(n778) );
  NOR2_X1 U866 ( .A1(G559), .A2(n778), .ZN(n781) );
  NOR2_X1 U867 ( .A1(G868), .A2(n779), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U869 ( .A1(G111), .A2(n896), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G135), .A2(n891), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n789) );
  NAND2_X1 U872 ( .A1(n892), .A2(G99), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n784), .B(KEYINPUT80), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G123), .A2(n895), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n785), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n933) );
  XNOR2_X1 U878 ( .A(n933), .B(G2096), .ZN(n791) );
  INV_X1 U879 ( .A(G2100), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(G156) );
  XOR2_X1 U881 ( .A(n972), .B(KEYINPUT81), .Z(n794) );
  NAND2_X1 U882 ( .A1(G559), .A2(n792), .ZN(n793) );
  XNOR2_X1 U883 ( .A(n794), .B(n793), .ZN(n815) );
  XOR2_X1 U884 ( .A(n815), .B(KEYINPUT82), .Z(n795) );
  NOR2_X1 U885 ( .A1(G860), .A2(n795), .ZN(n796) );
  XOR2_X1 U886 ( .A(KEYINPUT84), .B(n796), .Z(n808) );
  NAND2_X1 U887 ( .A1(G80), .A2(n797), .ZN(n800) );
  NAND2_X1 U888 ( .A1(G67), .A2(n798), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G93), .A2(n801), .ZN(n802) );
  XNOR2_X1 U891 ( .A(KEYINPUT83), .B(n802), .ZN(n803) );
  NOR2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n805), .A2(G55), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n819) );
  XNOR2_X1 U895 ( .A(n808), .B(n819), .ZN(G145) );
  XNOR2_X1 U896 ( .A(G166), .B(n819), .ZN(n813) );
  XOR2_X1 U897 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n809) );
  XNOR2_X1 U898 ( .A(G305), .B(n809), .ZN(n810) );
  XNOR2_X1 U899 ( .A(n920), .B(n810), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n811), .B(G290), .ZN(n812) );
  XNOR2_X1 U901 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n814), .B(G288), .ZN(n909) );
  XNOR2_X1 U903 ( .A(n815), .B(n909), .ZN(n816) );
  XNOR2_X1 U904 ( .A(KEYINPUT88), .B(n816), .ZN(n817) );
  NOR2_X1 U905 ( .A1(n818), .A2(n817), .ZN(n821) );
  NOR2_X1 U906 ( .A1(G868), .A2(n819), .ZN(n820) );
  NOR2_X1 U907 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U908 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U909 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n823), .ZN(n825) );
  XOR2_X1 U911 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n824) );
  XNOR2_X1 U912 ( .A(n825), .B(n824), .ZN(n826) );
  NAND2_X1 U913 ( .A1(G2072), .A2(n826), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n827) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U917 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U918 ( .A1(G96), .A2(n829), .ZN(n841) );
  NAND2_X1 U919 ( .A1(n841), .A2(G2106), .ZN(n833) );
  NAND2_X1 U920 ( .A1(G69), .A2(G120), .ZN(n830) );
  NOR2_X1 U921 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G108), .A2(n831), .ZN(n842) );
  NAND2_X1 U923 ( .A1(n842), .A2(G567), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n843) );
  NAND2_X1 U925 ( .A1(G483), .A2(G661), .ZN(n834) );
  NOR2_X1 U926 ( .A1(n843), .A2(n834), .ZN(n840) );
  NAND2_X1 U927 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n835), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT106), .B(n836), .Z(n837) );
  NAND2_X1 U931 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT107), .B(n838), .Z(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  INV_X1 U941 ( .A(n843), .ZN(G319) );
  XOR2_X1 U942 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2678), .B(KEYINPUT43), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(KEYINPUT42), .B(G2067), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2090), .B(G2072), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2096), .B(G2100), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U951 ( .A(G2078), .B(G2084), .Z(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G227) );
  XNOR2_X1 U953 ( .A(G1956), .B(KEYINPUT110), .ZN(n863) );
  XOR2_X1 U954 ( .A(G1986), .B(G1976), .Z(n855) );
  XNOR2_X1 U955 ( .A(G1961), .B(G1971), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U957 ( .A(G1981), .B(G1966), .Z(n857) );
  XNOR2_X1 U958 ( .A(G1991), .B(G1996), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U961 ( .A(G2474), .B(KEYINPUT41), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G124), .A2(n895), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n896), .A2(G112), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G136), .A2(n891), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G100), .A2(n892), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U971 ( .A1(n870), .A2(n869), .ZN(G162) );
  XOR2_X1 U972 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n872) );
  XNOR2_X1 U973 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(n873), .B(KEYINPUT112), .Z(n885) );
  NAND2_X1 U976 ( .A1(G118), .A2(n896), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G130), .A2(n895), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G142), .A2(n891), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G106), .A2(n892), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n878), .ZN(n879) );
  XNOR2_X1 U983 ( .A(KEYINPUT111), .B(n879), .ZN(n880) );
  NOR2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U985 ( .A(n883), .B(n882), .Z(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U987 ( .A(n886), .B(n933), .Z(n889) );
  XOR2_X1 U988 ( .A(G164), .B(n887), .Z(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U990 ( .A(n890), .B(G162), .Z(n905) );
  NAND2_X1 U991 ( .A1(G139), .A2(n891), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G103), .A2(n892), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n903) );
  XNOR2_X1 U994 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n901) );
  NAND2_X1 U995 ( .A1(n895), .A2(G127), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n896), .A2(G115), .ZN(n897) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(n897), .Z(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n927) );
  XNOR2_X1 U1001 ( .A(G160), .B(n927), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n907), .B(n906), .Z(n908) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n908), .ZN(G395) );
  XNOR2_X1 U1005 ( .A(G286), .B(n909), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(G171), .B(n978), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(n972), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n914) );
  XOR2_X1 U1011 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  XOR2_X1 U1015 ( .A(KEYINPUT117), .B(n917), .Z(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  INV_X1 U1019 ( .A(n920), .ZN(G299) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n923), .Z(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n932) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT118), .B(n926), .ZN(n929) );
  XOR2_X1 U1026 ( .A(G2072), .B(n927), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT50), .B(n930), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n942) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(G160), .B(G2084), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(KEYINPUT119), .B(n943), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n944), .ZN(n946) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(KEYINPUT120), .B(n948), .ZN(n1027) );
  XOR2_X1 U1042 ( .A(G2084), .B(G34), .Z(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT54), .B(n949), .ZN(n966) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n964) );
  XOR2_X1 U1045 ( .A(G2072), .B(G33), .Z(n950) );
  NAND2_X1 U1046 ( .A1(n950), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1047 ( .A(n951), .B(G32), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n952), .B(G27), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT121), .B(n955), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(G1991), .B(G25), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(G26), .B(G2067), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(n967), .B(KEYINPUT122), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n968), .B(KEYINPUT55), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(G29), .A2(n969), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(KEYINPUT123), .B(n970), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n971), .A2(G11), .ZN(n1025) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XOR2_X1 U1065 ( .A(n972), .B(G1341), .Z(n977) );
  XOR2_X1 U1066 ( .A(G1966), .B(G168), .Z(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(KEYINPUT57), .B(n975), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n993) );
  XNOR2_X1 U1070 ( .A(G301), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(n978), .B(G1348), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n986) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1956), .B(G299), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(n991), .B(KEYINPUT124), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n1023) );
  INV_X1 U1083 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1084 ( .A(G5), .B(n996), .ZN(n1009) );
  XNOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n997), .B(G4), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G20), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G6), .B(G1981), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT125), .B(G1341), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(G19), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1010), .ZN(n1018) );
  XOR2_X1 U1099 ( .A(G1976), .B(G23), .Z(n1014) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G24), .B(G1986), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

