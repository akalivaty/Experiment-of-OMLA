

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G2105), .A2(n522), .ZN(n976) );
  XNOR2_X1 U551 ( .A(n784), .B(n681), .ZN(n682) );
  OR2_X1 U552 ( .A1(n694), .A2(n971), .ZN(n693) );
  OR2_X1 U553 ( .A1(n720), .A2(n683), .ZN(n685) );
  INV_X1 U554 ( .A(KEYINPUT102), .ZN(n686) );
  XNOR2_X1 U555 ( .A(n687), .B(n686), .ZN(n694) );
  INV_X1 U556 ( .A(KEYINPUT100), .ZN(n681) );
  NOR2_X1 U557 ( .A1(n747), .A2(n746), .ZN(n802) );
  NAND2_X2 U558 ( .A1(n682), .A2(n785), .ZN(n720) );
  NOR2_X1 U559 ( .A1(n792), .A2(n791), .ZN(n795) );
  NOR2_X1 U560 ( .A1(G651), .A2(n629), .ZN(n641) );
  NOR2_X2 U561 ( .A1(n527), .A2(n526), .ZN(G160) );
  INV_X1 U562 ( .A(G2104), .ZN(n522) );
  INV_X1 U563 ( .A(G2105), .ZN(n517) );
  NOR2_X1 U564 ( .A1(n522), .A2(n517), .ZN(n981) );
  NAND2_X1 U565 ( .A1(G113), .A2(n981), .ZN(n519) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n517), .ZN(n982) );
  NAND2_X1 U567 ( .A1(G125), .A2(n982), .ZN(n518) );
  NAND2_X1 U568 ( .A1(n519), .A2(n518), .ZN(n527) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n520), .Z(n977) );
  NAND2_X1 U571 ( .A1(G137), .A2(n977), .ZN(n521) );
  XNOR2_X1 U572 ( .A(n521), .B(KEYINPUT64), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G101), .A2(n976), .ZN(n523) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X1 U576 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U577 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n529) );
  NAND2_X1 U578 ( .A1(G123), .A2(n982), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n529), .B(n528), .ZN(n536) );
  NAND2_X1 U580 ( .A1(G99), .A2(n976), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G135), .A2(n977), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n981), .A2(G111), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT80), .B(n532), .Z(n533) );
  NOR2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n991) );
  XNOR2_X1 U587 ( .A(G2096), .B(n991), .ZN(n537) );
  OR2_X1 U588 ( .A1(G2100), .A2(n537), .ZN(G156) );
  NOR2_X1 U589 ( .A1(G543), .A2(G651), .ZN(n632) );
  NAND2_X1 U590 ( .A1(G90), .A2(n632), .ZN(n539) );
  XOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .Z(n629) );
  INV_X1 U592 ( .A(G651), .ZN(n541) );
  NOR2_X1 U593 ( .A1(n629), .A2(n541), .ZN(n636) );
  NAND2_X1 U594 ( .A1(G77), .A2(n636), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n540), .B(KEYINPUT9), .ZN(n544) );
  NOR2_X1 U597 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n542), .Z(n633) );
  NAND2_X1 U599 ( .A1(G64), .A2(n633), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G52), .A2(n641), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT67), .B(n545), .ZN(n546) );
  NOR2_X1 U603 ( .A1(n547), .A2(n546), .ZN(G171) );
  NAND2_X1 U604 ( .A1(n632), .A2(G89), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G76), .A2(n636), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT5), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n641), .A2(G51), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT76), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G63), .A2(n633), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n558), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n561) );
  XNOR2_X1 U620 ( .A(G223), .B(KEYINPUT71), .ZN(n823) );
  NAND2_X1 U621 ( .A1(G567), .A2(n823), .ZN(n560) );
  XNOR2_X1 U622 ( .A(n561), .B(n560), .ZN(G234) );
  NAND2_X1 U623 ( .A1(G56), .A2(n633), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT14), .B(n562), .Z(n568) );
  NAND2_X1 U625 ( .A1(n632), .A2(G81), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G68), .A2(n636), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n566), .Z(n567) );
  NOR2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n641), .A2(G43), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n970) );
  XNOR2_X1 U633 ( .A(G860), .B(KEYINPUT73), .ZN(n593) );
  OR2_X1 U634 ( .A1(n970), .A2(n593), .ZN(G153) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G92), .A2(n632), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G66), .A2(n633), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT74), .B(n573), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G79), .A2(n636), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G54), .A2(n641), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT15), .B(n578), .Z(n971) );
  NOR2_X1 U645 ( .A1(n971), .A2(G868), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(KEYINPUT75), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U649 ( .A1(G91), .A2(n632), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G78), .A2(n636), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U652 ( .A(KEYINPUT68), .B(n584), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G65), .A2(n633), .ZN(n585) );
  XNOR2_X1 U654 ( .A(KEYINPUT69), .B(n585), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n641), .A2(G53), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(G299) );
  INV_X1 U658 ( .A(G299), .ZN(n703) );
  INV_X1 U659 ( .A(G868), .ZN(n644) );
  NAND2_X1 U660 ( .A1(n703), .A2(n644), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT77), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n644), .A2(G286), .ZN(n591) );
  NOR2_X1 U663 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U664 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n594), .A2(n971), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  AND2_X1 U667 ( .A1(n971), .A2(G868), .ZN(n596) );
  XOR2_X1 U668 ( .A(KEYINPUT78), .B(n596), .Z(n597) );
  NOR2_X1 U669 ( .A1(G559), .A2(n597), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G868), .A2(n970), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G559), .A2(n971), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT81), .B(n600), .Z(n601) );
  XNOR2_X1 U674 ( .A(n970), .B(n601), .ZN(n654) );
  NOR2_X1 U675 ( .A1(n654), .A2(G860), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G55), .A2(n641), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G67), .A2(n633), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U679 ( .A(KEYINPUT82), .B(n604), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G93), .A2(n632), .ZN(n606) );
  NAND2_X1 U681 ( .A1(G80), .A2(n636), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n645) );
  XNOR2_X1 U684 ( .A(n609), .B(n645), .ZN(G145) );
  NAND2_X1 U685 ( .A1(n636), .A2(G75), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n610), .B(KEYINPUT84), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G88), .A2(n632), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U689 ( .A(KEYINPUT85), .B(n613), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n641), .A2(G50), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G62), .A2(n633), .ZN(n614) );
  AND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(G303) );
  INV_X1 U694 ( .A(G303), .ZN(G166) );
  NAND2_X1 U695 ( .A1(G47), .A2(n641), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT66), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G85), .A2(n632), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G60), .A2(n633), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G72), .A2(n636), .ZN(n621) );
  XNOR2_X1 U701 ( .A(KEYINPUT65), .B(n621), .ZN(n622) );
  NOR2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(G290) );
  NAND2_X1 U704 ( .A1(G49), .A2(n641), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U707 ( .A1(n633), .A2(n628), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G86), .A2(n632), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G61), .A2(n633), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G73), .A2(n636), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n637), .B(KEYINPUT83), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(KEYINPUT2), .ZN(n639) );
  NOR2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n641), .A2(G48), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U719 ( .A1(n644), .A2(n645), .ZN(n657) );
  XOR2_X1 U720 ( .A(n645), .B(G166), .Z(n653) );
  XOR2_X1 U721 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n646) );
  XNOR2_X1 U722 ( .A(G288), .B(n646), .ZN(n647) );
  XOR2_X1 U723 ( .A(n647), .B(KEYINPUT86), .Z(n649) );
  XOR2_X1 U724 ( .A(G299), .B(KEYINPUT19), .Z(n648) );
  XNOR2_X1 U725 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U726 ( .A(n650), .B(G305), .Z(n651) );
  XNOR2_X1 U727 ( .A(G290), .B(n651), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n653), .B(n652), .ZN(n969) );
  XNOR2_X1 U729 ( .A(n969), .B(n654), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n655), .A2(G868), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(KEYINPUT89), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U735 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U736 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XOR2_X1 U738 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U740 ( .A1(G108), .A2(G120), .ZN(n663) );
  NOR2_X1 U741 ( .A1(G237), .A2(n663), .ZN(n664) );
  NAND2_X1 U742 ( .A1(G69), .A2(n664), .ZN(n945) );
  NAND2_X1 U743 ( .A1(G567), .A2(n945), .ZN(n665) );
  XNOR2_X1 U744 ( .A(KEYINPUT92), .B(n665), .ZN(n672) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n667) );
  NAND2_X1 U746 ( .A1(G132), .A2(G82), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT90), .ZN(n669) );
  NOR2_X1 U749 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G96), .A2(n670), .ZN(n946) );
  NAND2_X1 U751 ( .A1(G2106), .A2(n946), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n672), .A2(n671), .ZN(n947) );
  NAND2_X1 U753 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U754 ( .A1(n947), .A2(n673), .ZN(n826) );
  NAND2_X1 U755 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U756 ( .A1(G102), .A2(n976), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G138), .A2(n977), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U759 ( .A1(G114), .A2(n981), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G126), .A2(n982), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U762 ( .A1(n679), .A2(n678), .ZN(G164) );
  NOR2_X1 U763 ( .A1(G1971), .A2(G303), .ZN(n680) );
  XOR2_X1 U764 ( .A(n680), .B(KEYINPUT106), .Z(n749) );
  NOR2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n874) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n784) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n785) );
  INV_X1 U768 ( .A(G2067), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G1348), .A2(n720), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n687) );
  INV_X1 U771 ( .A(G1996), .ZN(n951) );
  NOR2_X1 U772 ( .A1(n720), .A2(n951), .ZN(n688) );
  XOR2_X1 U773 ( .A(n688), .B(KEYINPUT26), .Z(n690) );
  NAND2_X1 U774 ( .A1(n720), .A2(G1341), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U776 ( .A1(n970), .A2(n691), .ZN(n692) );
  NAND2_X1 U777 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U778 ( .A1(n694), .A2(n971), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U780 ( .A(n697), .B(KEYINPUT103), .ZN(n702) );
  INV_X1 U781 ( .A(n720), .ZN(n710) );
  NAND2_X1 U782 ( .A1(n710), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U783 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U784 ( .A(G1956), .ZN(n948) );
  NOR2_X1 U785 ( .A1(n948), .A2(n710), .ZN(n699) );
  NOR2_X1 U786 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n707) );
  NOR2_X1 U789 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U790 ( .A(n705), .B(KEYINPUT28), .Z(n706) );
  NAND2_X1 U791 ( .A1(n707), .A2(n706), .ZN(n709) );
  INV_X1 U792 ( .A(KEYINPUT29), .ZN(n708) );
  XNOR2_X1 U793 ( .A(n709), .B(n708), .ZN(n737) );
  XNOR2_X1 U794 ( .A(G1961), .B(KEYINPUT101), .ZN(n920) );
  NAND2_X1 U795 ( .A1(n720), .A2(n920), .ZN(n712) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n898) );
  NAND2_X1 U797 ( .A1(n710), .A2(n898), .ZN(n711) );
  NAND2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U799 ( .A1(n716), .A2(G171), .ZN(n735) );
  NAND2_X1 U800 ( .A1(n737), .A2(n735), .ZN(n726) );
  NAND2_X1 U801 ( .A1(G8), .A2(n720), .ZN(n799) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n799), .ZN(n738) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n720), .ZN(n742) );
  NOR2_X1 U804 ( .A1(n738), .A2(n742), .ZN(n713) );
  NAND2_X1 U805 ( .A1(G8), .A2(n713), .ZN(n714) );
  XNOR2_X1 U806 ( .A(KEYINPUT30), .B(n714), .ZN(n715) );
  NOR2_X1 U807 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U808 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U810 ( .A(n719), .B(KEYINPUT31), .Z(n739) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n799), .ZN(n722) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n723), .A2(G303), .ZN(n724) );
  XOR2_X1 U815 ( .A(KEYINPUT105), .B(n724), .Z(n727) );
  AND2_X1 U816 ( .A1(n739), .A2(n727), .ZN(n725) );
  NAND2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n731) );
  INV_X1 U818 ( .A(n727), .ZN(n728) );
  OR2_X1 U819 ( .A1(n728), .A2(G286), .ZN(n729) );
  AND2_X1 U820 ( .A1(n729), .A2(G8), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n733) );
  INV_X1 U822 ( .A(KEYINPUT32), .ZN(n732) );
  XNOR2_X1 U823 ( .A(n733), .B(n732), .ZN(n747) );
  INV_X1 U824 ( .A(n738), .ZN(n734) );
  AND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n741) );
  OR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n744) );
  NAND2_X1 U829 ( .A1(G8), .A2(n742), .ZN(n743) );
  NAND2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U831 ( .A(KEYINPUT104), .B(n745), .Z(n746) );
  NOR2_X1 U832 ( .A1(n874), .A2(n802), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n875) );
  NAND2_X1 U835 ( .A1(n750), .A2(n875), .ZN(n751) );
  XOR2_X1 U836 ( .A(KEYINPUT107), .B(n751), .Z(n792) );
  XOR2_X1 U837 ( .A(G1981), .B(G305), .Z(n870) );
  NAND2_X1 U838 ( .A1(n981), .A2(G117), .ZN(n752) );
  XOR2_X1 U839 ( .A(KEYINPUT97), .B(n752), .Z(n754) );
  NAND2_X1 U840 ( .A1(n982), .A2(G129), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U842 ( .A(KEYINPUT98), .B(n755), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n976), .A2(G105), .ZN(n756) );
  XOR2_X1 U844 ( .A(KEYINPUT38), .B(n756), .Z(n757) );
  NOR2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n977), .A2(G141), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U848 ( .A(KEYINPUT99), .B(n761), .Z(n1002) );
  NAND2_X1 U849 ( .A1(G1996), .A2(n1002), .ZN(n770) );
  NAND2_X1 U850 ( .A1(G95), .A2(n976), .ZN(n763) );
  NAND2_X1 U851 ( .A1(G119), .A2(n982), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n981), .A2(G107), .ZN(n764) );
  XOR2_X1 U854 ( .A(KEYINPUT96), .B(n764), .Z(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n977), .A2(G131), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n990) );
  NAND2_X1 U858 ( .A1(G1991), .A2(n990), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n835) );
  XNOR2_X1 U860 ( .A(G1986), .B(G290), .ZN(n873) );
  NOR2_X1 U861 ( .A1(n835), .A2(n873), .ZN(n783) );
  NAND2_X1 U862 ( .A1(n982), .A2(G128), .ZN(n771) );
  XNOR2_X1 U863 ( .A(KEYINPUT94), .B(n771), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n981), .A2(G116), .ZN(n772) );
  XOR2_X1 U865 ( .A(KEYINPUT95), .B(n772), .Z(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n775), .B(KEYINPUT35), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G104), .A2(n976), .ZN(n777) );
  NAND2_X1 U869 ( .A1(G140), .A2(n977), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U871 ( .A(KEYINPUT34), .B(n778), .Z(n779) );
  NAND2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U873 ( .A(n781), .B(KEYINPUT36), .Z(n1003) );
  XNOR2_X1 U874 ( .A(G2067), .B(KEYINPUT37), .ZN(n782) );
  XOR2_X1 U875 ( .A(n782), .B(KEYINPUT93), .Z(n814) );
  OR2_X1 U876 ( .A1(n1003), .A2(n814), .ZN(n852) );
  NAND2_X1 U877 ( .A1(n783), .A2(n852), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n816) );
  NAND2_X1 U879 ( .A1(n786), .A2(n816), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n870), .A2(n796), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n874), .A2(KEYINPUT33), .ZN(n787) );
  NOR2_X1 U882 ( .A1(n799), .A2(n787), .ZN(n788) );
  NOR2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n793) );
  INV_X1 U884 ( .A(n793), .ZN(n790) );
  OR2_X1 U885 ( .A1(n799), .A2(n790), .ZN(n791) );
  AND2_X1 U886 ( .A1(n793), .A2(KEYINPUT33), .ZN(n794) );
  NOR2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n821) );
  INV_X1 U888 ( .A(n796), .ZN(n808) );
  NOR2_X1 U889 ( .A1(G1981), .A2(G305), .ZN(n797) );
  XOR2_X1 U890 ( .A(n797), .B(KEYINPUT24), .Z(n798) );
  NOR2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n806) );
  INV_X1 U892 ( .A(n799), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G166), .A2(G8), .ZN(n800) );
  NOR2_X1 U894 ( .A1(G2090), .A2(n800), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n819) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n1002), .ZN(n856) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n990), .ZN(n851) );
  NOR2_X1 U902 ( .A1(n809), .A2(n851), .ZN(n810) );
  NOR2_X1 U903 ( .A1(n835), .A2(n810), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n856), .A2(n811), .ZN(n812) );
  XNOR2_X1 U905 ( .A(KEYINPUT39), .B(n812), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n813), .A2(n852), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n1003), .A2(n814), .ZN(n836) );
  NAND2_X1 U908 ( .A1(n815), .A2(n836), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  AND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U912 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(G188) );
  NAND2_X1 U919 ( .A1(G112), .A2(n981), .ZN(n833) );
  NAND2_X1 U920 ( .A1(G100), .A2(n976), .ZN(n828) );
  NAND2_X1 U921 ( .A1(G136), .A2(n977), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n982), .A2(G124), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT44), .B(n829), .Z(n830) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT111), .ZN(G162) );
  INV_X1 U928 ( .A(n835), .ZN(n837) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(n864) );
  NAND2_X1 U930 ( .A1(G103), .A2(n976), .ZN(n839) );
  NAND2_X1 U931 ( .A1(G139), .A2(n977), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U933 ( .A(KEYINPUT113), .B(n840), .Z(n845) );
  NAND2_X1 U934 ( .A1(G115), .A2(n981), .ZN(n842) );
  NAND2_X1 U935 ( .A1(G127), .A2(n982), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U937 ( .A(KEYINPUT47), .B(n843), .Z(n844) );
  NOR2_X1 U938 ( .A1(n845), .A2(n844), .ZN(n988) );
  XOR2_X1 U939 ( .A(G2072), .B(n988), .Z(n847) );
  XOR2_X1 U940 ( .A(G164), .B(G2078), .Z(n846) );
  NOR2_X1 U941 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT50), .B(n848), .ZN(n862) );
  XNOR2_X1 U943 ( .A(G160), .B(G2084), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n849), .A2(n991), .ZN(n850) );
  NOR2_X1 U945 ( .A1(n851), .A2(n850), .ZN(n853) );
  NAND2_X1 U946 ( .A1(n853), .A2(n852), .ZN(n860) );
  XOR2_X1 U947 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n858) );
  XNOR2_X1 U948 ( .A(G2090), .B(G162), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n854), .B(KEYINPUT117), .ZN(n855) );
  NOR2_X1 U950 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U951 ( .A(n858), .B(n857), .Z(n859) );
  NOR2_X1 U952 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U953 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U954 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U955 ( .A(KEYINPUT52), .B(n865), .Z(n866) );
  NOR2_X1 U956 ( .A1(KEYINPUT55), .A2(n866), .ZN(n867) );
  XNOR2_X1 U957 ( .A(KEYINPUT119), .B(n867), .ZN(n868) );
  NAND2_X1 U958 ( .A1(n868), .A2(G29), .ZN(n919) );
  XOR2_X1 U959 ( .A(G16), .B(KEYINPUT122), .Z(n869) );
  XNOR2_X1 U960 ( .A(KEYINPUT56), .B(n869), .ZN(n894) );
  XNOR2_X1 U961 ( .A(G1966), .B(G168), .ZN(n871) );
  NAND2_X1 U962 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U963 ( .A(n872), .B(KEYINPUT57), .ZN(n891) );
  XNOR2_X1 U964 ( .A(n970), .B(G1341), .ZN(n889) );
  NOR2_X1 U965 ( .A1(n874), .A2(n873), .ZN(n876) );
  NAND2_X1 U966 ( .A1(n876), .A2(n875), .ZN(n880) );
  XOR2_X1 U967 ( .A(G303), .B(G1971), .Z(n878) );
  XOR2_X1 U968 ( .A(G299), .B(G1956), .Z(n877) );
  NAND2_X1 U969 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U970 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U971 ( .A(KEYINPUT124), .B(n881), .ZN(n883) );
  XNOR2_X1 U972 ( .A(n971), .B(G1348), .ZN(n882) );
  NAND2_X1 U973 ( .A1(n883), .A2(n882), .ZN(n886) );
  XNOR2_X1 U974 ( .A(G1961), .B(G171), .ZN(n884) );
  XNOR2_X1 U975 ( .A(KEYINPUT123), .B(n884), .ZN(n885) );
  NOR2_X1 U976 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U977 ( .A(KEYINPUT125), .B(n887), .ZN(n888) );
  NOR2_X1 U978 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U979 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U980 ( .A(KEYINPUT126), .B(n892), .Z(n893) );
  NOR2_X1 U981 ( .A1(n894), .A2(n893), .ZN(n917) );
  XOR2_X1 U982 ( .A(KEYINPUT120), .B(G29), .Z(n913) );
  XNOR2_X1 U983 ( .A(G2072), .B(G33), .ZN(n896) );
  XNOR2_X1 U984 ( .A(G2067), .B(G26), .ZN(n895) );
  NOR2_X1 U985 ( .A1(n896), .A2(n895), .ZN(n904) );
  XOR2_X1 U986 ( .A(G1991), .B(G25), .Z(n897) );
  NAND2_X1 U987 ( .A1(n897), .A2(G28), .ZN(n902) );
  XOR2_X1 U988 ( .A(G1996), .B(G32), .Z(n900) );
  XNOR2_X1 U989 ( .A(n898), .B(G27), .ZN(n899) );
  NAND2_X1 U990 ( .A1(n900), .A2(n899), .ZN(n901) );
  NOR2_X1 U991 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U992 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U993 ( .A(n905), .B(KEYINPUT53), .ZN(n908) );
  XOR2_X1 U994 ( .A(G2084), .B(KEYINPUT54), .Z(n906) );
  XNOR2_X1 U995 ( .A(G34), .B(n906), .ZN(n907) );
  NAND2_X1 U996 ( .A1(n908), .A2(n907), .ZN(n910) );
  XNOR2_X1 U997 ( .A(G35), .B(G2090), .ZN(n909) );
  NOR2_X1 U998 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U999 ( .A(KEYINPUT55), .B(n911), .ZN(n912) );
  NAND2_X1 U1000 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1001 ( .A1(G11), .A2(n914), .ZN(n915) );
  XOR2_X1 U1002 ( .A(KEYINPUT121), .B(n915), .Z(n916) );
  NOR2_X1 U1003 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1004 ( .A1(n919), .A2(n918), .ZN(n943) );
  XNOR2_X1 U1005 ( .A(G5), .B(n920), .ZN(n932) );
  XOR2_X1 U1006 ( .A(G20), .B(G1956), .Z(n924) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G19), .ZN(n922) );
  XNOR2_X1 U1008 ( .A(G1981), .B(G6), .ZN(n921) );
  NOR2_X1 U1009 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1010 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1011 ( .A(KEYINPUT59), .B(G1348), .Z(n925) );
  XNOR2_X1 U1012 ( .A(G4), .B(n925), .ZN(n926) );
  NOR2_X1 U1013 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1014 ( .A(KEYINPUT60), .B(n928), .Z(n930) );
  XNOR2_X1 U1015 ( .A(G1966), .B(G21), .ZN(n929) );
  NOR2_X1 U1016 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1017 ( .A1(n932), .A2(n931), .ZN(n939) );
  XNOR2_X1 U1018 ( .A(G1971), .B(G22), .ZN(n934) );
  XNOR2_X1 U1019 ( .A(G23), .B(G1976), .ZN(n933) );
  NOR2_X1 U1020 ( .A1(n934), .A2(n933), .ZN(n936) );
  XOR2_X1 U1021 ( .A(G1986), .B(G24), .Z(n935) );
  NAND2_X1 U1022 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1023 ( .A(KEYINPUT58), .B(n937), .ZN(n938) );
  NOR2_X1 U1024 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1025 ( .A(KEYINPUT61), .B(n940), .Z(n941) );
  NOR2_X1 U1026 ( .A1(G16), .A2(n941), .ZN(n942) );
  NOR2_X1 U1027 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1028 ( .A(n944), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1029 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1030 ( .A(G132), .ZN(G219) );
  INV_X1 U1031 ( .A(G120), .ZN(G236) );
  INV_X1 U1032 ( .A(G108), .ZN(G238) );
  INV_X1 U1033 ( .A(G96), .ZN(G221) );
  INV_X1 U1034 ( .A(G82), .ZN(G220) );
  INV_X1 U1035 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(G325) );
  INV_X1 U1037 ( .A(G325), .ZN(G261) );
  INV_X1 U1038 ( .A(n947), .ZN(G319) );
  XOR2_X1 U1039 ( .A(n948), .B(G1986), .Z(n959) );
  XOR2_X1 U1040 ( .A(KEYINPUT110), .B(G1981), .Z(n950) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G1971), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n950), .B(n949), .ZN(n955) );
  XOR2_X1 U1043 ( .A(KEYINPUT41), .B(G1991), .Z(n953) );
  XOR2_X1 U1044 ( .A(G1961), .B(n951), .Z(n952) );
  XNOR2_X1 U1045 ( .A(n953), .B(n952), .ZN(n954) );
  XOR2_X1 U1046 ( .A(n955), .B(n954), .Z(n957) );
  XNOR2_X1 U1047 ( .A(G1976), .B(G2474), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n957), .B(n956), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n959), .B(n958), .ZN(G229) );
  XOR2_X1 U1050 ( .A(G2678), .B(G2084), .Z(n961) );
  XNOR2_X1 U1051 ( .A(G2078), .B(G2067), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n961), .B(n960), .ZN(n962) );
  XOR2_X1 U1053 ( .A(n962), .B(KEYINPUT109), .Z(n964) );
  XNOR2_X1 U1054 ( .A(G2072), .B(KEYINPUT42), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n964), .B(n963), .ZN(n968) );
  XOR2_X1 U1056 ( .A(G2100), .B(G2096), .Z(n966) );
  XNOR2_X1 U1057 ( .A(G2090), .B(KEYINPUT43), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n966), .B(n965), .ZN(n967) );
  XOR2_X1 U1059 ( .A(n968), .B(n967), .Z(G227) );
  XNOR2_X1 U1060 ( .A(n970), .B(n969), .ZN(n973) );
  XOR2_X1 U1061 ( .A(G301), .B(n971), .Z(n972) );
  XNOR2_X1 U1062 ( .A(n973), .B(n972), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(n974), .B(G286), .ZN(n975) );
  NOR2_X1 U1064 ( .A1(G37), .A2(n975), .ZN(G397) );
  NAND2_X1 U1065 ( .A1(G106), .A2(n976), .ZN(n979) );
  NAND2_X1 U1066 ( .A1(G142), .A2(n977), .ZN(n978) );
  NAND2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(n980), .B(KEYINPUT45), .ZN(n987) );
  NAND2_X1 U1069 ( .A1(G118), .A2(n981), .ZN(n984) );
  NAND2_X1 U1070 ( .A1(G130), .A2(n982), .ZN(n983) );
  NAND2_X1 U1071 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1072 ( .A(KEYINPUT112), .B(n985), .Z(n986) );
  NAND2_X1 U1073 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(n989), .B(n988), .ZN(n1000) );
  XNOR2_X1 U1075 ( .A(G162), .B(n990), .ZN(n992) );
  XNOR2_X1 U1076 ( .A(n992), .B(n991), .ZN(n996) );
  XOR2_X1 U1077 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n994) );
  XNOR2_X1 U1078 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(n994), .B(n993), .ZN(n995) );
  XOR2_X1 U1080 ( .A(n996), .B(n995), .Z(n998) );
  XNOR2_X1 U1081 ( .A(G164), .B(G160), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(n998), .B(n997), .ZN(n999) );
  XOR2_X1 U1083 ( .A(n1000), .B(n999), .Z(n1001) );
  XNOR2_X1 U1084 ( .A(n1002), .B(n1001), .ZN(n1004) );
  XNOR2_X1 U1085 ( .A(n1004), .B(n1003), .ZN(n1005) );
  NOR2_X1 U1086 ( .A1(G37), .A2(n1005), .ZN(n1006) );
  XNOR2_X1 U1087 ( .A(KEYINPUT116), .B(n1006), .ZN(G395) );
  XOR2_X1 U1088 ( .A(KEYINPUT108), .B(G2446), .Z(n1008) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G2454), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(n1008), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1091 ( .A(n1009), .B(G2451), .Z(n1011) );
  XNOR2_X1 U1092 ( .A(G2430), .B(G2438), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(n1011), .B(n1010), .ZN(n1015) );
  XOR2_X1 U1094 ( .A(G2443), .B(G2435), .Z(n1013) );
  XNOR2_X1 U1095 ( .A(G1348), .B(G2427), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1013), .B(n1012), .ZN(n1014) );
  XOR2_X1 U1097 ( .A(n1015), .B(n1014), .Z(n1016) );
  NAND2_X1 U1098 ( .A1(G14), .A2(n1016), .ZN(n1022) );
  NAND2_X1 U1099 ( .A1(G319), .A2(n1022), .ZN(n1019) );
  NOR2_X1 U1100 ( .A1(G229), .A2(G227), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(KEYINPUT49), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  NOR2_X1 U1103 ( .A1(G397), .A2(G395), .ZN(n1020) );
  NAND2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(G225) );
  INV_X1 U1105 ( .A(G225), .ZN(G308) );
  INV_X1 U1106 ( .A(n1022), .ZN(G401) );
endmodule

