

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X2 U323 ( .A(n361), .B(n360), .ZN(n375) );
  XOR2_X2 U324 ( .A(G29GAT), .B(G43GAT), .Z(n361) );
  XNOR2_X2 U325 ( .A(n353), .B(n352), .ZN(n393) );
  NOR2_X1 U326 ( .A1(n561), .A2(n567), .ZN(n563) );
  NOR2_X1 U327 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U328 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n439) );
  XNOR2_X1 U329 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U330 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n417) );
  XNOR2_X1 U331 ( .A(n303), .B(n302), .ZN(n306) );
  AND2_X1 U332 ( .A1(n488), .A2(n581), .ZN(n489) );
  NOR2_X1 U333 ( .A1(n514), .A2(n506), .ZN(n511) );
  XOR2_X1 U334 ( .A(n423), .B(n422), .Z(n291) );
  XOR2_X1 U335 ( .A(KEYINPUT13), .B(G57GAT), .Z(n343) );
  XNOR2_X1 U336 ( .A(n430), .B(n429), .ZN(n431) );
  INV_X1 U337 ( .A(n374), .ZN(n348) );
  INV_X1 U338 ( .A(KEYINPUT15), .ZN(n300) );
  XNOR2_X1 U339 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U340 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U341 ( .A(n301), .B(n300), .ZN(n302) );
  NOR2_X1 U342 ( .A1(n475), .A2(n474), .ZN(n487) );
  XNOR2_X1 U343 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U344 ( .A(n401), .B(KEYINPUT48), .ZN(n545) );
  XNOR2_X1 U345 ( .A(n342), .B(n341), .ZN(n413) );
  NOR2_X1 U346 ( .A1(n516), .A2(n419), .ZN(n572) );
  XNOR2_X1 U347 ( .A(n440), .B(n439), .ZN(n456) );
  XNOR2_X1 U348 ( .A(n489), .B(KEYINPUT37), .ZN(n515) );
  XOR2_X1 U349 ( .A(n438), .B(n437), .Z(n472) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n581) );
  XOR2_X1 U351 ( .A(n455), .B(n454), .Z(n533) );
  XNOR2_X1 U352 ( .A(KEYINPUT38), .B(n491), .ZN(n500) );
  XNOR2_X1 U353 ( .A(n457), .B(KEYINPUT122), .ZN(n458) );
  XNOR2_X1 U354 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  XOR2_X1 U355 ( .A(G78GAT), .B(G155GAT), .Z(n293) );
  XNOR2_X1 U356 ( .A(G22GAT), .B(G211GAT), .ZN(n292) );
  XNOR2_X1 U357 ( .A(n293), .B(n292), .ZN(n308) );
  XOR2_X1 U358 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n295) );
  XNOR2_X1 U359 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n294) );
  XNOR2_X1 U360 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U361 ( .A(n343), .B(G71GAT), .Z(n297) );
  XOR2_X1 U362 ( .A(G15GAT), .B(G1GAT), .Z(n364) );
  XNOR2_X1 U363 ( .A(n364), .B(G127GAT), .ZN(n296) );
  XNOR2_X1 U364 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U365 ( .A(n299), .B(n298), .Z(n303) );
  NAND2_X1 U366 ( .A1(G231GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U367 ( .A(G8GAT), .B(G183GAT), .ZN(n304) );
  XNOR2_X1 U368 ( .A(n304), .B(KEYINPUT76), .ZN(n406) );
  XNOR2_X1 U369 ( .A(n406), .B(KEYINPUT77), .ZN(n305) );
  XNOR2_X1 U370 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U371 ( .A(G127GAT), .B(KEYINPUT79), .Z(n310) );
  XNOR2_X1 U372 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n309) );
  XNOR2_X1 U373 ( .A(n310), .B(n309), .ZN(n447) );
  XOR2_X1 U374 ( .A(G155GAT), .B(KEYINPUT3), .Z(n312) );
  XNOR2_X1 U375 ( .A(KEYINPUT83), .B(KEYINPUT2), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n423) );
  XNOR2_X1 U377 ( .A(n447), .B(n423), .ZN(n331) );
  XOR2_X1 U378 ( .A(G57GAT), .B(G148GAT), .Z(n314) );
  XNOR2_X1 U379 ( .A(G1GAT), .B(G141GAT), .ZN(n313) );
  XNOR2_X1 U380 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U381 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n316) );
  XNOR2_X1 U382 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n315) );
  XNOR2_X1 U383 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U384 ( .A(n318), .B(n317), .Z(n329) );
  XOR2_X1 U385 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n320) );
  XNOR2_X1 U386 ( .A(KEYINPUT86), .B(KEYINPUT6), .ZN(n319) );
  XNOR2_X1 U387 ( .A(n320), .B(n319), .ZN(n327) );
  XOR2_X1 U388 ( .A(G134GAT), .B(KEYINPUT75), .Z(n378) );
  XOR2_X1 U389 ( .A(G85GAT), .B(G162GAT), .Z(n322) );
  XNOR2_X1 U390 ( .A(G29GAT), .B(G120GAT), .ZN(n321) );
  XNOR2_X1 U391 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U392 ( .A(n378), .B(n323), .Z(n325) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U394 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U395 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U396 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n516) );
  INV_X1 U398 ( .A(n581), .ZN(n554) );
  XOR2_X1 U399 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n333) );
  NAND2_X1 U400 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U401 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U402 ( .A(KEYINPUT32), .B(n334), .ZN(n353) );
  INV_X1 U403 ( .A(G204GAT), .ZN(n342) );
  XOR2_X1 U404 ( .A(G92GAT), .B(KEYINPUT70), .Z(n335) );
  XNOR2_X1 U405 ( .A(G176GAT), .B(G64GAT), .ZN(n336) );
  NAND2_X1 U406 ( .A1(n335), .A2(n336), .ZN(n340) );
  INV_X1 U407 ( .A(n335), .ZN(n338) );
  INV_X1 U408 ( .A(n336), .ZN(n337) );
  NAND2_X1 U409 ( .A1(n338), .A2(n337), .ZN(n339) );
  NAND2_X1 U410 ( .A1(n340), .A2(n339), .ZN(n341) );
  XNOR2_X1 U411 ( .A(n413), .B(n343), .ZN(n345) );
  XOR2_X1 U412 ( .A(KEYINPUT67), .B(KEYINPUT31), .Z(n344) );
  XNOR2_X1 U413 ( .A(n345), .B(n344), .ZN(n351) );
  XOR2_X1 U414 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  XOR2_X1 U415 ( .A(G148GAT), .B(G78GAT), .Z(n427) );
  XNOR2_X1 U416 ( .A(n450), .B(n427), .ZN(n349) );
  XOR2_X1 U417 ( .A(G85GAT), .B(KEYINPUT68), .Z(n347) );
  XNOR2_X1 U418 ( .A(G99GAT), .B(G106GAT), .ZN(n346) );
  XNOR2_X1 U419 ( .A(n347), .B(n346), .ZN(n374) );
  XNOR2_X1 U420 ( .A(n393), .B(KEYINPUT41), .ZN(n505) );
  XOR2_X1 U421 ( .A(G8GAT), .B(G197GAT), .Z(n355) );
  XNOR2_X1 U422 ( .A(G169GAT), .B(G113GAT), .ZN(n354) );
  XNOR2_X1 U423 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U424 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n357) );
  XNOR2_X1 U425 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n369) );
  XNOR2_X1 U428 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n360) );
  XOR2_X1 U429 ( .A(G141GAT), .B(G22GAT), .Z(n429) );
  XOR2_X1 U430 ( .A(n375), .B(n429), .Z(n363) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U433 ( .A(n365), .B(n364), .Z(n367) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(G50GAT), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U436 ( .A(n369), .B(n368), .Z(n547) );
  NAND2_X1 U437 ( .A1(n505), .A2(n547), .ZN(n371) );
  XOR2_X1 U438 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n370) );
  XOR2_X1 U439 ( .A(n371), .B(n370), .Z(n372) );
  NOR2_X1 U440 ( .A1(n554), .A2(n372), .ZN(n373) );
  XNOR2_X1 U441 ( .A(KEYINPUT112), .B(n373), .ZN(n391) );
  XOR2_X1 U442 ( .A(n375), .B(n374), .Z(n390) );
  XOR2_X1 U443 ( .A(KEYINPUT71), .B(KEYINPUT73), .Z(n377) );
  XNOR2_X1 U444 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n377), .B(n376), .ZN(n382) );
  XOR2_X1 U446 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n380) );
  XOR2_X1 U447 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XNOR2_X1 U448 ( .A(n422), .B(n378), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U450 ( .A(n382), .B(n381), .Z(n384) );
  NAND2_X1 U451 ( .A1(G232GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U453 ( .A(n385), .B(KEYINPUT74), .Z(n388) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(G190GAT), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n386), .B(G218GAT), .ZN(n409) );
  XNOR2_X1 U456 ( .A(n409), .B(KEYINPUT72), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n556) );
  INV_X1 U459 ( .A(n556), .ZN(n568) );
  NAND2_X1 U460 ( .A1(n391), .A2(n568), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n392), .B(KEYINPUT47), .ZN(n400) );
  XOR2_X1 U462 ( .A(KEYINPUT36), .B(n556), .Z(n584) );
  NOR2_X1 U463 ( .A1(n581), .A2(n584), .ZN(n396) );
  XOR2_X1 U464 ( .A(KEYINPUT113), .B(KEYINPUT45), .Z(n394) );
  XNOR2_X1 U465 ( .A(KEYINPUT64), .B(n394), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n393), .A2(n397), .ZN(n398) );
  NOR2_X1 U468 ( .A1(n547), .A2(n398), .ZN(n399) );
  XOR2_X1 U469 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n403) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U472 ( .A(n404), .B(KEYINPUT90), .Z(n408) );
  XNOR2_X1 U473 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n405), .B(G211GAT), .ZN(n434) );
  XNOR2_X1 U475 ( .A(n434), .B(n406), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U477 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U478 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n412) );
  XNOR2_X1 U479 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n445) );
  XNOR2_X1 U481 ( .A(n445), .B(n413), .ZN(n414) );
  XOR2_X1 U482 ( .A(n415), .B(n414), .Z(n520) );
  XOR2_X1 U483 ( .A(n520), .B(KEYINPUT118), .Z(n416) );
  NOR2_X1 U484 ( .A1(n545), .A2(n416), .ZN(n418) );
  XOR2_X1 U485 ( .A(KEYINPUT82), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U486 ( .A(KEYINPUT81), .B(KEYINPUT22), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n438) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n291), .B(n424), .ZN(n432) );
  XOR2_X1 U490 ( .A(G204GAT), .B(KEYINPUT23), .Z(n426) );
  XNOR2_X1 U491 ( .A(G218GAT), .B(G106GAT), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U493 ( .A(n428), .B(n427), .Z(n430) );
  XOR2_X1 U494 ( .A(n433), .B(KEYINPUT85), .Z(n436) );
  XNOR2_X1 U495 ( .A(n434), .B(KEYINPUT84), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U497 ( .A1(n572), .A2(n472), .ZN(n440) );
  XOR2_X1 U498 ( .A(G183GAT), .B(KEYINPUT80), .Z(n442) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(G99GAT), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n455) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT20), .Z(n444) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U504 ( .A(n446), .B(n445), .Z(n449) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U507 ( .A(n451), .B(n450), .Z(n453) );
  XNOR2_X1 U508 ( .A(G190GAT), .B(G134GAT), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U510 ( .A1(n456), .A2(n533), .ZN(n567) );
  NOR2_X1 U511 ( .A1(n581), .A2(n567), .ZN(n459) );
  INV_X1 U512 ( .A(G183GAT), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n393), .A2(n547), .ZN(n490) );
  NOR2_X1 U514 ( .A1(n556), .A2(n581), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT16), .ZN(n477) );
  NAND2_X1 U516 ( .A1(n520), .A2(n533), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n461), .A2(n472), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT96), .ZN(n463) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(n463), .ZN(n468) );
  XNOR2_X1 U520 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n533), .A2(n472), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n465), .B(n464), .ZN(n571) );
  XNOR2_X1 U523 ( .A(n520), .B(KEYINPUT27), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n571), .A2(n470), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(KEYINPUT95), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n516), .A2(n469), .ZN(n475) );
  NAND2_X1 U528 ( .A1(n470), .A2(n516), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT93), .ZN(n543) );
  XOR2_X1 U530 ( .A(n472), .B(KEYINPUT28), .Z(n526) );
  INV_X1 U531 ( .A(n526), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n543), .A2(n473), .ZN(n531) );
  NOR2_X1 U533 ( .A1(n533), .A2(n531), .ZN(n474) );
  INV_X1 U534 ( .A(n487), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n506) );
  NOR2_X1 U536 ( .A1(n490), .A2(n506), .ZN(n485) );
  NAND2_X1 U537 ( .A1(n485), .A2(n516), .ZN(n480) );
  XOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT34), .Z(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT97), .B(n478), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n520), .A2(n485), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U544 ( .A1(n485), .A2(n533), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n485), .A2(n526), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NOR2_X1 U550 ( .A1(n487), .A2(n584), .ZN(n488) );
  NOR2_X1 U551 ( .A1(n515), .A2(n490), .ZN(n491) );
  NAND2_X1 U552 ( .A1(n516), .A2(n500), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n495) );
  NAND2_X1 U555 ( .A1(n500), .A2(n520), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n498) );
  NAND2_X1 U559 ( .A1(n533), .A2(n500), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G43GAT), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n500), .A2(n526), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT102), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(KEYINPUT103), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(n504), .Z(n508) );
  INV_X1 U568 ( .A(n547), .ZN(n573) );
  INV_X1 U569 ( .A(n505), .ZN(n561) );
  NAND2_X1 U570 ( .A1(n573), .A2(n505), .ZN(n514) );
  NAND2_X1 U571 ( .A1(n511), .A2(n516), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n520), .A2(n511), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n511), .A2(n533), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U578 ( .A1(n511), .A2(n526), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n518) );
  NOR2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n527), .A2(n516), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT107), .Z(n522) );
  NAND2_X1 U586 ( .A1(n527), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1337GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n524) );
  NAND2_X1 U589 ( .A1(n527), .A2(n533), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n529) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  NOR2_X1 U596 ( .A1(n545), .A2(n531), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n573), .A2(n540), .ZN(n534) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  NOR2_X1 U600 ( .A1(n561), .A2(n540), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n581), .A2(n540), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U607 ( .A1(n568), .A2(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n571), .A2(n543), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT115), .B(n546), .Z(n557) );
  NAND2_X1 U613 ( .A1(n547), .A2(n557), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT116), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n551) );
  NAND2_X1 U617 ( .A1(n557), .A2(n505), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .Z(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n557), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n558), .ZN(G1347GAT) );
  NOR2_X1 U625 ( .A1(n573), .A2(n567), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n564), .ZN(G1349GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(G1351GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n583) );
  NOR2_X1 U637 ( .A1(n573), .A2(n583), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT125), .B(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n393), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

