//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  AOI21_X1  g006(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  AOI211_X1 g011(.A(new_n195), .B(G146), .C1(new_n191), .C2(new_n192), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT24), .B(G110), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n207), .B(new_n203), .C1(new_n208), .C2(KEYINPUT23), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n206), .B1(G110), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n197), .A2(new_n199), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(new_n205), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n209), .B2(G110), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT73), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n212), .B(new_n215), .C1(new_n209), .C2(G110), .ZN(new_n216));
  XNOR2_X1  g030(.A(G125), .B(G140), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n196), .A3(new_n216), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT74), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G137), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n211), .A2(new_n220), .A3(new_n226), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G217), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(G234), .B2(new_n232), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n230), .A2(G902), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n228), .A2(new_n232), .A3(new_n229), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n228), .A2(KEYINPUT75), .A3(new_n232), .A4(new_n229), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n238), .A2(KEYINPUT76), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n233), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n236), .B2(new_n239), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT25), .B1(new_n236), .B2(new_n237), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n235), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G472), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  INV_X1    g063(.A(G237), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n222), .A3(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n249), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT2), .B(G113), .Z(new_n256));
  XNOR2_X1  g070(.A(G116), .B(G119), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n202), .A2(G116), .ZN(new_n259));
  INV_X1    g073(.A(G116), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G119), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(KEYINPUT67), .A3(new_n264), .ZN(new_n265));
  OR3_X1    g079(.A1(new_n256), .A2(KEYINPUT67), .A3(new_n257), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(G137), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n270), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n269), .A2(G137), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n271), .A2(G134), .ZN(new_n277));
  OAI21_X1  g091(.A(G131), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G143), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n283), .A3(G146), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n280), .A2(G146), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n289));
  OAI21_X1  g103(.A(G128), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G146), .B1(new_n281), .B2(new_n283), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n218), .A2(G143), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n279), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  NOR2_X1   g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n282), .A2(G143), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n218), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n292), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT64), .B(G143), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n285), .B1(new_n305), .B2(G146), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT65), .B1(new_n306), .B2(new_n296), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n284), .A2(KEYINPUT65), .A3(new_n286), .A4(new_n296), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n304), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G131), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n275), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(KEYINPUT66), .A3(G131), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n295), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT30), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n284), .A2(new_n286), .A3(new_n296), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n308), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n322), .A2(new_n315), .A3(new_n314), .A4(new_n304), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n295), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n267), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n267), .B(new_n295), .C1(new_n310), .C2(new_n316), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n255), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(KEYINPUT70), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n267), .B1(new_n323), .B2(new_n295), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n334));
  INV_X1    g148(.A(new_n267), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n317), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n327), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n327), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n344), .A3(new_n254), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n329), .B(new_n330), .C1(new_n339), .C2(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n342), .A2(new_n344), .A3(new_n254), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n317), .A2(new_n335), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n340), .B1(new_n348), .B2(new_n327), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(new_n330), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n248), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G472), .A2(G902), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT32), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n314), .A2(new_n315), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n303), .B1(new_n321), .B2(new_n308), .ZN(new_n359));
  AOI211_X1 g173(.A(KEYINPUT30), .B(new_n294), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n324), .B1(new_n323), .B2(new_n295), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n335), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n327), .A3(new_n254), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT31), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n362), .A2(KEYINPUT31), .A3(new_n327), .A4(new_n254), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n344), .B(new_n342), .C1(new_n333), .C2(new_n338), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n255), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n357), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n352), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n365), .A2(new_n366), .B1(new_n368), .B2(new_n255), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n355), .B1(new_n372), .B2(new_n354), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n247), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G469), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n288), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n284), .A2(KEYINPUT78), .A3(new_n286), .A4(new_n287), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n200), .B1(new_n301), .B2(KEYINPUT1), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n306), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G104), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G107), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n390));
  OAI22_X1  g204(.A1(new_n390), .A2(KEYINPUT3), .B1(new_n385), .B2(G104), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n386), .B1(KEYINPUT77), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n390), .A2(new_n385), .A3(KEYINPUT3), .A4(G104), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n389), .B1(new_n395), .B2(new_n384), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(KEYINPUT77), .A2(new_n392), .B1(new_n387), .B2(G107), .ZN(new_n398));
  AND4_X1   g212(.A1(new_n390), .A2(new_n385), .A3(KEYINPUT3), .A4(G104), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n390), .A2(KEYINPUT3), .B1(new_n385), .B2(G104), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n384), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n389), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n288), .A3(new_n293), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT12), .B1(new_n405), .B2(new_n358), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT12), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n407), .B(new_n316), .C1(new_n397), .C2(new_n404), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT80), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G128), .B1(new_n291), .B2(new_n289), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n284), .A2(new_n286), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n410), .A2(new_n411), .B1(new_n288), .B2(new_n379), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n403), .B1(new_n412), .B2(new_n381), .ZN(new_n413));
  INV_X1    g227(.A(new_n404), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n358), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n405), .A2(KEYINPUT12), .A3(new_n358), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G140), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n222), .A2(G227), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n293), .A2(new_n288), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n396), .A2(new_n423), .A3(KEYINPUT10), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G101), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n395), .A2(new_n384), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n424), .B1(new_n430), .B2(new_n310), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT10), .B1(new_n383), .B2(new_n396), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n422), .B1(new_n433), .B2(new_n316), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n409), .A2(new_n419), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n422), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n397), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(G101), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n359), .A2(new_n441), .A3(new_n427), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n438), .A2(new_n439), .A3(new_n442), .A4(new_n424), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT79), .B1(new_n431), .B2(new_n432), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n358), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n438), .A2(new_n316), .A3(new_n442), .A4(new_n424), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n436), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n378), .B(new_n232), .C1(new_n435), .C2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n406), .B2(new_n408), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n449), .A2(new_n422), .B1(new_n445), .B2(new_n434), .ZN(new_n450));
  OAI21_X1  g264(.A(G469), .B1(new_n450), .B2(G902), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n377), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n262), .A2(new_n263), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT5), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(G113), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n455), .B1(new_n458), .B2(KEYINPUT81), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n460), .A3(new_n457), .A4(G113), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n396), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G122), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n428), .A2(new_n429), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n427), .A2(new_n266), .A3(new_n265), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n462), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT6), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n463), .B(KEYINPUT82), .Z(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n310), .A2(KEYINPUT83), .A3(G125), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n359), .B2(new_n189), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n423), .B2(G125), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n293), .A2(KEYINPUT84), .A3(new_n189), .A4(new_n288), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G224), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(G953), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n473), .A2(new_n475), .A3(new_n479), .A4(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n471), .A2(new_n472), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n459), .A2(new_n403), .A3(new_n461), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n458), .A2(new_n258), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n396), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n463), .B(KEYINPUT8), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n477), .A2(new_n478), .B1(new_n310), .B2(G125), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT85), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n484), .B1(new_n493), .B2(KEYINPUT7), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n493), .B2(KEYINPUT7), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n466), .B(new_n491), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n484), .A2(KEYINPUT7), .ZN(new_n497));
  AND4_X1   g311(.A1(new_n475), .A2(new_n473), .A3(new_n479), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n232), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n454), .B1(new_n486), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n466), .A2(new_n491), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n310), .A2(G125), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n495), .B1(new_n479), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n189), .B1(new_n322), .B2(new_n304), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n505), .A2(KEYINPUT83), .B1(new_n477), .B2(new_n478), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n475), .A3(new_n497), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n484), .B1(new_n506), .B2(new_n475), .ZN(new_n509));
  INV_X1    g323(.A(new_n485), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n466), .A2(KEYINPUT6), .B1(new_n468), .B2(new_n469), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n513), .A3(new_n453), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n500), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G214), .B1(G237), .B2(G902), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G475), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n250), .A2(new_n222), .A3(G214), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n305), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n250), .A2(new_n222), .A3(G143), .A4(G214), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n273), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n281), .A2(new_n283), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n250), .A2(new_n222), .A3(G214), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G131), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n520), .A2(new_n273), .A3(new_n521), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n196), .A2(new_n195), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n193), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n523), .B(new_n530), .C1(new_n532), .C2(new_n198), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n188), .A2(new_n190), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G146), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n219), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n273), .ZN(new_n538));
  OAI221_X1 g352(.A(new_n536), .B1(new_n526), .B2(new_n538), .C1(new_n527), .C2(new_n537), .ZN(new_n539));
  XOR2_X1   g353(.A(G113), .B(G122), .Z(new_n540));
  XOR2_X1   g354(.A(KEYINPUT90), .B(G104), .Z(new_n541));
  XOR2_X1   g355(.A(new_n540), .B(new_n541), .Z(new_n542));
  AND3_X1   g356(.A1(new_n533), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n533), .B2(new_n539), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n232), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n518), .B1(new_n545), .B2(KEYINPUT91), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n232), .C1(new_n543), .C2(new_n544), .ZN(new_n548));
  NOR2_X1   g362(.A1(G475), .A2(G902), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT19), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT88), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n534), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n217), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n553));
  AOI21_X1  g367(.A(G146), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n196), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT89), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n526), .A2(G131), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT87), .B1(new_n557), .B2(new_n522), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT19), .B1(new_n217), .B2(KEYINPUT88), .ZN(new_n559));
  AND4_X1   g373(.A1(KEYINPUT88), .A2(new_n188), .A3(new_n190), .A4(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n218), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n196), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT87), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n527), .A2(new_n564), .A3(new_n529), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n556), .A2(new_n558), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n542), .B1(new_n566), .B2(new_n539), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n549), .B1(new_n567), .B2(new_n543), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT20), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n572), .B(new_n549), .C1(new_n567), .C2(new_n543), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n546), .A2(new_n548), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(G234), .A2(G237), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n575), .A2(G952), .A3(new_n222), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n575), .A2(G902), .A3(G953), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT21), .B(G898), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n581));
  INV_X1    g395(.A(G122), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(G116), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n260), .A2(KEYINPUT92), .A3(G122), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(G116), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n385), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(KEYINPUT93), .A3(new_n385), .A4(new_n586), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n281), .A2(new_n283), .A3(G128), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n200), .A2(G143), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n269), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n269), .B1(new_n591), .B2(new_n592), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n589), .B(new_n590), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n585), .A2(KEYINPUT14), .B1(G116), .B2(new_n582), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT14), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n583), .A2(new_n598), .A3(new_n584), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n385), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n591), .A2(new_n592), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT13), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G134), .B1(new_n591), .B2(KEYINPUT13), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n585), .A2(new_n385), .A3(new_n586), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n385), .B1(new_n585), .B2(new_n586), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n593), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n596), .A2(new_n600), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n375), .A2(new_n231), .A3(G953), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI221_X1 g426(.A(new_n610), .B1(new_n605), .B2(new_n608), .C1(new_n596), .C2(new_n600), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G478), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(KEYINPUT15), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(G902), .B(new_n616), .C1(new_n612), .C2(new_n613), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n574), .A2(new_n580), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n517), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n374), .A2(new_n452), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  NAND2_X1  g438(.A1(new_n448), .A2(new_n451), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n241), .A2(new_n233), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n245), .A2(new_n240), .ZN(new_n627));
  INV_X1    g441(.A(new_n244), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n234), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n625), .A2(new_n630), .A3(new_n376), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n367), .A2(new_n369), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n232), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n633), .A2(G472), .B1(new_n353), .B2(new_n632), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT94), .Z(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n515), .A2(new_n516), .A3(new_n580), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(G475), .A3(new_n548), .ZN(new_n640));
  INV_X1    g454(.A(new_n549), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n566), .A2(new_n539), .ZN(new_n642));
  INV_X1    g456(.A(new_n542), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n533), .A2(new_n539), .A3(new_n542), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n573), .B1(new_n646), .B2(new_n569), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n612), .A2(new_n613), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT33), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n612), .A2(new_n613), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(G478), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n615), .A2(new_n232), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n614), .B2(new_n615), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n637), .B1(new_n638), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n516), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n660), .B(new_n579), .C1(new_n500), .C2(new_n514), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n574), .A2(new_n656), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(KEYINPUT95), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n636), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT96), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  XNOR2_X1  g483(.A(new_n614), .B(new_n617), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n644), .A2(new_n645), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n569), .B1(new_n671), .B2(new_n549), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n549), .B(new_n569), .C1(new_n567), .C2(new_n543), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n640), .B(new_n670), .C1(new_n672), .C2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n638), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n636), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NOR2_X1   g493(.A1(new_n227), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n221), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n233), .A2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n242), .B2(new_n246), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n634), .A2(new_n452), .A3(new_n622), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT37), .B(G110), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT97), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT98), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n685), .B(new_n688), .ZN(G12));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n640), .A2(new_n670), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n577), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n576), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n672), .B2(new_n674), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n690), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n695), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n571), .B2(new_n673), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n699), .A2(KEYINPUT99), .A3(new_n640), .A4(new_n670), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n697), .A2(new_n684), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n346), .A2(new_n351), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G472), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n632), .A2(new_n356), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n373), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n660), .B1(new_n500), .B2(new_n514), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n701), .A2(new_n705), .A3(new_n452), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  NOR2_X1   g522(.A1(new_n326), .A2(new_n328), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n255), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n348), .A2(new_n327), .A3(new_n255), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n232), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n373), .A2(new_n704), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n373), .A2(new_n704), .A3(KEYINPUT100), .A4(new_n713), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n684), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n515), .B(KEYINPUT38), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n620), .B1(new_n640), .B2(new_n647), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n516), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n695), .B(KEYINPUT39), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n452), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n723), .B1(new_n725), .B2(KEYINPUT40), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n720), .B(new_n726), .C1(KEYINPUT40), .C2(new_n725), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n524), .ZN(G45));
  INV_X1    g542(.A(new_n684), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n648), .A2(new_n657), .A3(new_n695), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n705), .A3(new_n452), .A4(new_n706), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  INV_X1    g547(.A(new_n448), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n409), .A2(new_n419), .A3(new_n434), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n442), .B(new_n424), .C1(new_n413), .C2(KEYINPUT10), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n316), .B1(new_n736), .B2(KEYINPUT79), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n737), .A2(new_n443), .B1(new_n316), .B2(new_n433), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n735), .B1(new_n738), .B2(new_n436), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n378), .B1(new_n739), .B2(new_n232), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n705), .A2(new_n741), .A3(new_n630), .A4(new_n376), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n664), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT41), .B(G113), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  NOR3_X1   g559(.A1(new_n734), .A2(new_n740), .A3(new_n377), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n705), .A3(new_n630), .A4(new_n676), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  OAI21_X1  g562(.A(new_n436), .B1(new_n736), .B2(new_n358), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n416), .A2(new_n417), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n749), .B1(new_n750), .B2(KEYINPUT80), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n445), .A2(new_n446), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n419), .A2(new_n751), .B1(new_n752), .B2(new_n422), .ZN(new_n753));
  OAI21_X1  g567(.A(G469), .B1(new_n753), .B2(G902), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n376), .A2(new_n754), .A3(new_n448), .A4(new_n706), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n729), .A2(new_n621), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n705), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G119), .ZN(G21));
  NAND2_X1  g572(.A1(new_n342), .A2(new_n344), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n255), .B1(new_n759), .B2(new_n349), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n354), .B1(new_n367), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT101), .B(G472), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n761), .B1(new_n633), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n722), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n638), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n746), .A2(new_n630), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  INV_X1    g581(.A(new_n761), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n574), .A2(new_n656), .A3(new_n698), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n762), .B1(new_n372), .B2(G902), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n684), .A2(new_n768), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n755), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  INV_X1    g587(.A(KEYINPUT102), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n705), .A2(new_n630), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n500), .A2(new_n514), .A3(new_n516), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n730), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n452), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n774), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n776), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n376), .A2(new_n625), .A3(new_n769), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n374), .A3(KEYINPUT102), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT42), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n373), .A2(new_n704), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT103), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT103), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n373), .A2(new_n704), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n703), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT42), .A3(new_n630), .A4(new_n781), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G131), .ZN(G33));
  AND2_X1   g606(.A1(new_n697), .A2(new_n700), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n776), .A2(new_n377), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n374), .A2(new_n625), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT106), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n574), .A2(new_n657), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT105), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n648), .A2(new_n656), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT105), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT43), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n802), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT104), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n799), .B2(new_n800), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n798), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n805), .B(KEYINPUT106), .C1(new_n807), .C2(new_n809), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n634), .A2(new_n729), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n797), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n449), .A2(new_n422), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n445), .A2(new_n434), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n378), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  NAND2_X1  g636(.A1(G469), .A2(G902), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT46), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n734), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(KEYINPUT46), .A3(new_n823), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n377), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n776), .B(KEYINPUT107), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n827), .A2(new_n724), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n813), .A4(new_n814), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n816), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  NAND4_X1  g646(.A1(new_n777), .A2(new_n371), .A3(new_n373), .A4(new_n247), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n827), .A2(KEYINPUT47), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n827), .A2(KEYINPUT47), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  NOR2_X1   g653(.A1(G952), .A2(G953), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT117), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n806), .A2(new_n810), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n763), .A2(new_n630), .A3(new_n576), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n721), .A2(new_n516), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n746), .A3(new_n845), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT50), .Z(new_n847));
  NAND3_X1  g661(.A1(new_n741), .A2(new_n576), .A3(new_n794), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n684), .A3(new_n763), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n848), .A2(new_n247), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n719), .A2(new_n574), .A3(new_n656), .A4(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n837), .ZN(new_n855));
  INV_X1    g669(.A(new_n741), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT114), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT114), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n377), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n835), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n828), .A3(new_n844), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT51), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n847), .A2(KEYINPUT51), .A3(new_n853), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n860), .A2(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n844), .A2(new_n828), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n860), .B2(KEYINPUT115), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n849), .A2(new_n630), .A3(new_n789), .ZN(new_n868));
  XOR2_X1   g682(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n719), .A2(new_n662), .A3(new_n851), .ZN(new_n871));
  INV_X1    g685(.A(G952), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n872), .B(G953), .C1(new_n844), .C2(new_n755), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  OR3_X1    g688(.A1(new_n862), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n763), .A2(new_n452), .A3(new_n684), .A4(new_n777), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n699), .A2(new_n640), .A3(new_n620), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n776), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n705), .A2(new_n452), .A3(new_n684), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n794), .A2(new_n625), .A3(new_n697), .A4(new_n700), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n877), .B(new_n880), .C1(new_n775), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT112), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n795), .A2(new_n884), .A3(new_n877), .A4(new_n880), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n883), .A2(new_n885), .B1(new_n784), .B2(new_n790), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT110), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT109), .B1(new_n574), .B2(new_n656), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT109), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n648), .A2(new_n657), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n891), .B2(new_n638), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n661), .A2(KEYINPUT110), .A3(new_n888), .A4(new_n890), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n634), .A3(new_n631), .A4(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n894), .A2(KEYINPUT111), .A3(new_n623), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT111), .B1(new_n894), .B2(new_n623), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n640), .A2(new_n670), .A3(new_n647), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n638), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n634), .A2(new_n899), .A3(new_n630), .A4(new_n452), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n747), .B(new_n900), .C1(new_n664), .C2(new_n742), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n757), .A2(new_n766), .A3(new_n685), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n886), .A2(new_n897), .A3(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n722), .A2(new_n515), .A3(new_n516), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n452), .A3(new_n695), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n714), .A2(new_n715), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n684), .B(new_n906), .C1(new_n907), .C2(new_n717), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n772), .A2(new_n707), .A3(new_n732), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT52), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n697), .A2(new_n684), .A3(new_n700), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n373), .B2(new_n371), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n452), .A2(new_n706), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n912), .A2(new_n913), .B1(new_n755), .B2(new_n771), .ZN(new_n914));
  INV_X1    g728(.A(new_n906), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n729), .B(new_n915), .C1(new_n716), .C2(new_n718), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT52), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n914), .A2(new_n916), .A3(new_n917), .A4(new_n732), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n876), .B1(new_n904), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n772), .A2(new_n707), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT52), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n910), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n894), .A2(new_n623), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT111), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n894), .A2(new_n623), .A3(KEYINPUT111), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n903), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n923), .A2(KEYINPUT53), .A3(new_n928), .A4(new_n886), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n920), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n904), .A2(new_n876), .A3(new_n919), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT113), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n883), .A2(new_n885), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n791), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n903), .A2(new_n926), .A3(new_n927), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT53), .B1(new_n939), .B2(new_n923), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n931), .B1(new_n941), .B2(new_n930), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n841), .B1(new_n875), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n630), .A2(new_n376), .A3(new_n516), .A4(new_n802), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n856), .B2(KEYINPUT49), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT108), .Z(new_n946));
  INV_X1    g760(.A(KEYINPUT49), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n721), .B1(new_n947), .B2(new_n741), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n719), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n943), .A2(new_n949), .ZN(G75));
  NOR2_X1   g764(.A1(new_n222), .A2(G952), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n920), .A2(new_n929), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n232), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n955), .B2(G210), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n511), .A2(new_n512), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n483), .A3(new_n485), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n513), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT55), .Z(new_n960));
  OAI21_X1  g774(.A(new_n952), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n956), .B2(new_n960), .ZN(G51));
  INV_X1    g776(.A(KEYINPUT119), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n954), .A2(new_n232), .A3(new_n822), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n823), .B(KEYINPUT57), .Z(new_n965));
  AOI21_X1  g779(.A(new_n930), .B1(new_n920), .B2(new_n929), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT118), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n931), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g782(.A(KEYINPUT118), .B(new_n930), .C1(new_n920), .C2(new_n929), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n964), .B1(new_n970), .B2(new_n739), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n963), .B1(new_n971), .B2(new_n951), .ZN(new_n972));
  INV_X1    g786(.A(new_n919), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT53), .B1(new_n939), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n910), .A2(new_n918), .A3(new_n922), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n904), .A2(new_n876), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT54), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT118), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n966), .A2(new_n967), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n931), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n753), .B1(new_n980), .B2(new_n965), .ZN(new_n981));
  OAI211_X1 g795(.A(KEYINPUT119), .B(new_n952), .C1(new_n981), .C2(new_n964), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n972), .A2(new_n982), .ZN(G54));
  NAND2_X1  g797(.A1(KEYINPUT58), .A2(G475), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT120), .Z(new_n985));
  AND3_X1   g799(.A1(new_n955), .A2(new_n671), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n671), .B1(new_n955), .B2(new_n985), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n986), .A2(new_n987), .A3(new_n951), .ZN(G60));
  NAND2_X1  g802(.A1(new_n650), .A2(new_n652), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n654), .B(KEYINPUT59), .Z(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n942), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n980), .A2(new_n989), .A3(new_n990), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n951), .ZN(G63));
  OAI21_X1  g807(.A(new_n952), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n994));
  XNOR2_X1  g808(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n231), .A2(new_n232), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n995), .B(new_n996), .Z(new_n997));
  NOR2_X1   g811(.A1(new_n954), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n994), .B1(new_n998), .B2(new_n681), .ZN(new_n999));
  INV_X1    g813(.A(new_n230), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n998), .ZN(new_n1001));
  NAND2_X1  g815(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n578), .B2(new_n481), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n928), .B2(G953), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n957), .B1(G898), .B2(new_n222), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT123), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1005), .B(new_n1007), .ZN(G69));
  NAND2_X1  g822(.A1(new_n318), .A2(new_n325), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n559), .A2(new_n560), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT124), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1009), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n838), .A2(new_n831), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n789), .A2(new_n630), .A3(new_n905), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1017), .A2(new_n724), .A3(new_n827), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT125), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1017), .A2(KEYINPUT125), .A3(new_n724), .A4(new_n827), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n795), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n1023), .B(new_n909), .C1(new_n784), .C2(new_n790), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1015), .A2(new_n1016), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1022), .A2(new_n831), .A3(new_n838), .A4(new_n1024), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(KEYINPUT126), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n222), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n222), .A2(G900), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1014), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(G953), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1033), .A2(KEYINPUT127), .A3(new_n1030), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1013), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n222), .B1(G227), .B2(G900), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n727), .A2(new_n732), .A3(new_n914), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT62), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n776), .B1(new_n891), .B2(new_n898), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n374), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1040), .B1(new_n725), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1015), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1012), .B1(new_n1045), .B2(G953), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1035), .A2(new_n1037), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1029), .A2(new_n1014), .A3(new_n1031), .ZN(new_n1048));
  OAI21_X1  g862(.A(KEYINPUT127), .B1(new_n1033), .B2(new_n1030), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1012), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g864(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1013), .B1(new_n1051), .B2(new_n222), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1036), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1047), .A2(new_n1053), .ZN(G72));
  NAND2_X1  g868(.A1(new_n329), .A2(new_n363), .ZN(new_n1055));
  NAND2_X1  g869(.A1(G472), .A2(G902), .ZN(new_n1056));
  XOR2_X1   g870(.A(new_n1056), .B(KEYINPUT63), .Z(new_n1057));
  NAND2_X1  g871(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1057), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1059), .B1(new_n1045), .B2(new_n928), .ZN(new_n1060));
  INV_X1    g874(.A(new_n710), .ZN(new_n1061));
  OAI221_X1 g875(.A(new_n952), .B1(new_n941), .B2(new_n1058), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g876(.A(new_n1057), .B1(new_n1028), .B2(new_n938), .ZN(new_n1063));
  AND3_X1   g877(.A1(new_n1063), .A2(new_n255), .A3(new_n709), .ZN(new_n1064));
  NOR2_X1   g878(.A1(new_n1062), .A2(new_n1064), .ZN(G57));
endmodule


