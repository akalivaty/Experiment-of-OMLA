

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(G1966), .A2(n830), .ZN(n761) );
  NOR2_X1 U556 ( .A1(n761), .A2(n758), .ZN(n734) );
  XNOR2_X1 U557 ( .A(n700), .B(KEYINPUT64), .ZN(n705) );
  NAND2_X1 U558 ( .A1(n733), .A2(G8), .ZN(n830) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  XOR2_X1 U560 ( .A(KEYINPUT29), .B(n731), .Z(n521) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n537), .Z(n904) );
  BUF_X1 U562 ( .A(n733), .Z(n742) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n796) );
  NOR2_X1 U564 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U565 ( .A1(n774), .A2(n771), .ZN(n772) );
  INV_X1 U566 ( .A(KEYINPUT33), .ZN(n771) );
  INV_X1 U567 ( .A(KEYINPUT102), .ZN(n780) );
  INV_X1 U568 ( .A(n992), .ZN(n766) );
  OR2_X1 U569 ( .A1(n830), .A2(n829), .ZN(n522) );
  AND2_X1 U570 ( .A1(n831), .A2(n522), .ZN(n523) );
  NOR2_X1 U571 ( .A1(n764), .A2(n763), .ZN(n782) );
  AND2_X1 U572 ( .A1(n767), .A2(n766), .ZN(n768) );
  INV_X1 U573 ( .A(n701), .ZN(n733) );
  INV_X1 U574 ( .A(KEYINPUT70), .ZN(n591) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n539), .ZN(n907) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n664) );
  XNOR2_X1 U577 ( .A(n592), .B(n591), .ZN(n593) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n909) );
  XNOR2_X1 U579 ( .A(n605), .B(KEYINPUT15), .ZN(n999) );
  NOR2_X1 U580 ( .A1(n595), .A2(n594), .ZN(n984) );
  INV_X1 U581 ( .A(G543), .ZN(n524) );
  XOR2_X1 U582 ( .A(KEYINPUT66), .B(G651), .Z(n532) );
  NOR2_X1 U583 ( .A1(G543), .A2(n532), .ZN(n525) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n525), .Z(n660) );
  NAND2_X1 U585 ( .A1(G60), .A2(n660), .ZN(n531) );
  INV_X1 U586 ( .A(KEYINPUT0), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n526), .A2(G543), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n524), .A2(KEYINPUT0), .ZN(n527) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n645) );
  NOR2_X1 U590 ( .A1(n645), .A2(G651), .ZN(n529) );
  XOR2_X1 U591 ( .A(KEYINPUT65), .B(n529), .Z(n596) );
  BUF_X1 U592 ( .A(n596), .Z(n661) );
  NAND2_X1 U593 ( .A1(G47), .A2(n661), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G85), .A2(n664), .ZN(n534) );
  NOR2_X1 U596 ( .A1(n645), .A2(n532), .ZN(n665) );
  NAND2_X1 U597 ( .A1(G72), .A2(n665), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  OR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(G290) );
  NAND2_X1 U600 ( .A1(n904), .A2(G137), .ZN(n698) );
  INV_X1 U601 ( .A(G2105), .ZN(n539) );
  AND2_X1 U602 ( .A1(n539), .A2(G2104), .ZN(n626) );
  NAND2_X1 U603 ( .A1(G101), .A2(n626), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT23), .B(n538), .ZN(n543) );
  NAND2_X1 U605 ( .A1(G125), .A2(n907), .ZN(n541) );
  NAND2_X1 U606 ( .A1(G113), .A2(n909), .ZN(n540) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n696) );
  AND2_X1 U609 ( .A1(n698), .A2(n696), .ZN(G160) );
  XNOR2_X1 U610 ( .A(KEYINPUT104), .B(G2451), .ZN(n553) );
  XOR2_X1 U611 ( .A(G2446), .B(G2430), .Z(n545) );
  XNOR2_X1 U612 ( .A(G2454), .B(G2435), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n549) );
  XOR2_X1 U614 ( .A(G2438), .B(G2427), .Z(n547) );
  XNOR2_X1 U615 ( .A(G1348), .B(G1341), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U617 ( .A(n549), .B(n548), .Z(n551) );
  XNOR2_X1 U618 ( .A(G2443), .B(KEYINPUT105), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  AND2_X1 U621 ( .A1(n554), .A2(G14), .ZN(G401) );
  AND2_X1 U622 ( .A1(G452), .A2(G94), .ZN(G173) );
  AND2_X1 U623 ( .A1(n904), .A2(G138), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G114), .A2(n909), .ZN(n555) );
  XOR2_X1 U625 ( .A(KEYINPUT87), .B(n555), .Z(n557) );
  NAND2_X1 U626 ( .A1(G102), .A2(n626), .ZN(n556) );
  AND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U628 ( .A1(G126), .A2(n907), .ZN(n558) );
  NAND2_X1 U629 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U630 ( .A1(n561), .A2(n560), .ZN(G164) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  INV_X1 U632 ( .A(G82), .ZN(G220) );
  NAND2_X1 U633 ( .A1(G64), .A2(n660), .ZN(n563) );
  NAND2_X1 U634 ( .A1(G52), .A2(n661), .ZN(n562) );
  NAND2_X1 U635 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n665), .A2(G77), .ZN(n564) );
  XOR2_X1 U637 ( .A(KEYINPUT67), .B(n564), .Z(n566) );
  NAND2_X1 U638 ( .A1(n664), .A2(G90), .ZN(n565) );
  NAND2_X1 U639 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U640 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U641 ( .A1(n569), .A2(n568), .ZN(G171) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G63), .A2(n660), .ZN(n571) );
  NAND2_X1 U644 ( .A1(G51), .A2(n661), .ZN(n570) );
  NAND2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U646 ( .A(n572), .B(KEYINPUT6), .ZN(n573) );
  XNOR2_X1 U647 ( .A(n573), .B(KEYINPUT75), .ZN(n580) );
  XNOR2_X1 U648 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n664), .A2(G89), .ZN(n574) );
  XNOR2_X1 U650 ( .A(n574), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U651 ( .A1(G76), .A2(n665), .ZN(n575) );
  NAND2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U653 ( .A(n578), .B(n577), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U655 ( .A(KEYINPUT7), .B(n581), .ZN(G168) );
  XOR2_X1 U656 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n582), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U659 ( .A(G223), .ZN(n845) );
  NAND2_X1 U660 ( .A1(n845), .A2(G567), .ZN(n583) );
  XNOR2_X1 U661 ( .A(n583), .B(KEYINPUT11), .ZN(n584) );
  XNOR2_X1 U662 ( .A(KEYINPUT69), .B(n584), .ZN(G234) );
  NAND2_X1 U663 ( .A1(n660), .A2(G56), .ZN(n585) );
  XNOR2_X1 U664 ( .A(n585), .B(KEYINPUT14), .ZN(n587) );
  NAND2_X1 U665 ( .A1(G43), .A2(n661), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n664), .A2(G81), .ZN(n588) );
  XNOR2_X1 U668 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U669 ( .A1(G68), .A2(n665), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U671 ( .A(KEYINPUT13), .B(n593), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n984), .A2(G860), .ZN(G153) );
  NAND2_X1 U673 ( .A1(n596), .A2(G54), .ZN(n597) );
  XOR2_X1 U674 ( .A(KEYINPUT71), .B(n597), .Z(n599) );
  NAND2_X1 U675 ( .A1(n665), .A2(G79), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U677 ( .A(KEYINPUT72), .B(n600), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G66), .A2(n660), .ZN(n602) );
  NAND2_X1 U679 ( .A1(G92), .A2(n664), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U682 ( .A(n999), .ZN(n658) );
  NOR2_X1 U683 ( .A1(n658), .A2(G868), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT73), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G868), .A2(G301), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G284) );
  AND2_X1 U687 ( .A1(n660), .A2(G65), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G53), .A2(n661), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G91), .A2(n664), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n665), .A2(G78), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(G299) );
  INV_X1 U694 ( .A(G868), .ZN(n678) );
  XNOR2_X1 U695 ( .A(KEYINPUT76), .B(n678), .ZN(n615) );
  NOR2_X1 U696 ( .A1(G286), .A2(n615), .ZN(n617) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(G297) );
  INV_X1 U699 ( .A(G860), .ZN(n852) );
  NAND2_X1 U700 ( .A1(n852), .A2(G559), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n618), .A2(n658), .ZN(n619) );
  XNOR2_X1 U702 ( .A(n619), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U703 ( .A1(n658), .A2(G868), .ZN(n620) );
  NOR2_X1 U704 ( .A1(G559), .A2(n620), .ZN(n622) );
  AND2_X1 U705 ( .A1(n678), .A2(n984), .ZN(n621) );
  NOR2_X1 U706 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U707 ( .A1(n907), .A2(G123), .ZN(n623) );
  XNOR2_X1 U708 ( .A(n623), .B(KEYINPUT18), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G111), .A2(n909), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G99), .A2(n626), .ZN(n628) );
  NAND2_X1 U712 ( .A1(G135), .A2(n904), .ZN(n627) );
  NAND2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n933) );
  XNOR2_X1 U715 ( .A(n933), .B(G2096), .ZN(n632) );
  INV_X1 U716 ( .A(G2100), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U718 ( .A1(G61), .A2(n660), .ZN(n634) );
  NAND2_X1 U719 ( .A1(G86), .A2(n664), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U721 ( .A(n635), .B(KEYINPUT79), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n637) );
  NAND2_X1 U723 ( .A1(G73), .A2(n665), .ZN(n636) );
  XNOR2_X1 U724 ( .A(n637), .B(n636), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G48), .A2(n661), .ZN(n638) );
  XNOR2_X1 U726 ( .A(KEYINPUT81), .B(n638), .ZN(n639) );
  NOR2_X1 U727 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U729 ( .A(n643), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G74), .A2(G651), .ZN(n644) );
  XNOR2_X1 U731 ( .A(n644), .B(KEYINPUT78), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G49), .A2(n661), .ZN(n647) );
  NAND2_X1 U733 ( .A1(G87), .A2(n645), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U735 ( .A1(n660), .A2(n648), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U737 ( .A1(G88), .A2(n664), .ZN(n652) );
  NAND2_X1 U738 ( .A1(G75), .A2(n665), .ZN(n651) );
  NAND2_X1 U739 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U740 ( .A(KEYINPUT83), .B(n653), .ZN(n657) );
  NAND2_X1 U741 ( .A1(G62), .A2(n660), .ZN(n655) );
  NAND2_X1 U742 ( .A1(G50), .A2(n661), .ZN(n654) );
  AND2_X1 U743 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U744 ( .A1(n657), .A2(n656), .ZN(G303) );
  INV_X1 U745 ( .A(G303), .ZN(G166) );
  NAND2_X1 U746 ( .A1(G559), .A2(n658), .ZN(n659) );
  XNOR2_X1 U747 ( .A(n659), .B(n984), .ZN(n851) );
  NAND2_X1 U748 ( .A1(G67), .A2(n660), .ZN(n663) );
  NAND2_X1 U749 ( .A1(G55), .A2(n661), .ZN(n662) );
  NAND2_X1 U750 ( .A1(n663), .A2(n662), .ZN(n669) );
  NAND2_X1 U751 ( .A1(G93), .A2(n664), .ZN(n667) );
  NAND2_X1 U752 ( .A1(G80), .A2(n665), .ZN(n666) );
  NAND2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U755 ( .A(KEYINPUT77), .B(n670), .ZN(n853) );
  XOR2_X1 U756 ( .A(G305), .B(n853), .Z(n676) );
  XOR2_X1 U757 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n671) );
  XNOR2_X1 U758 ( .A(G288), .B(n671), .ZN(n672) );
  XNOR2_X1 U759 ( .A(G290), .B(n672), .ZN(n674) );
  INV_X1 U760 ( .A(G299), .ZN(n989) );
  XNOR2_X1 U761 ( .A(n989), .B(G166), .ZN(n673) );
  XNOR2_X1 U762 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U763 ( .A(n676), .B(n675), .ZN(n920) );
  XNOR2_X1 U764 ( .A(n851), .B(n920), .ZN(n677) );
  NAND2_X1 U765 ( .A1(n677), .A2(G868), .ZN(n680) );
  NAND2_X1 U766 ( .A1(n678), .A2(n853), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U768 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U769 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U770 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U771 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XOR2_X1 U773 ( .A(KEYINPUT85), .B(G44), .Z(n685) );
  XNOR2_X1 U774 ( .A(KEYINPUT3), .B(n685), .ZN(G218) );
  XOR2_X1 U775 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NOR2_X1 U776 ( .A1(G219), .A2(G220), .ZN(n686) );
  XOR2_X1 U777 ( .A(KEYINPUT86), .B(n686), .Z(n687) );
  XNOR2_X1 U778 ( .A(n687), .B(KEYINPUT22), .ZN(n688) );
  NOR2_X1 U779 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U780 ( .A1(G96), .A2(n689), .ZN(n849) );
  NAND2_X1 U781 ( .A1(G2106), .A2(n849), .ZN(n693) );
  NAND2_X1 U782 ( .A1(G69), .A2(G120), .ZN(n690) );
  NOR2_X1 U783 ( .A1(G237), .A2(n690), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G108), .A2(n691), .ZN(n850) );
  NAND2_X1 U785 ( .A1(G567), .A2(n850), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n876) );
  NAND2_X1 U787 ( .A1(G661), .A2(G483), .ZN(n694) );
  NOR2_X1 U788 ( .A1(n876), .A2(n694), .ZN(n848) );
  NAND2_X1 U789 ( .A1(n848), .A2(G36), .ZN(G176) );
  XOR2_X1 U790 ( .A(G2078), .B(KEYINPUT25), .Z(n965) );
  AND2_X1 U791 ( .A1(n696), .A2(G40), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n797) );
  INV_X1 U793 ( .A(n797), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n796), .A2(n699), .ZN(n700) );
  INV_X1 U795 ( .A(n705), .ZN(n701) );
  INV_X1 U796 ( .A(n733), .ZN(n721) );
  NAND2_X1 U797 ( .A1(n965), .A2(n721), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n742), .A2(G1961), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n737) );
  NOR2_X1 U800 ( .A1(G301), .A2(n737), .ZN(n704) );
  XNOR2_X1 U801 ( .A(n704), .B(KEYINPUT93), .ZN(n732) );
  NAND2_X1 U802 ( .A1(n705), .A2(G1348), .ZN(n706) );
  XOR2_X1 U803 ( .A(KEYINPUT95), .B(n706), .Z(n708) );
  NAND2_X1 U804 ( .A1(G2067), .A2(n721), .ZN(n707) );
  NAND2_X1 U805 ( .A1(n708), .A2(n707), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n717), .A2(n999), .ZN(n711) );
  NAND2_X1 U807 ( .A1(G1341), .A2(n733), .ZN(n709) );
  XNOR2_X1 U808 ( .A(n709), .B(KEYINPUT94), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n716) );
  INV_X1 U810 ( .A(G1996), .ZN(n712) );
  OR2_X1 U811 ( .A1(n733), .A2(n712), .ZN(n713) );
  XNOR2_X1 U812 ( .A(n713), .B(KEYINPUT26), .ZN(n714) );
  NAND2_X1 U813 ( .A1(n714), .A2(n984), .ZN(n715) );
  NOR2_X1 U814 ( .A1(n716), .A2(n715), .ZN(n719) );
  NOR2_X1 U815 ( .A1(n717), .A2(n999), .ZN(n718) );
  NOR2_X1 U816 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U817 ( .A(n720), .B(KEYINPUT96), .ZN(n726) );
  NAND2_X1 U818 ( .A1(G2072), .A2(n721), .ZN(n722) );
  XNOR2_X1 U819 ( .A(n722), .B(KEYINPUT27), .ZN(n724) );
  INV_X1 U820 ( .A(G1956), .ZN(n1014) );
  NOR2_X1 U821 ( .A1(n721), .A2(n1014), .ZN(n723) );
  NOR2_X1 U822 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n727), .A2(n989), .ZN(n725) );
  NAND2_X1 U824 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U825 ( .A1(n727), .A2(n989), .ZN(n728) );
  XOR2_X1 U826 ( .A(n728), .B(KEYINPUT28), .Z(n729) );
  NAND2_X1 U827 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U828 ( .A1(n732), .A2(n521), .ZN(n757) );
  NOR2_X1 U829 ( .A1(n742), .A2(G2084), .ZN(n758) );
  NAND2_X1 U830 ( .A1(G8), .A2(n734), .ZN(n735) );
  XNOR2_X1 U831 ( .A(KEYINPUT30), .B(n735), .ZN(n736) );
  NOR2_X1 U832 ( .A1(n736), .A2(G168), .ZN(n740) );
  NAND2_X1 U833 ( .A1(G301), .A2(n737), .ZN(n738) );
  XNOR2_X1 U834 ( .A(n738), .B(KEYINPUT97), .ZN(n739) );
  XOR2_X1 U835 ( .A(KEYINPUT31), .B(n741), .Z(n756) );
  INV_X1 U836 ( .A(G8), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n742), .A2(G2090), .ZN(n744) );
  NOR2_X1 U838 ( .A1(G1971), .A2(n830), .ZN(n743) );
  NOR2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U840 ( .A(n745), .B(KEYINPUT98), .ZN(n746) );
  NAND2_X1 U841 ( .A1(n746), .A2(G303), .ZN(n747) );
  OR2_X1 U842 ( .A1(n748), .A2(n747), .ZN(n750) );
  AND2_X1 U843 ( .A1(n756), .A2(n750), .ZN(n749) );
  NAND2_X1 U844 ( .A1(n757), .A2(n749), .ZN(n753) );
  INV_X1 U845 ( .A(n750), .ZN(n751) );
  OR2_X1 U846 ( .A1(n751), .A2(G286), .ZN(n752) );
  NAND2_X1 U847 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U848 ( .A(KEYINPUT32), .B(KEYINPUT99), .ZN(n754) );
  XNOR2_X1 U849 ( .A(n755), .B(n754), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n757), .A2(n756), .ZN(n760) );
  NAND2_X1 U851 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n762) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  INV_X1 U854 ( .A(n782), .ZN(n769) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n765) );
  XOR2_X1 U856 ( .A(n765), .B(KEYINPUT100), .Z(n767) );
  NOR2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n992) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NAND2_X1 U860 ( .A1(n770), .A2(n993), .ZN(n773) );
  INV_X1 U861 ( .A(n830), .ZN(n774) );
  OR2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n992), .A2(n774), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n775), .A2(KEYINPUT33), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT101), .B(n778), .ZN(n779) );
  XNOR2_X1 U867 ( .A(G305), .B(G1981), .ZN(n982) );
  NOR2_X1 U868 ( .A1(n779), .A2(n982), .ZN(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(n780), .ZN(n832) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G8), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n769), .A2(n784), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n830), .A2(n785), .ZN(n827) );
  NAND2_X1 U874 ( .A1(n626), .A2(G104), .ZN(n786) );
  XOR2_X1 U875 ( .A(KEYINPUT89), .B(n786), .Z(n788) );
  NAND2_X1 U876 ( .A1(n904), .A2(G140), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n789), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G128), .A2(n907), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G116), .A2(n909), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U882 ( .A(KEYINPUT35), .B(n792), .Z(n793) );
  NOR2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U884 ( .A(KEYINPUT36), .B(n795), .Z(n916) );
  XOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .Z(n824) );
  AND2_X1 U886 ( .A1(n916), .A2(n824), .ZN(n949) );
  NOR2_X1 U887 ( .A1(n796), .A2(n797), .ZN(n836) );
  NAND2_X1 U888 ( .A1(n949), .A2(n836), .ZN(n838) );
  INV_X1 U889 ( .A(n838), .ZN(n823) );
  NAND2_X1 U890 ( .A1(G105), .A2(n626), .ZN(n798) );
  XNOR2_X1 U891 ( .A(n798), .B(KEYINPUT92), .ZN(n799) );
  XNOR2_X1 U892 ( .A(KEYINPUT38), .B(n799), .ZN(n802) );
  NAND2_X1 U893 ( .A1(G129), .A2(n907), .ZN(n800) );
  XOR2_X1 U894 ( .A(KEYINPUT91), .B(n800), .Z(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G117), .A2(n909), .ZN(n804) );
  NAND2_X1 U897 ( .A1(G141), .A2(n904), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n885) );
  AND2_X1 U900 ( .A1(n712), .A2(n885), .ZN(n936) );
  NAND2_X1 U901 ( .A1(G119), .A2(n907), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G131), .A2(n904), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U904 ( .A1(G107), .A2(n909), .ZN(n810) );
  NAND2_X1 U905 ( .A1(G95), .A2(n626), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n901) );
  NAND2_X1 U908 ( .A1(G1991), .A2(n901), .ZN(n813) );
  XOR2_X1 U909 ( .A(KEYINPUT90), .B(n813), .Z(n815) );
  NOR2_X1 U910 ( .A1(n885), .A2(n712), .ZN(n814) );
  NOR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n835) );
  INV_X1 U912 ( .A(n835), .ZN(n943) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n901), .ZN(n934) );
  NOR2_X1 U915 ( .A1(n816), .A2(n934), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n943), .A2(n817), .ZN(n818) );
  XOR2_X1 U917 ( .A(KEYINPUT103), .B(n818), .Z(n819) );
  NOR2_X1 U918 ( .A1(n936), .A2(n819), .ZN(n820) );
  XNOR2_X1 U919 ( .A(KEYINPUT39), .B(n820), .ZN(n821) );
  NAND2_X1 U920 ( .A1(n821), .A2(n836), .ZN(n822) );
  OR2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n916), .A2(n824), .ZN(n953) );
  NAND2_X1 U923 ( .A1(n953), .A2(n836), .ZN(n825) );
  AND2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n833) );
  AND2_X1 U925 ( .A1(n827), .A2(n833), .ZN(n831) );
  NOR2_X1 U926 ( .A1(G305), .A2(G1981), .ZN(n828) );
  XOR2_X1 U927 ( .A(n828), .B(KEYINPUT24), .Z(n829) );
  NAND2_X1 U928 ( .A1(n832), .A2(n523), .ZN(n843) );
  INV_X1 U929 ( .A(n833), .ZN(n841) );
  XOR2_X1 U930 ( .A(KEYINPUT88), .B(G1986), .Z(n834) );
  XNOR2_X1 U931 ( .A(G290), .B(n834), .ZN(n985) );
  NAND2_X1 U932 ( .A1(n835), .A2(n985), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(n839) );
  AND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  OR2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  AND2_X1 U936 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U937 ( .A(n844), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U940 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U942 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U944 ( .A(G120), .ZN(G236) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n854), .B(n853), .ZN(G145) );
  XOR2_X1 U950 ( .A(G2474), .B(G1981), .Z(n856) );
  XNOR2_X1 U951 ( .A(G1966), .B(G1961), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U953 ( .A(n857), .B(KEYINPUT109), .Z(n859) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U956 ( .A(G1986), .B(G1976), .Z(n861) );
  XNOR2_X1 U957 ( .A(G1956), .B(G1971), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U959 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U960 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(G229) );
  XOR2_X1 U962 ( .A(G2100), .B(KEYINPUT108), .Z(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT107), .B(G2678), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U965 ( .A(KEYINPUT42), .B(G2090), .Z(n869) );
  XNOR2_X1 U966 ( .A(G2067), .B(G2072), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U968 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U969 ( .A(KEYINPUT43), .B(G2096), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U971 ( .A(G2078), .B(G2084), .Z(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(G227) );
  XOR2_X1 U973 ( .A(KEYINPUT106), .B(n876), .Z(G319) );
  NAND2_X1 U974 ( .A1(G124), .A2(n907), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n877), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G100), .A2(n626), .ZN(n878) );
  XOR2_X1 U977 ( .A(KEYINPUT111), .B(n878), .Z(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G112), .A2(n909), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G136), .A2(n904), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(G162) );
  XOR2_X1 U983 ( .A(n933), .B(n885), .Z(n887) );
  XNOR2_X1 U984 ( .A(G164), .B(G160), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n900) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n898) );
  NAND2_X1 U987 ( .A1(G106), .A2(n626), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G142), .A2(n904), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n890), .B(KEYINPUT45), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G130), .A2(n907), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n909), .A2(G118), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT112), .B(n893), .Z(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n896), .B(KEYINPUT113), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n901), .B(G162), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n918) );
  NAND2_X1 U1001 ( .A1(G103), .A2(n626), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(G139), .A2(n904), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n914) );
  NAND2_X1 U1004 ( .A1(n907), .A2(G127), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(KEYINPUT114), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n909), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(KEYINPUT47), .B(n912), .Z(n913) );
  NOR2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1010 ( .A(KEYINPUT115), .B(n915), .Z(n944) );
  XOR2_X1 U1011 ( .A(n944), .B(n916), .Z(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n919), .ZN(G395) );
  XOR2_X1 U1014 ( .A(n920), .B(G286), .Z(n922) );
  XNOR2_X1 U1015 ( .A(n984), .B(G171), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(n922), .B(n921), .ZN(n923) );
  XOR2_X1 U1017 ( .A(n923), .B(n999), .Z(n924) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n924), .ZN(G397) );
  NOR2_X1 U1019 ( .A1(G229), .A2(G227), .ZN(n925) );
  XOR2_X1 U1020 ( .A(KEYINPUT49), .B(n925), .Z(n926) );
  XNOR2_X1 U1021 ( .A(KEYINPUT117), .B(n926), .ZN(n930) );
  INV_X1 U1022 ( .A(G319), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n927), .A2(G401), .ZN(n928) );
  XOR2_X1 U1024 ( .A(KEYINPUT116), .B(n928), .Z(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n932) );
  NOR2_X1 U1026 ( .A1(G395), .A2(G397), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1028 ( .A(G225), .ZN(G308) );
  INV_X1 U1029 ( .A(G96), .ZN(G221) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n941) );
  XOR2_X1 U1032 ( .A(G160), .B(G2084), .Z(n939) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT51), .B(n937), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n951) );
  XOR2_X1 U1039 ( .A(G2072), .B(n944), .Z(n946) );
  XOR2_X1 U1040 ( .A(G164), .B(G2078), .Z(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1042 ( .A(KEYINPUT50), .B(n947), .Z(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n976), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n956), .A2(G29), .ZN(n1040) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G35), .ZN(n971) );
  XNOR2_X1 U1051 ( .A(G2072), .B(G33), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G1991), .B(G25), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(G32), .B(n712), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n959), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT118), .B(G2067), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G26), .B(n960), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n968) );
  XOR2_X1 U1060 ( .A(G27), .B(n965), .Z(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT119), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n969), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1069 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n979), .ZN(n1038) );
  INV_X1 U1072 ( .A(G16), .ZN(n1034) );
  XOR2_X1 U1073 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n980) );
  XNOR2_X1 U1074 ( .A(n1034), .B(n980), .ZN(n1005) );
  XOR2_X1 U1075 ( .A(G168), .B(G1966), .Z(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1077 ( .A(KEYINPUT57), .B(n983), .Z(n1003) );
  XNOR2_X1 U1078 ( .A(n984), .B(G1341), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G301), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n998) );
  XNOR2_X1 U1082 ( .A(G166), .B(G1971), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n989), .B(G1956), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n766), .A2(n993), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT121), .B(n996), .Z(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G1348), .B(n999), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1036) );
  XNOR2_X1 U1093 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n1032) );
  XNOR2_X1 U1094 ( .A(G1986), .B(G24), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G1976), .B(G23), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT125), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1011), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT58), .ZN(n1030) );
  XOR2_X1 U1102 ( .A(G1961), .B(KEYINPUT122), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(G5), .B(n1013), .ZN(n1026) );
  XNOR2_X1 U1104 ( .A(KEYINPUT123), .B(G20), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(n1014), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G19), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(G6), .B(G1981), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1109 ( .A(KEYINPUT124), .B(n1018), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(G1348), .B(G4), .ZN(n1019) );
  XNOR2_X1 U1111 ( .A(n1019), .B(KEYINPUT59), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(n1024), .B(KEYINPUT60), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(G21), .B(G1966), .ZN(n1027) );
  NOR2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(n1032), .B(n1031), .ZN(n1033) );
  NAND2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1123 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

