//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n548, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT67), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n469), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  AOI21_X1  g052(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n466), .B2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  AND2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NOR2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(G138), .B(new_n469), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n468), .A2(new_n490), .A3(G138), .A4(new_n469), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n469), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n496), .A2(new_n500), .B1(new_n480), .B2(G126), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n504), .A2(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n512), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g098(.A(KEYINPUT70), .B(new_n519), .C1(new_n510), .C2(new_n520), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT5), .B(G543), .Z(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n514), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n505), .A2(new_n506), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT69), .B(G51), .Z(new_n530));
  AOI22_X1  g105(.A1(new_n526), .A2(G63), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n523), .A2(new_n524), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(G90), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT71), .B(G52), .Z(new_n535));
  OAI22_X1  g110(.A1(new_n510), .A2(new_n534), .B1(new_n508), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n540), .A2(new_n508), .B1(new_n510), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n514), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g122(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n548));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n525), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n525), .A2(new_n527), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n554), .A2(G651), .B1(new_n555), .B2(G91), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(KEYINPUT74), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n558), .B(G543), .C1(new_n506), .C2(new_n505), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  AOI22_X1  g140(.A1(new_n555), .A2(G87), .B1(new_n529), .B2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(KEYINPUT76), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(G288));
  AOI22_X1  g145(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n514), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n555), .A2(G86), .B1(new_n529), .B2(G48), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(G72), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G60), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n525), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n514), .B1(new_n577), .B2(KEYINPUT77), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n578), .B1(KEYINPUT77), .B2(new_n577), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n555), .A2(G85), .B1(new_n529), .B2(G47), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G290));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n582));
  INV_X1    g157(.A(G92), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n510), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n525), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n529), .B2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(G171), .ZN(G284));
  OAI21_X1  g169(.A(new_n593), .B1(new_n592), .B2(G171), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(new_n556), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n600), .B2(G868), .ZN(G297));
  OAI21_X1  g176(.A(new_n596), .B1(new_n600), .B2(G868), .ZN(G280));
  INV_X1    g177(.A(new_n591), .ZN(new_n603));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G860), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT78), .ZN(G148));
  OAI21_X1  g181(.A(KEYINPUT79), .B1(new_n545), .B2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n604), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  MUX2_X1   g184(.A(KEYINPUT79), .B(new_n607), .S(new_n609), .Z(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n468), .A2(new_n463), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT12), .Z(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  INV_X1    g189(.A(G2100), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n478), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n480), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n469), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT80), .Z(G156));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT81), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(G14), .B1(new_n637), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT83), .Z(G401));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(new_n615), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n623), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n665), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G22), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G166), .B2(new_n676), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G1971), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(G6), .ZN(new_n680));
  INV_X1    g255(.A(G305), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n676), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT32), .B(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n682), .B(new_n684), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n676), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n676), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT33), .ZN(new_n690));
  INV_X1    g265(.A(G1976), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(KEYINPUT34), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n686), .A2(new_n692), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n478), .A2(G131), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n480), .A2(G119), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n469), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT84), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n699), .B1(new_n706), .B2(new_n698), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT85), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G24), .B(G290), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT86), .B(G1986), .Z(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  NAND4_X1  g288(.A1(new_n695), .A2(new_n697), .A3(new_n710), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT36), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT98), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n478), .A2(G141), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT91), .Z(new_n719));
  AND2_X1   g294(.A1(new_n463), .A2(G105), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT26), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n720), .B(new_n722), .C1(G129), .C2(new_n480), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n698), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n727));
  INV_X1    g302(.A(G32), .ZN(new_n728));
  AOI21_X1  g303(.A(KEYINPUT93), .B1(new_n698), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n725), .B2(new_n698), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n717), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G171), .A2(new_n676), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G5), .B2(new_n676), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  NOR2_X1   g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n698), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT90), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G160), .B2(G29), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n734), .A2(G1961), .B1(G2084), .B2(new_n739), .ZN(new_n740));
  OR3_X1    g315(.A1(new_n731), .A2(KEYINPUT96), .A3(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n676), .A2(G20), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n600), .B2(new_n676), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n727), .A2(new_n730), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n717), .ZN(new_n748));
  OAI21_X1  g323(.A(KEYINPUT96), .B1(new_n731), .B2(new_n740), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT25), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n468), .A2(G127), .ZN(new_n752));
  NAND2_X1  g327(.A1(G115), .A2(G2104), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n469), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n751), .B(new_n754), .C1(G139), .C2(new_n478), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n698), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n698), .B2(G33), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n757), .A2(new_n758), .B1(G2084), .B2(new_n739), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n603), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G4), .B2(G16), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n698), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n698), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT29), .B(G2090), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n759), .A2(new_n763), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n545), .B2(G16), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT88), .B(G1341), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n698), .A2(G27), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G164), .B2(new_n698), .ZN(new_n775));
  INV_X1    g350(.A(G2078), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n773), .B(new_n777), .C1(new_n757), .C2(new_n758), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n478), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n480), .A2(G128), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n469), .A2(G116), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT89), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n698), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2067), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n769), .A2(new_n778), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n741), .A2(new_n748), .A3(new_n749), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n676), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n676), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n793), .A2(KEYINPUT94), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(KEYINPUT94), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n794), .A2(new_n795), .A3(G1966), .ZN(new_n796));
  OAI21_X1  g371(.A(G1966), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT30), .B(G28), .ZN(new_n798));
  OR2_X1    g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  NAND2_X1  g374(.A1(KEYINPUT31), .A2(G11), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n798), .A2(new_n698), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n622), .B2(new_n698), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n734), .B2(G1961), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n796), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT95), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n791), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n715), .A2(new_n716), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n716), .B1(new_n715), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(G311));
  NAND2_X1  g384(.A1(new_n715), .A2(new_n806), .ZN(G150));
  AOI22_X1  g385(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(new_n514), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n555), .A2(G93), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n529), .A2(G55), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n814), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n603), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  INV_X1    g397(.A(new_n545), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n545), .B(new_n812), .C1(new_n816), .C2(new_n817), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n822), .A2(new_n826), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(KEYINPUT39), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT100), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT39), .B1(new_n827), .B2(new_n828), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n831), .B1(new_n830), .B2(new_n833), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n820), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT102), .ZN(G145));
  XOR2_X1   g412(.A(new_n783), .B(KEYINPUT104), .Z(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT105), .ZN(new_n840));
  OR3_X1    g415(.A1(new_n840), .A2(new_n469), .A3(G118), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n469), .B2(G118), .ZN(new_n842));
  OR2_X1    g417(.A1(G106), .A2(G2105), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n841), .A2(G2104), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n480), .A2(G130), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n478), .A2(G142), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n704), .B(KEYINPUT106), .ZN(new_n848));
  INV_X1    g423(.A(new_n613), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  INV_X1    g429(.A(new_n847), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n856), .A3(new_n502), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n502), .B1(new_n853), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n839), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n853), .A2(new_n856), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G164), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(new_n838), .A3(new_n857), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n725), .A2(new_n755), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n724), .B2(new_n755), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n860), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n860), .B2(new_n863), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(G160), .B(KEYINPUT103), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G162), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n622), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n866), .B2(new_n867), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g451(.A1(new_n818), .A2(new_n592), .ZN(new_n877));
  XOR2_X1   g452(.A(G303), .B(KEYINPUT108), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G288), .ZN(new_n879));
  XNOR2_X1  g454(.A(G290), .B(G305), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n878), .B(new_n688), .ZN(new_n882));
  INV_X1    g457(.A(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n826), .B(new_n608), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(new_n600), .B2(new_n591), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(G299), .A2(new_n603), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n600), .A2(new_n888), .A3(new_n591), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT41), .B1(new_n895), .B2(new_n889), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n890), .A2(new_n897), .A3(new_n891), .A4(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n894), .B1(new_n899), .B2(new_n887), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n886), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n877), .B1(new_n901), .B2(new_n592), .ZN(G295));
  OAI21_X1  g477(.A(new_n877), .B1(new_n901), .B2(new_n592), .ZN(G331));
  AND2_X1   g478(.A1(new_n881), .A2(new_n884), .ZN(new_n904));
  NOR2_X1   g479(.A1(G301), .A2(KEYINPUT109), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT109), .B1(new_n536), .B2(new_n538), .ZN(new_n906));
  NAND2_X1  g481(.A1(G286), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT110), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n909));
  NAND3_X1  g484(.A1(G286), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n824), .A3(new_n825), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n826), .A2(new_n908), .A3(new_n910), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n905), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n905), .A3(new_n913), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n915), .A2(new_n893), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n899), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n904), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n893), .A3(new_n916), .ZN(new_n921));
  INV_X1    g496(.A(new_n916), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(new_n914), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n885), .B(new_n921), .C1(new_n923), .C2(new_n899), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n919), .A2(new_n924), .A3(new_n927), .A4(new_n920), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(KEYINPUT111), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n931), .A3(KEYINPUT43), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n926), .A2(KEYINPUT44), .A3(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G397));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n489), .A2(new_n491), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n496), .A2(new_n500), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n480), .A2(G126), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n936), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n476), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n945), .A3(G40), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n948), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT46), .B1(new_n948), .B2(G1996), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n783), .B(G2067), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n951), .A2(new_n724), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n949), .A2(new_n950), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT47), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(G1996), .B2(new_n724), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n725), .B2(G1996), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n947), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n706), .A2(new_n708), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n958), .A2(new_n959), .B1(G2067), .B2(new_n783), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT125), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n947), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n704), .B(new_n708), .Z(new_n964));
  OAI21_X1  g539(.A(new_n947), .B1(new_n956), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n948), .A2(G290), .A3(G1986), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT48), .Z(new_n967));
  AOI211_X1 g542(.A(new_n954), .B(new_n963), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT45), .B1(new_n502), .B2(new_n936), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n942), .A2(G1384), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT113), .B1(new_n502), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G40), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n472), .A2(new_n476), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n502), .A2(KEYINPUT113), .A3(new_n970), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT56), .B(G2072), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n972), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n597), .A2(new_n561), .A3(KEYINPUT57), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(G299), .B2(KEYINPUT57), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n941), .A2(KEYINPUT50), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n492), .B2(new_n501), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n974), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1956), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n977), .A2(new_n979), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n974), .A2(new_n981), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(G2067), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n984), .B2(new_n762), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n591), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n979), .B1(new_n977), .B2(new_n986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n591), .B1(new_n990), .B2(KEYINPUT60), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n946), .B1(new_n941), .B2(KEYINPUT50), .ZN(new_n995));
  AOI21_X1  g570(.A(G1348), .B1(new_n995), .B2(new_n983), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT60), .ZN(new_n997));
  NOR4_X1   g572(.A1(new_n996), .A2(new_n997), .A3(new_n603), .A4(new_n989), .ZN(new_n998));
  OAI22_X1  g573(.A1(new_n994), .A2(new_n998), .B1(KEYINPUT60), .B2(new_n990), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT61), .ZN(new_n1000));
  INV_X1    g575(.A(new_n987), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n992), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n823), .A2(KEYINPUT121), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n970), .B1(new_n937), .B2(new_n940), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n943), .A2(new_n1006), .A3(new_n974), .A4(new_n975), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(G1996), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT58), .B(G1341), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n974), .B2(new_n981), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT59), .B(new_n1003), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n999), .A2(new_n1002), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n987), .B1(new_n992), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n977), .A2(new_n979), .A3(new_n986), .A4(KEYINPUT122), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(KEYINPUT61), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n993), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2084), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n980), .A2(new_n1021), .A3(new_n974), .A4(new_n983), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1966), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1004), .A2(new_n974), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n969), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n995), .A2(KEYINPUT119), .A3(new_n1021), .A4(new_n983), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1024), .A2(G168), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(KEYINPUT123), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT123), .B(KEYINPUT51), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(G8), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1024), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1027), .ZN(new_n1037));
  OAI211_X1 g612(.A(G8), .B(G286), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1026), .A2(new_n969), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n776), .ZN(new_n1041));
  INV_X1    g616(.A(G1961), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n984), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1007), .A2(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n972), .A2(new_n1045), .A3(new_n974), .A4(new_n975), .ZN(new_n1046));
  AOI21_X1  g621(.A(G2078), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1041), .B(new_n1043), .C1(new_n1047), .C2(KEYINPUT53), .ZN(new_n1048));
  XOR2_X1   g623(.A(G171), .B(KEYINPUT54), .Z(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n972), .A2(new_n975), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n776), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1054));
  NOR4_X1   g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n476), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1049), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1043), .B(new_n1056), .C1(new_n1047), .C2(KEYINPUT53), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1039), .A2(new_n1050), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n988), .B2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1060), .B(new_n1061), .C1(new_n974), .C2(new_n981), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n691), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1064), .B(new_n1065), .C1(new_n691), .C2(G288), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT117), .B(G1981), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n681), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n681), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1064), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1063), .B1(G1976), .B2(new_n688), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1066), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1971), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1044), .A2(new_n1078), .A3(new_n1046), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n984), .A2(G2090), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1079), .A2(KEYINPUT115), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT115), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1061), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G303), .A2(G8), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT55), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1077), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1085), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1061), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT118), .B1(new_n1092), .B2(new_n1086), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1020), .A2(new_n1058), .A3(new_n1087), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1048), .A2(G171), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1039), .B2(KEYINPUT62), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1033), .A2(new_n1098), .A3(new_n1035), .A4(new_n1038), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1087), .A2(new_n1097), .A3(new_n1094), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1088), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1079), .A2(KEYINPUT115), .A3(new_n1080), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(G8), .A3(new_n1086), .A4(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1077), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1074), .A2(new_n691), .A3(new_n688), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1063), .B1(new_n1106), .B2(new_n1068), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1095), .A2(new_n1100), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1077), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1104), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1082), .A2(new_n1061), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1086), .B1(new_n1112), .B2(new_n1103), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n1061), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1111), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1090), .B1(new_n1089), .B2(new_n1085), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1092), .A2(KEYINPUT118), .A3(new_n1086), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1110), .B(new_n1104), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1115), .A2(G168), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT120), .B(new_n1118), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1109), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(G290), .A2(G1986), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n966), .B1(new_n947), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT112), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n965), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n968), .B1(new_n1127), .B2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g707(.A1(G227), .A2(new_n460), .ZN(new_n1134));
  OAI21_X1  g708(.A(new_n1134), .B1(new_n642), .B2(new_n643), .ZN(new_n1135));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n1136));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g711(.A(KEYINPUT126), .B(new_n1134), .C1(new_n642), .C2(new_n643), .ZN(new_n1138));
  NAND3_X1  g712(.A1(new_n674), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g713(.A(new_n1139), .B1(new_n873), .B2(new_n874), .ZN(new_n1140));
  AND3_X1   g714(.A1(new_n1140), .A2(new_n929), .A3(new_n932), .ZN(G308));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n929), .A3(new_n932), .ZN(G225));
endmodule


