//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n212));
  AOI21_X1  g011(.A(G190gat), .B1(new_n212), .B2(KEYINPUT64), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT28), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  NOR4_X1   g014(.A1(new_n208), .A2(new_n210), .A3(new_n215), .A4(G190gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n217), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n218), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n219), .B1(new_n218), .B2(new_n224), .ZN(new_n226));
  OAI22_X1  g025(.A1(new_n214), .A2(new_n216), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  AND2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n229), .A2(new_n230), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n220), .A3(new_n221), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n209), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT24), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n231), .A2(new_n235), .A3(new_n239), .A4(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n207), .A2(G183gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT64), .B1(new_n212), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(new_n207), .B2(G183gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n236), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n215), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n208), .A2(new_n210), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT28), .A3(new_n236), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT26), .ZN(new_n253));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n238), .B(new_n253), .C1(new_n256), .C2(new_n217), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n218), .A2(new_n224), .A3(new_n219), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n252), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n228), .A2(new_n244), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G134gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G127gat), .ZN(new_n265));
  INV_X1    g064(.A(G127gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G134gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(KEYINPUT1), .ZN(new_n270));
  INV_X1    g069(.A(G120gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G113gat), .ZN(new_n272));
  INV_X1    g071(.A(G113gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n270), .A2(new_n278), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n228), .A2(new_n281), .A3(new_n244), .A4(new_n262), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n205), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n204), .B1(new_n283), .B2(KEYINPUT33), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT32), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n282), .ZN(new_n288));
  INV_X1    g087(.A(new_n205), .ZN(new_n289));
  AOI221_X4 g088(.A(new_n285), .B1(KEYINPUT33), .B2(new_n204), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n280), .A2(new_n205), .A3(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT34), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n280), .A2(new_n293), .A3(new_n205), .A4(new_n282), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  OAI22_X1  g095(.A1(new_n287), .A2(new_n290), .B1(new_n296), .B2(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n288), .A2(new_n289), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n301), .A3(new_n204), .ZN(new_n302));
  INV_X1    g101(.A(new_n290), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT67), .B1(new_n292), .B2(new_n294), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT31), .B(G50gat), .ZN(new_n307));
  INV_X1    g106(.A(G106gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G228gat), .ZN(new_n311));
  INV_X1    g110(.A(G233gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316));
  INV_X1    g115(.A(G211gat), .ZN(new_n317));
  INV_X1    g116(.A(G218gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G211gat), .B(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n315), .A3(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(KEYINPUT71), .A2(G155gat), .A3(G162gat), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G141gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n326), .A2(KEYINPUT2), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT72), .B1(new_n334), .B2(new_n336), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n332), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(KEYINPUT74), .A2(G155gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT74), .A2(G155gat), .ZN(new_n343));
  OAI21_X1  g142(.A(G162gat), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT2), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n335), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(G141gat), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n334), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n331), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n326), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n345), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n341), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n325), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n336), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n338), .A3(new_n337), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n349), .A2(new_n334), .B1(new_n326), .B2(new_n351), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n361), .A2(new_n332), .B1(new_n362), .B2(new_n345), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT3), .B1(new_n325), .B2(new_n356), .ZN(new_n364));
  OAI22_X1  g163(.A1(new_n357), .A2(KEYINPUT80), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n357), .A2(KEYINPUT80), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n314), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n323), .A2(new_n324), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n354), .B1(new_n368), .B2(KEYINPUT29), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n341), .A2(new_n353), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n314), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n357), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT81), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n313), .B1(new_n364), .B2(new_n363), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n357), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G22gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n367), .B2(new_n377), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n380), .A2(G78gat), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G78gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n377), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G22gat), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n385), .B2(new_n379), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n310), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(G78gat), .B1(new_n380), .B2(new_n381), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n383), .A3(new_n379), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n309), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n306), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n392));
  XOR2_X1   g191(.A(G1gat), .B(G29gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT0), .ZN(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n370), .A2(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n279), .A3(new_n355), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n281), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n281), .A2(new_n341), .A3(new_n353), .ZN(new_n401));
  XOR2_X1   g200(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n370), .A2(new_n279), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n401), .ZN(new_n407));
  INV_X1    g206(.A(new_n399), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT76), .B(new_n399), .C1(new_n406), .C2(new_n401), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n404), .B(KEYINPUT5), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n355), .A2(new_n279), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n354), .B1(new_n341), .B2(new_n353), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(new_n399), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n363), .A2(new_n281), .A3(new_n402), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n401), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n396), .B1(new_n411), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n396), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n416), .B2(new_n422), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n429), .B2(KEYINPUT78), .ZN(new_n430));
  AOI211_X1 g229(.A(KEYINPUT78), .B(KEYINPUT6), .C1(new_n411), .C2(new_n426), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n430), .A2(new_n432), .B1(KEYINPUT6), .B2(new_n424), .ZN(new_n433));
  XNOR2_X1  g232(.A(G8gat), .B(G36gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n262), .A2(new_n244), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n261), .B1(new_n252), .B2(new_n260), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n356), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G226gat), .A2(G233gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT69), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n227), .A2(new_n244), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI211_X1 g245(.A(KEYINPUT69), .B(new_n441), .C1(new_n227), .C2(new_n244), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n325), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n228), .A2(new_n445), .A3(new_n244), .A4(new_n262), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n356), .A3(new_n441), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n368), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n437), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n445), .B1(new_n263), .B2(new_n356), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n252), .A2(new_n260), .B1(new_n242), .B2(new_n243), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT69), .B1(new_n455), .B2(new_n441), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n444), .A2(new_n443), .A3(new_n445), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n368), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n452), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(KEYINPUT30), .A3(new_n460), .A4(new_n436), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT70), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n460), .A3(new_n436), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n453), .A2(new_n467), .A3(new_n461), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n392), .B1(new_n433), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n466), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n467), .B1(new_n453), .B2(new_n461), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n424), .A2(KEYINPUT6), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n409), .A2(new_n410), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n399), .B1(new_n413), .B2(new_n414), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n403), .A2(new_n400), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT5), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n423), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n425), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT6), .B1(new_n411), .B2(new_n426), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n474), .B1(new_n483), .B2(new_n431), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n473), .A2(KEYINPUT79), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n391), .A2(new_n470), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n453), .A3(new_n461), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n396), .B(KEYINPUT82), .Z(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n479), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n481), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT35), .B1(new_n493), .B2(new_n474), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n387), .A2(new_n489), .A3(new_n390), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n302), .A2(new_n303), .A3(new_n296), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT68), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n295), .B1(new_n287), .B2(new_n290), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n302), .A2(new_n499), .A3(new_n303), .A4(new_n296), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n387), .A2(new_n390), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n468), .A2(new_n466), .ZN(new_n506));
  AND4_X1   g305(.A1(KEYINPUT79), .A2(new_n484), .A3(new_n463), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT79), .B1(new_n473), .B2(new_n484), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n399), .B1(new_n422), .B2(new_n398), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT39), .B1(new_n407), .B2(new_n408), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n421), .A2(new_n420), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT77), .B1(new_n401), .B2(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n398), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT39), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n408), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n490), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n520), .A3(new_n490), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n512), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n492), .B(new_n488), .C1(new_n522), .C2(KEYINPUT40), .ZN(new_n523));
  INV_X1    g322(.A(new_n512), .ZN(new_n524));
  INV_X1    g323(.A(new_n521), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n520), .B1(new_n517), .B2(new_n490), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n524), .B(KEYINPUT40), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT84), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n387), .A2(new_n390), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n459), .A2(new_n460), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n437), .B1(new_n531), .B2(KEYINPUT37), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT37), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n459), .B2(new_n460), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT38), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT87), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n532), .A2(KEYINPUT38), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n450), .A2(new_n368), .A3(new_n451), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n454), .A2(new_n458), .A3(new_n368), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(KEYINPUT85), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT37), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n493), .A2(new_n474), .A3(new_n464), .ZN(new_n547));
  OAI211_X1 g346(.A(KEYINPUT87), .B(KEYINPUT38), .C1(new_n532), .C2(new_n534), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n537), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n453), .A2(new_n461), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n550), .A2(new_n466), .B1(new_n479), .B2(new_n491), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT40), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT84), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n551), .A2(new_n554), .A3(new_n555), .A4(new_n527), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n529), .A2(new_n530), .A3(new_n549), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n306), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT36), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n497), .A2(new_n560), .A3(new_n498), .A4(new_n500), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n509), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n504), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NOR3_X1   g365(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n567));
  INV_X1    g366(.A(G29gat), .ZN(new_n568));
  INV_X1    g367(.A(G36gat), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n566), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G43gat), .B(G50gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT15), .A3(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(KEYINPUT15), .B2(new_n571), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT89), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n567), .A2(new_n575), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n566), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n572), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT90), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n579), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n585), .B(new_n589), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n590), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n582), .A2(new_n583), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n592), .B(new_n593), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT41), .ZN(new_n598));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n595), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT97), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n598), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT95), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n603), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n603), .A2(new_n609), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G57gat), .B(G64gat), .Z(new_n614));
  INV_X1    g413(.A(G71gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n383), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(KEYINPUT9), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G71gat), .B(G78gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  XOR2_X1   g418(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n266), .ZN(new_n624));
  XNOR2_X1  g423(.A(G15gat), .B(G22gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(G1gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(G8gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT16), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n625), .B1(new_n629), .B2(G1gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT92), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n627), .A2(KEYINPUT91), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT91), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n630), .B1(new_n626), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(G8gat), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT93), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n617), .B(new_n618), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(KEYINPUT21), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n624), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G155gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n641), .B(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n613), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n594), .A2(new_n619), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT10), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n596), .A2(new_n639), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n594), .A2(new_n619), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n649), .A2(KEYINPUT10), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT99), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n648), .B(new_n651), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n654), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(G230gat), .A3(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n647), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n638), .A2(new_n580), .ZN(new_n670));
  NAND2_X1  g469(.A1(G229gat), .A2(G233gat), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n582), .A2(new_n636), .A3(new_n632), .A4(new_n583), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT93), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n637), .B(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n580), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n670), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n671), .B(KEYINPUT13), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n670), .A2(KEYINPUT18), .A3(new_n671), .A4(new_n672), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n675), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G113gat), .B(G141gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(G169gat), .B(G197gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT12), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n682), .A3(new_n683), .A4(new_n690), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n669), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n564), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n484), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(G1gat), .Z(G1324gat));
  INV_X1    g498(.A(new_n697), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n628), .B1(new_n700), .B2(new_n488), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT16), .B(G8gat), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n697), .A2(new_n489), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT42), .B2(new_n703), .ZN(G1325gat));
  OAI21_X1  g504(.A(G15gat), .B1(new_n697), .B2(new_n562), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n501), .A2(G15gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n697), .B2(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n697), .A2(new_n530), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(new_n613), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n504), .B2(new_n563), .ZN(new_n713));
  INV_X1    g512(.A(new_n646), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(new_n695), .A3(new_n667), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n568), .A3(new_n433), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n720));
  AND3_X1   g519(.A1(new_n509), .A2(new_n557), .A3(new_n562), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n502), .B1(new_n486), .B2(KEYINPUT35), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n613), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n723), .B(new_n715), .C1(new_n713), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT101), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n613), .B1(new_n721), .B2(new_n722), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n724), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n729), .A2(new_n730), .A3(new_n723), .A4(new_n715), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n727), .A2(new_n433), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n719), .B1(new_n568), .B2(new_n732), .ZN(G1328gat));
  NOR3_X1   g532(.A1(new_n716), .A2(G36gat), .A3(new_n489), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n727), .A2(new_n488), .A3(new_n731), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n569), .ZN(G1329gat));
  NOR3_X1   g536(.A1(new_n716), .A2(G43gat), .A3(new_n501), .ZN(new_n738));
  INV_X1    g537(.A(new_n562), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n727), .A2(new_n739), .A3(new_n731), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(G43gat), .ZN(new_n741));
  INV_X1    g540(.A(G43gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n726), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n739), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n741), .A2(KEYINPUT47), .B1(new_n744), .B2(new_n746), .ZN(G1330gat));
  NOR3_X1   g546(.A1(new_n716), .A2(G50gat), .A3(new_n530), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G50gat), .B1(new_n726), .B2(new_n530), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT103), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n727), .A2(new_n505), .A3(new_n731), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n754), .A2(KEYINPUT102), .A3(G50gat), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT102), .B1(new_n754), .B2(G50gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n755), .A2(new_n756), .A3(new_n748), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n757), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g557(.A1(new_n564), .A2(new_n695), .A3(new_n647), .A4(new_n667), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT104), .Z(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n433), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT105), .B(G57gat), .Z(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1332gat));
  AOI21_X1  g562(.A(new_n489), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n760), .B(new_n764), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(G1333gat));
  INV_X1    g571(.A(new_n501), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n760), .A2(new_n615), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n760), .A2(new_n739), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n615), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(KEYINPUT50), .B(new_n774), .C1(new_n775), .C2(new_n615), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n505), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT108), .B(G78gat), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n695), .A2(new_n646), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT109), .Z(new_n785));
  NAND4_X1  g584(.A1(new_n729), .A2(new_n667), .A3(new_n723), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n484), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n713), .A2(new_n785), .ZN(new_n788));
  AND2_X1   g587(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n788), .B2(new_n790), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n433), .A2(new_n587), .A3(new_n667), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  OAI21_X1  g594(.A(G92gat), .B1(new_n786), .B2(new_n489), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n667), .A2(new_n588), .A3(new_n488), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT111), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n788), .B1(KEYINPUT112), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n713), .B2(new_n785), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n797), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n793), .B2(new_n799), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n806), .A2(new_n807), .B1(new_n797), .B2(new_n808), .ZN(G1337gat));
  XOR2_X1   g608(.A(KEYINPUT113), .B(G99gat), .Z(new_n810));
  NAND3_X1  g609(.A1(new_n773), .A2(new_n667), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT114), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n786), .A2(new_n562), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n793), .A2(new_n812), .B1(new_n813), .B2(new_n810), .ZN(G1338gat));
  NOR3_X1   g613(.A1(new_n530), .A2(G106gat), .A3(new_n668), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n792), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G106gat), .B1(new_n786), .B2(new_n530), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n815), .B1(new_n802), .B2(new_n804), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n817), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT115), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n817), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n820), .A2(new_n817), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(new_n819), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1339gat));
  NOR2_X1   g626(.A1(new_n484), .A2(new_n488), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  OAI211_X1 g629(.A(KEYINPUT99), .B(new_n656), .C1(new_n659), .C2(KEYINPUT10), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n648), .A4(new_n651), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n658), .A2(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n648), .B1(new_n831), .B2(new_n651), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n664), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n665), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n835), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n658), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n833), .A2(new_n664), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT55), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n830), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n841), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n836), .A2(new_n837), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT116), .A4(new_n665), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n694), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n680), .A2(new_n681), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n671), .B1(new_n670), .B2(new_n672), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n689), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n693), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n667), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n613), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  AND4_X1   g652(.A1(new_n613), .A2(new_n851), .A3(new_n843), .A4(new_n846), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n646), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n647), .A2(new_n695), .A3(new_n668), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n829), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n391), .ZN(new_n858));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n694), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n773), .A2(new_n530), .A3(new_n828), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n855), .B2(new_n856), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n695), .A2(new_n273), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(G1340gat));
  AOI21_X1  g662(.A(new_n271), .B1(new_n861), .B2(new_n667), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT117), .Z(new_n865));
  NAND3_X1  g664(.A1(new_n858), .A2(new_n271), .A3(new_n667), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(G1341gat));
  NAND3_X1  g668(.A1(new_n858), .A2(new_n266), .A3(new_n714), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n861), .A2(new_n714), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n266), .ZN(G1342gat));
  NAND3_X1  g671(.A1(new_n858), .A2(new_n264), .A3(new_n613), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT56), .Z(new_n874));
  AOI21_X1  g673(.A(new_n264), .B1(new_n861), .B2(new_n613), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT119), .Z(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n739), .A2(new_n829), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n838), .A2(new_n842), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n852), .B1(new_n695), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n712), .ZN(new_n882));
  INV_X1    g681(.A(new_n854), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n714), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n856), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT57), .B(new_n505), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n855), .A2(new_n856), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n505), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT120), .B(KEYINPUT57), .C1(new_n887), .C2(new_n505), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n694), .B(new_n878), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n857), .A2(new_n505), .A3(new_n562), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n333), .A3(new_n694), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n893), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n347), .A2(new_n348), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n668), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n505), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT57), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n530), .A2(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n613), .A2(new_n851), .A3(new_n879), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n714), .B1(new_n882), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n909), .B2(new_n885), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(new_n667), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n335), .B1(new_n912), .B2(new_n878), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n904), .B1(new_n901), .B2(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n894), .A2(new_n347), .A3(new_n348), .A4(new_n667), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1345gat));
  INV_X1    g715(.A(new_n903), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n342), .A2(new_n343), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n646), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n894), .A2(new_n714), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n917), .A2(new_n920), .B1(new_n918), .B2(new_n921), .ZN(G1346gat));
  NAND3_X1  g721(.A1(new_n894), .A2(new_n331), .A3(new_n613), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n903), .B2(new_n712), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G162gat), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n903), .A2(new_n924), .A3(new_n712), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n433), .A2(new_n489), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n887), .A2(new_n530), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n558), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n694), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n930), .A2(new_n501), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n695), .A2(new_n220), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  NOR4_X1   g734(.A1(new_n930), .A2(new_n221), .A3(new_n501), .A4(new_n668), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n931), .A2(new_n667), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n221), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT123), .ZN(G1349gat));
  NAND3_X1  g738(.A1(new_n931), .A2(new_n250), .A3(new_n714), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n930), .A2(new_n501), .A3(new_n646), .ZN(new_n943));
  OAI221_X1 g742(.A(new_n940), .B1(new_n941), .B2(new_n942), .C1(new_n209), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(G1350gat));
  AOI21_X1  g745(.A(new_n236), .B1(new_n933), .B2(new_n613), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT61), .Z(new_n948));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n236), .A3(new_n613), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1351gat));
  NAND2_X1  g749(.A1(new_n562), .A2(new_n929), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n906), .A2(new_n910), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n694), .A2(G197gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n905), .A2(new_n695), .A3(new_n951), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n953), .A2(new_n954), .B1(G197gat), .B2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n905), .A2(new_n951), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  AOI21_X1  g758(.A(G204gat), .B1(new_n959), .B2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n667), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n911), .B2(new_n951), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n911), .A2(new_n964), .A3(new_n951), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n958), .A2(new_n317), .A3(new_n714), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n953), .A2(new_n646), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  OAI21_X1  g773(.A(G218gat), .B1(new_n953), .B2(new_n712), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n318), .A3(new_n613), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n977), .B(new_n978), .ZN(G1355gat));
endmodule


