//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n190), .A3(G104), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(KEYINPUT78), .A3(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n193), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G101), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT79), .B(G101), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n198), .B(KEYINPUT4), .C1(new_n200), .C2(new_n197), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G116), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT2), .B(G113), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n197), .A2(new_n209), .A3(G101), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n201), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  AND4_X1   g025(.A1(new_n191), .A2(new_n193), .A3(new_n195), .A4(new_n196), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n192), .A2(G107), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n192), .A2(KEYINPUT81), .A3(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT81), .B1(new_n192), .B2(G107), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n212), .A2(new_n199), .B1(new_n217), .B2(G101), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT5), .ZN(new_n219));
  OAI21_X1  g033(.A(G113), .B1(new_n203), .B2(KEYINPUT5), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n219), .A2(new_n220), .B1(new_n206), .B2(new_n207), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G110), .B(G122), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT86), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n226), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n211), .A2(new_n228), .A3(new_n223), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(KEYINPUT6), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n231), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G125), .ZN(new_n242));
  INV_X1    g056(.A(G125), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n234), .A2(new_n236), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n243), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G224), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(G953), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n250), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n254));
  AND4_X1   g068(.A1(KEYINPUT87), .A2(new_n224), .A3(new_n254), .A4(new_n226), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n228), .B1(new_n211), .B2(new_n223), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT87), .B1(new_n256), .B2(new_n254), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n230), .B(new_n253), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT7), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(KEYINPUT90), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n250), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n260), .ZN(new_n263));
  OAI221_X1 g077(.A(new_n263), .B1(KEYINPUT90), .B2(new_n259), .C1(new_n242), .C2(new_n249), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n208), .A2(new_n210), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n265), .A2(new_n201), .B1(new_n218), .B2(new_n222), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n262), .A2(new_n264), .B1(new_n266), .B2(new_n228), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT88), .B(KEYINPUT8), .Z(new_n268));
  XNOR2_X1  g082(.A(new_n226), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n223), .A2(KEYINPUT89), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n218), .B2(new_n222), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n223), .A2(KEYINPUT89), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(G902), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n258), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(G210), .B1(G237), .B2(G902), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n258), .A2(new_n274), .A3(new_n276), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n188), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT9), .B(G234), .ZN(new_n281));
  OAI21_X1  g095(.A(G221), .B1(new_n281), .B2(G902), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n190), .B2(G104), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n192), .A2(KEYINPUT81), .A3(G107), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n213), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G101), .ZN(new_n287));
  OAI22_X1  g101(.A1(new_n197), .A2(new_n200), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n289), .A2(G128), .B1(new_n234), .B2(new_n236), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT10), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n289), .A2(KEYINPUT82), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n234), .A2(new_n295), .A3(KEYINPUT1), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n231), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n237), .B1(new_n297), .B2(new_n239), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n218), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT11), .ZN(new_n302));
  INV_X1    g116(.A(G134), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(G137), .ZN(new_n304));
  INV_X1    g118(.A(G137), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT11), .A3(G134), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(G137), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G131), .ZN(new_n309));
  INV_X1    g123(.A(G131), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n304), .A2(new_n306), .A3(new_n310), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n197), .A2(G101), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT4), .B1(new_n197), .B2(new_n200), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n246), .A2(new_n248), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n210), .A2(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n210), .A2(new_n318), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT80), .B1(new_n321), .B2(new_n201), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n301), .B(new_n313), .C1(new_n320), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT84), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n317), .B1(new_n316), .B2(new_n319), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n201), .A3(KEYINPUT80), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n324), .B(new_n313), .C1(new_n327), .C2(new_n301), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n301), .B1(new_n320), .B2(new_n322), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT84), .B1(new_n329), .B2(new_n312), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n323), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G140), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G227), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n288), .A2(new_n241), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n313), .B1(new_n299), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n313), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n339), .A2(new_n342), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n323), .B(new_n335), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT85), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n339), .B(new_n342), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n348), .A2(KEYINPUT85), .A3(new_n323), .A4(new_n335), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI211_X1 g164(.A(G469), .B(G902), .C1(new_n337), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G469), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n323), .B(new_n335), .C1(new_n328), .C2(new_n330), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n323), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n335), .B(KEYINPUT77), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G902), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n352), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n280), .B(new_n282), .C1(new_n351), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n235), .A2(G128), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n231), .A2(G143), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n303), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G116), .B(G122), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n190), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n204), .A2(G122), .ZN(new_n367));
  INV_X1    g181(.A(G122), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G116), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n364), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(new_n361), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n362), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n376), .B2(new_n361), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n372), .B1(new_n377), .B2(new_n303), .ZN(new_n378));
  INV_X1    g192(.A(G217), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n281), .A2(new_n379), .A3(G953), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n231), .A2(G143), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n235), .A2(G128), .ZN(new_n382));
  OAI21_X1  g196(.A(G134), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n383), .A2(new_n363), .B1(new_n190), .B2(new_n365), .ZN(new_n384));
  OAI211_X1 g198(.A(KEYINPUT93), .B(KEYINPUT14), .C1(new_n368), .C2(G116), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n204), .A3(G122), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n369), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT93), .B1(new_n367), .B2(KEYINPUT14), .ZN(new_n389));
  OAI21_X1  g203(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n384), .A2(new_n390), .A3(KEYINPUT94), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT94), .B1(new_n384), .B2(new_n390), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n378), .B(new_n380), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n385), .A2(new_n369), .A3(new_n387), .ZN(new_n397));
  INV_X1    g211(.A(new_n389), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n190), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n303), .B1(new_n361), .B2(new_n362), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n366), .B1(new_n364), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n384), .A2(new_n390), .A3(KEYINPUT94), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(KEYINPUT95), .A3(new_n378), .A4(new_n380), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n378), .B1(new_n391), .B2(new_n392), .ZN(new_n406));
  INV_X1    g220(.A(new_n380), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n395), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n358), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(KEYINPUT96), .A3(new_n358), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  AOI211_X1 g230(.A(KEYINPUT96), .B(new_n415), .C1(new_n409), .C2(new_n358), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G952), .ZN(new_n420));
  AOI211_X1 g234(.A(G953), .B(new_n420), .C1(G234), .C2(G237), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n358), .B(new_n333), .C1(G234), .C2(G237), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G237), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n333), .A3(G214), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n235), .ZN(new_n428));
  NOR2_X1   g242(.A1(G237), .A2(G953), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G143), .A3(G214), .ZN(new_n430));
  NAND2_X1  g244(.A1(KEYINPUT18), .A2(G131), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G140), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G125), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n243), .A2(G140), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G146), .ZN(new_n437));
  XNOR2_X1  g251(.A(G125), .B(G140), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n233), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n428), .A2(new_n430), .ZN(new_n441));
  INV_X1    g255(.A(new_n431), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(KEYINPUT91), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT91), .B1(new_n441), .B2(new_n442), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n432), .B(new_n440), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G113), .B(G122), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(new_n192), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT72), .B1(new_n243), .B2(G140), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT72), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n433), .A3(G125), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT16), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(KEYINPUT72), .A2(KEYINPUT16), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n434), .B2(new_n435), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n457), .A3(new_n233), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT16), .B1(new_n449), .B2(new_n451), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n461), .A2(new_n456), .A3(G146), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT73), .ZN(new_n463));
  OAI21_X1  g277(.A(G146), .B1(new_n461), .B2(new_n456), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n441), .A2(G131), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT17), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n428), .A2(new_n310), .A3(new_n430), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n441), .A2(KEYINPUT17), .A3(G131), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n446), .B(new_n448), .C1(new_n465), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n448), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n468), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n438), .A2(KEYINPUT19), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n438), .A2(KEYINPUT19), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n233), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n474), .A2(new_n477), .A3(new_n464), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n440), .A2(new_n432), .ZN(new_n479));
  INV_X1    g293(.A(new_n445), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n443), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n473), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(G475), .A2(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT20), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n487), .A3(new_n484), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n464), .B1(new_n462), .B2(KEYINPUT73), .ZN(new_n489));
  NOR4_X1   g303(.A1(new_n461), .A2(new_n456), .A3(new_n459), .A4(G146), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n471), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n448), .B1(new_n493), .B2(new_n446), .ZN(new_n494));
  INV_X1    g308(.A(new_n472), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n358), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n486), .A2(new_n488), .B1(new_n496), .B2(G475), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n419), .A2(new_n425), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n360), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT26), .B(G101), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n429), .A2(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n312), .A2(new_n318), .ZN(new_n506));
  INV_X1    g320(.A(new_n208), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n305), .A2(G134), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n307), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT65), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(G131), .ZN(new_n511));
  XNOR2_X1  g325(.A(G134), .B(G137), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT65), .B1(new_n512), .B2(new_n310), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n240), .A2(new_n311), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n506), .A2(new_n507), .A3(new_n514), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n506), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n309), .A2(new_n311), .B1(new_n246), .B2(new_n248), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT64), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n518), .B1(new_n523), .B2(new_n208), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n505), .B(new_n517), .C1(new_n524), .C2(new_n516), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n514), .B1(new_n521), .B2(KEYINPUT64), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n312), .A2(KEYINPUT64), .A3(new_n318), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n208), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n515), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT28), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(KEYINPUT68), .A3(new_n505), .A4(new_n517), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n520), .A2(new_n535), .A3(new_n514), .A4(new_n522), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n506), .A2(new_n514), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT30), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n507), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n504), .B1(new_n539), .B2(new_n518), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n527), .A2(new_n528), .A3(new_n534), .A4(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n507), .B1(new_n506), .B2(new_n514), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT28), .B1(new_n518), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n504), .A2(new_n528), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n517), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n358), .B1(new_n545), .B2(KEYINPUT69), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n545), .B2(KEYINPUT69), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G472), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n536), .A2(new_n538), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n208), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n505), .A3(new_n515), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT31), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n539), .A2(new_n504), .A3(new_n518), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n516), .B1(new_n531), .B2(new_n515), .ZN(new_n557));
  INV_X1    g371(.A(new_n517), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n504), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT32), .ZN(new_n561));
  NOR2_X1   g375(.A1(G472), .A2(G902), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT67), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n560), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n549), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT25), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT71), .B(KEYINPUT23), .C1(new_n231), .C2(G119), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n231), .B(G119), .C1(KEYINPUT71), .C2(KEYINPUT23), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT70), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n202), .B2(G128), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n231), .A2(KEYINPUT70), .A3(G119), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n202), .A2(G128), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT24), .B(G110), .Z(new_n578));
  AOI22_X1  g392(.A1(new_n572), .A2(G110), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n489), .B2(new_n490), .ZN(new_n580));
  OAI22_X1  g394(.A1(new_n572), .A2(G110), .B1(new_n577), .B2(new_n578), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n439), .A3(new_n464), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(KEYINPUT74), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT22), .B(G137), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT74), .B1(new_n580), .B2(new_n582), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n582), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT74), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n586), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n569), .B(new_n358), .C1(new_n590), .C2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n379), .B1(G234), .B2(new_n358), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n591), .A2(new_n592), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n587), .A3(new_n583), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n593), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n569), .B1(new_n600), .B2(new_n358), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT75), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n358), .B1(new_n590), .B2(new_n594), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT25), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n595), .A4(new_n596), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n596), .A2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT76), .B1(new_n568), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n559), .B1(new_n554), .B2(new_n555), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n552), .A2(KEYINPUT31), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n564), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT32), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n614), .A2(new_n565), .B1(G472), .B2(new_n548), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT76), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n499), .B1(new_n610), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n200), .ZN(G3));
  NAND3_X1  g434(.A1(new_n408), .A2(KEYINPUT33), .A3(new_n393), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n414), .A2(G902), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n409), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n623), .B1(new_n409), .B2(new_n624), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n621), .B(new_n622), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n410), .A2(new_n414), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n497), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n279), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n276), .B1(new_n258), .B2(new_n274), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n425), .B(new_n187), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT99), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n634), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n637), .A3(new_n630), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n560), .A2(new_n358), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(KEYINPUT97), .A3(G472), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n643), .A2(new_n644), .B1(new_n564), .B2(new_n560), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n282), .B1(new_n351), .B2(new_n359), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n616), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n639), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  NAND3_X1  g464(.A1(new_n647), .A2(new_n645), .A3(new_n636), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n413), .A2(new_n415), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT96), .B1(new_n409), .B2(new_n358), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n417), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n497), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n587), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n591), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n607), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n602), .A2(new_n606), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n602), .A2(new_n606), .A3(KEYINPUT100), .A4(new_n662), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n499), .A2(new_n667), .A3(new_n645), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n421), .B1(new_n422), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n655), .A2(KEYINPUT101), .A3(new_n497), .A4(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n416), .A2(new_n497), .A3(new_n418), .A4(new_n673), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n677), .A3(new_n280), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n646), .A2(new_n615), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n674), .A2(new_n677), .A3(KEYINPUT102), .A4(new_n280), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n680), .A2(new_n667), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  NOR2_X1   g498(.A1(new_n518), .A2(new_n542), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n505), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n358), .B1(new_n554), .B2(new_n686), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n614), .A2(new_n565), .B1(G472), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT103), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n667), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n419), .A2(new_n497), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n187), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n632), .A2(new_n633), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT38), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n672), .B(KEYINPUT39), .Z(new_n695));
  OAI211_X1 g509(.A(new_n282), .B(new_n695), .C1(new_n351), .C2(new_n359), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n692), .B(new_n694), .C1(KEYINPUT40), .C2(new_n696), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n690), .B(new_n697), .C1(KEYINPUT40), .C2(new_n696), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NOR2_X1   g513(.A1(new_n360), .A2(new_n615), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n630), .A2(new_n673), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n667), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  NOR2_X1   g518(.A1(new_n615), .A2(new_n616), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n331), .A2(new_n336), .B1(new_n347), .B2(new_n349), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n337), .A2(new_n350), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n352), .A3(new_n358), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n709), .A3(new_n282), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n639), .A2(new_n705), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NOR2_X1   g528(.A1(new_n656), .A2(new_n634), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n705), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND4_X1  g531(.A1(new_n707), .A2(new_n709), .A3(new_n280), .A4(new_n282), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n615), .A3(new_n498), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT104), .B1(new_n719), .B2(new_n667), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(KEYINPUT104), .A3(new_n667), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND2_X1  g538(.A1(new_n691), .A2(new_n280), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n710), .A2(new_n725), .A3(new_n424), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n543), .A2(new_n517), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n553), .B1(new_n505), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n564), .B1(new_n728), .B2(new_n612), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n641), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n616), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NOR2_X1   g547(.A1(new_n718), .A2(new_n701), .ZN(new_n734));
  INV_X1    g548(.A(new_n730), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n667), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n632), .A2(new_n188), .A3(new_n633), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n739), .B(new_n282), .C1(new_n351), .C2(new_n359), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n740), .A2(new_n615), .A3(new_n616), .A4(new_n701), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n740), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n705), .A3(new_n702), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NAND4_X1  g562(.A1(new_n744), .A2(new_n705), .A3(new_n677), .A4(new_n674), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n353), .A2(new_n752), .A3(new_n356), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n353), .B2(new_n356), .ZN(new_n754));
  OAI21_X1  g568(.A(G469), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT106), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n757), .B(G469), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(G469), .A2(G902), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n751), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n351), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n759), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n760), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n282), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n695), .ZN(new_n768));
  INV_X1    g582(.A(new_n739), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n665), .A2(new_n666), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n628), .A2(new_n629), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n497), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(KEYINPUT43), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(KEYINPUT43), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n770), .A2(new_n645), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n769), .B1(new_n775), .B2(KEYINPUT44), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(KEYINPUT44), .B2(new_n775), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n305), .ZN(G39));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n766), .A2(new_n282), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n783), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n766), .A2(new_n282), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n568), .A2(new_n609), .A3(new_n701), .A4(new_n769), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND3_X1  g604(.A1(new_n694), .A2(new_n187), .A3(new_n282), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n616), .A3(new_n772), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n707), .A2(new_n709), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT49), .Z(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n689), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n784), .B(new_n786), .C1(new_n282), .C2(new_n793), .ZN(new_n797));
  INV_X1    g611(.A(new_n421), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n773), .A2(new_n774), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n731), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n769), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT116), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n710), .A2(new_n616), .A3(new_n769), .A4(new_n798), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n689), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n497), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n771), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT119), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n710), .A2(new_n769), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n799), .A2(KEYINPUT118), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT118), .B1(new_n799), .B2(new_n811), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n667), .A3(new_n735), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n187), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n711), .A2(new_n694), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n800), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n816), .A2(new_n817), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n810), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n796), .B1(new_n803), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n800), .A2(new_n718), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n420), .A3(G953), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT48), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n814), .A2(new_n827), .A3(new_n705), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n814), .B2(new_n705), .ZN(new_n829));
  OAI221_X1 g643(.A(new_n826), .B1(new_n631), .B2(new_n805), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n823), .B1(new_n797), .B2(new_n802), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(KEYINPUT51), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n654), .A2(KEYINPUT110), .A3(new_n417), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n416), .B2(new_n418), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n497), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n621), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n409), .A2(new_n624), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT98), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(new_n625), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n842), .A2(new_n622), .B1(new_n414), .B2(new_n410), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT109), .B1(new_n843), .B2(new_n497), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT109), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n630), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n838), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n647), .A2(new_n847), .A3(new_n645), .A4(new_n636), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n619), .A2(new_n668), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT111), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n619), .A2(new_n848), .A3(new_n668), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OR3_X1    g667(.A1(new_n835), .A2(new_n837), .A3(new_n806), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n854), .A2(new_n615), .B1(new_n631), .B2(new_n730), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n667), .A3(new_n673), .A4(new_n744), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n746), .A2(new_n743), .A3(new_n749), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n712), .A2(new_n732), .A3(new_n716), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n722), .B2(new_n721), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n853), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n568), .A2(new_n609), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n710), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n864), .A2(new_n639), .B1(new_n726), .B2(new_n731), .ZN(new_n865));
  INV_X1    g679(.A(new_n722), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n865), .B(new_n716), .C1(new_n866), .C2(new_n720), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n852), .B2(new_n850), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(KEYINPUT112), .A3(new_n857), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n646), .A2(new_n725), .A3(new_n672), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n688), .A2(new_n663), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT113), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n683), .A2(new_n874), .A3(new_n736), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n683), .B2(new_n736), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n703), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n871), .A2(new_n872), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n683), .A2(new_n703), .A3(new_n736), .A4(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n862), .A2(new_n869), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n860), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n870), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n360), .A2(new_n615), .A3(new_n701), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n888), .A2(new_n667), .B1(new_n871), .B2(new_n872), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(KEYINPUT52), .A3(new_n683), .A4(new_n736), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n886), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n891), .A2(new_n853), .A3(new_n859), .A4(new_n857), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n884), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n834), .B1(new_n885), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n882), .A2(new_n868), .A3(KEYINPUT53), .A4(new_n857), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n884), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n899), .A3(new_n834), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n833), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n795), .B1(new_n902), .B2(new_n903), .ZN(G75));
  NOR2_X1   g718(.A1(new_n333), .A2(G952), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n358), .B1(new_n898), .B2(new_n899), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT56), .B1(new_n907), .B2(G210), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n230), .B1(new_n255), .B2(new_n257), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT120), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n253), .B(KEYINPUT55), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n906), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n908), .B2(new_n912), .ZN(G51));
  AOI21_X1  g728(.A(new_n834), .B1(new_n898), .B2(new_n899), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n901), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n760), .B(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n708), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n907), .A2(new_n758), .A3(new_n756), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n905), .B1(new_n918), .B2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  INV_X1    g735(.A(new_n483), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n905), .ZN(G60));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n842), .B(KEYINPUT121), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n926), .B(new_n906), .C1(new_n916), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n898), .A2(new_n899), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT54), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n934), .B2(new_n900), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT122), .B1(new_n935), .B2(new_n905), .ZN(new_n936));
  INV_X1    g750(.A(new_n929), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n897), .B2(new_n901), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n932), .A2(new_n936), .B1(new_n938), .B2(new_n927), .ZN(G63));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n379), .A2(new_n358), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n898), .B2(new_n899), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n940), .B(new_n906), .C1(new_n945), .C2(new_n600), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n894), .A2(new_n884), .ZN(new_n949));
  INV_X1    g763(.A(new_n881), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n683), .A2(new_n736), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT113), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n683), .A2(new_n874), .A3(new_n736), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n952), .A2(new_n953), .B1(new_n667), .B2(new_n888), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n954), .B2(new_n873), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n853), .A2(new_n857), .A3(KEYINPUT53), .A4(new_n859), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n943), .B1(new_n949), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n600), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n905), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND4_X1   g774(.A1(KEYINPUT124), .A2(new_n933), .A3(new_n661), .A4(new_n943), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT124), .B1(new_n945), .B2(new_n661), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n948), .A2(new_n963), .ZN(new_n964));
  OAI221_X1 g778(.A(new_n960), .B1(new_n940), .B2(KEYINPUT61), .C1(new_n961), .C2(new_n962), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(G66));
  NOR3_X1   g780(.A1(new_n423), .A2(new_n251), .A3(new_n333), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n868), .B2(new_n333), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n910), .B1(G898), .B2(new_n333), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G69));
  NAND3_X1  g784(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n954), .A2(new_n698), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n696), .A2(new_n769), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n847), .C1(new_n610), .C2(new_n618), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n778), .B1(new_n787), .B2(new_n788), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n971), .B1(new_n977), .B2(G953), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n475), .A2(new_n476), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n550), .B(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n954), .A2(new_n747), .A3(new_n749), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n863), .A2(new_n725), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n767), .A2(new_n695), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n333), .A3(new_n976), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n671), .A2(KEYINPUT127), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT127), .B1(new_n671), .B2(G227), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n333), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  AOI22_X1  g805(.A1(new_n978), .A2(new_n980), .B1(new_n987), .B2(new_n991), .ZN(G72));
  NOR2_X1   g806(.A1(new_n539), .A2(new_n518), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(new_n505), .ZN(new_n994));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n885), .B2(new_n896), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n906), .B1(new_n994), .B2(new_n996), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n993), .A2(new_n504), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n973), .A2(new_n975), .A3(new_n976), .A4(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n986), .A2(new_n504), .A3(new_n993), .A4(new_n976), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n998), .B(new_n999), .C1(new_n1003), .C2(new_n868), .ZN(G57));
endmodule


