

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(n694), .B(KEYINPUT103), .ZN(n695) );
  XOR2_X1 U555 ( .A(KEYINPUT1), .B(n524), .Z(n660) );
  NOR2_X2 U556 ( .A1(n556), .A2(n555), .ZN(G164) );
  XNOR2_X1 U557 ( .A(n548), .B(KEYINPUT65), .ZN(G160) );
  NOR2_X1 U558 ( .A1(n812), .A2(n523), .ZN(n521) );
  NOR2_X1 U559 ( .A1(n771), .A2(n770), .ZN(n522) );
  AND2_X1 U560 ( .A1(n811), .A2(n825), .ZN(n523) );
  INV_X1 U561 ( .A(KEYINPUT30), .ZN(n694) );
  INV_X1 U562 ( .A(KEYINPUT28), .ZN(n728) );
  XNOR2_X1 U563 ( .A(n696), .B(n695), .ZN(n697) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n702) );
  NOR2_X1 U565 ( .A1(G1966), .A2(n771), .ZN(n751) );
  NAND2_X1 U566 ( .A1(n794), .A2(n691), .ZN(n710) );
  AND2_X1 U567 ( .A1(n813), .A2(n521), .ZN(n815) );
  NOR2_X2 U568 ( .A1(G2105), .A2(n542), .ZN(n883) );
  NOR2_X1 U569 ( .A1(G651), .A2(n661), .ZN(n655) );
  XOR2_X1 U570 ( .A(KEYINPUT74), .B(n536), .Z(G299) );
  INV_X1 U571 ( .A(G651), .ZN(n529) );
  NOR2_X1 U572 ( .A1(G543), .A2(n529), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n660), .A2(G65), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n525), .B(KEYINPUT72), .ZN(n527) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n661) );
  NAND2_X1 U576 ( .A1(G53), .A2(n655), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U578 ( .A(n528), .B(KEYINPUT73), .ZN(n531) );
  NOR2_X1 U579 ( .A1(n661), .A2(n529), .ZN(n649) );
  NAND2_X1 U580 ( .A1(G78), .A2(n649), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n535) );
  NOR2_X1 U582 ( .A1(G543), .A2(G651), .ZN(n532) );
  XNOR2_X1 U583 ( .A(n532), .B(KEYINPUT64), .ZN(n646) );
  NAND2_X1 U584 ( .A1(G91), .A2(n646), .ZN(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT71), .B(n533), .ZN(n534) );
  NOR2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  INV_X1 U587 ( .A(G2105), .ZN(n539) );
  NOR2_X1 U588 ( .A1(n539), .A2(G2104), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n537), .B(KEYINPUT66), .ZN(n887) );
  NAND2_X1 U590 ( .A1(n887), .A2(G125), .ZN(n547) );
  NOR2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  XOR2_X2 U592 ( .A(KEYINPUT17), .B(n538), .Z(n884) );
  NAND2_X1 U593 ( .A1(G137), .A2(n884), .ZN(n541) );
  INV_X1 U594 ( .A(G2104), .ZN(n542) );
  NOR2_X1 U595 ( .A1(n542), .A2(n539), .ZN(n889) );
  NAND2_X1 U596 ( .A1(G113), .A2(n889), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G101), .A2(n883), .ZN(n543) );
  XNOR2_X1 U599 ( .A(KEYINPUT23), .B(n543), .ZN(n544) );
  NOR2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U602 ( .A1(G102), .A2(n883), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G138), .A2(n884), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U605 ( .A(KEYINPUT92), .B(n551), .Z(n553) );
  NAND2_X1 U606 ( .A1(G126), .A2(n887), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U608 ( .A1(G114), .A2(n889), .ZN(n554) );
  XNOR2_X1 U609 ( .A(KEYINPUT91), .B(n554), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G64), .A2(n660), .ZN(n558) );
  NAND2_X1 U611 ( .A1(G52), .A2(n655), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT69), .B(n559), .Z(n565) );
  NAND2_X1 U614 ( .A1(G90), .A2(n646), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n560), .B(KEYINPUT70), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G77), .A2(n649), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U619 ( .A1(n565), .A2(n564), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U621 ( .A1(G99), .A2(n883), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G111), .A2(n889), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U624 ( .A1(n887), .A2(G123), .ZN(n568) );
  XNOR2_X1 U625 ( .A(n568), .B(KEYINPUT18), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n884), .A2(G135), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U628 ( .A1(n572), .A2(n571), .ZN(n1000) );
  XNOR2_X1 U629 ( .A(n1000), .B(G2096), .ZN(n573) );
  XNOR2_X1 U630 ( .A(n573), .B(KEYINPUT83), .ZN(n574) );
  OR2_X1 U631 ( .A1(G2100), .A2(n574), .ZN(G156) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  NAND2_X1 U633 ( .A1(G75), .A2(n649), .ZN(n575) );
  XNOR2_X1 U634 ( .A(n575), .B(KEYINPUT86), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G88), .A2(n646), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G62), .A2(n660), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G50), .A2(n655), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U640 ( .A1(n581), .A2(n580), .ZN(G166) );
  NAND2_X1 U641 ( .A1(G89), .A2(n646), .ZN(n582) );
  XNOR2_X1 U642 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G76), .A2(n649), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U645 ( .A(KEYINPUT5), .B(n585), .ZN(n593) );
  NAND2_X1 U646 ( .A1(n655), .A2(G51), .ZN(n586) );
  XNOR2_X1 U647 ( .A(KEYINPUT79), .B(n586), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n660), .A2(G63), .ZN(n587) );
  XOR2_X1 U649 ( .A(n587), .B(KEYINPUT78), .Z(n588) );
  NOR2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U651 ( .A(KEYINPUT80), .B(n590), .Z(n591) );
  XOR2_X1 U652 ( .A(KEYINPUT6), .B(n591), .Z(n592) );
  NAND2_X1 U653 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U654 ( .A(KEYINPUT7), .B(n594), .ZN(G168) );
  XOR2_X1 U655 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n595) );
  XNOR2_X1 U657 ( .A(n595), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U658 ( .A(G223), .ZN(n830) );
  NAND2_X1 U659 ( .A1(n830), .A2(G567), .ZN(n596) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n596), .Z(G234) );
  NAND2_X1 U661 ( .A1(n646), .A2(G81), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n597), .B(KEYINPUT12), .ZN(n598) );
  XNOR2_X1 U663 ( .A(n598), .B(KEYINPUT76), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G68), .A2(n649), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U666 ( .A(KEYINPUT13), .B(n601), .Z(n605) );
  NAND2_X1 U667 ( .A1(G56), .A2(n660), .ZN(n602) );
  XNOR2_X1 U668 ( .A(n602), .B(KEYINPUT14), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n603), .B(KEYINPUT75), .ZN(n604) );
  NOR2_X1 U670 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U671 ( .A1(n655), .A2(G43), .ZN(n606) );
  NAND2_X1 U672 ( .A1(n607), .A2(n606), .ZN(n923) );
  INV_X1 U673 ( .A(n923), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n608), .A2(G860), .ZN(G153) );
  INV_X1 U675 ( .A(G171), .ZN(G301) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n618) );
  NAND2_X1 U677 ( .A1(n649), .A2(G79), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G92), .A2(n646), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U680 ( .A1(G66), .A2(n660), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G54), .A2(n655), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n616) );
  XNOR2_X1 U684 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n616), .B(n615), .ZN(n922) );
  OR2_X1 U686 ( .A1(n922), .A2(G868), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n618), .A2(n617), .ZN(G284) );
  INV_X1 U688 ( .A(G868), .ZN(n664) );
  NOR2_X1 U689 ( .A1(G286), .A2(n664), .ZN(n620) );
  NOR2_X1 U690 ( .A1(G299), .A2(G868), .ZN(n619) );
  NOR2_X1 U691 ( .A1(n620), .A2(n619), .ZN(G297) );
  INV_X1 U692 ( .A(G559), .ZN(n621) );
  NOR2_X1 U693 ( .A1(G860), .A2(n621), .ZN(n622) );
  XNOR2_X1 U694 ( .A(KEYINPUT81), .B(n622), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n623), .A2(n922), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n624), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G868), .A2(n923), .ZN(n625) );
  XNOR2_X1 U698 ( .A(KEYINPUT82), .B(n625), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G868), .A2(n922), .ZN(n626) );
  NOR2_X1 U700 ( .A1(G559), .A2(n626), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U702 ( .A1(G559), .A2(n922), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n629), .B(n923), .ZN(n673) );
  NOR2_X1 U704 ( .A1(G860), .A2(n673), .ZN(n637) );
  NAND2_X1 U705 ( .A1(G67), .A2(n660), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G55), .A2(n655), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n649), .A2(G80), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G93), .A2(n646), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n666) );
  XOR2_X1 U712 ( .A(n666), .B(KEYINPUT84), .Z(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(G145) );
  NAND2_X1 U714 ( .A1(G60), .A2(n660), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G47), .A2(n655), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U717 ( .A(KEYINPUT68), .B(n640), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G85), .A2(n646), .ZN(n641) );
  XNOR2_X1 U719 ( .A(KEYINPUT67), .B(n641), .ZN(n642) );
  NOR2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n649), .A2(G72), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U723 ( .A1(G61), .A2(n660), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G86), .A2(n646), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n649), .A2(G73), .ZN(n650) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(G48), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G49), .A2(n655), .ZN(n657) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U734 ( .A(KEYINPUT85), .B(n658), .Z(n659) );
  NOR2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n661), .A2(G87), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n663), .A2(n662), .ZN(G288) );
  NAND2_X1 U738 ( .A1(n664), .A2(n666), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n665), .B(KEYINPUT88), .ZN(n676) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n667) );
  XOR2_X1 U741 ( .A(n667), .B(n666), .Z(n668) );
  XNOR2_X1 U742 ( .A(n668), .B(G290), .ZN(n671) );
  XNOR2_X1 U743 ( .A(G166), .B(G299), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n669), .B(G305), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n672), .B(G288), .ZN(n901) );
  XNOR2_X1 U747 ( .A(n901), .B(n673), .ZN(n674) );
  NAND2_X1 U748 ( .A1(G868), .A2(n674), .ZN(n675) );
  NAND2_X1 U749 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U754 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n682) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U759 ( .A1(n683), .A2(G218), .ZN(n684) );
  NAND2_X1 U760 ( .A1(G96), .A2(n684), .ZN(n836) );
  NAND2_X1 U761 ( .A1(n836), .A2(G2106), .ZN(n689) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U763 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U764 ( .A1(G108), .A2(n686), .ZN(n835) );
  NAND2_X1 U765 ( .A1(G567), .A2(n835), .ZN(n687) );
  XNOR2_X1 U766 ( .A(KEYINPUT90), .B(n687), .ZN(n688) );
  NAND2_X1 U767 ( .A1(n689), .A2(n688), .ZN(n837) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n690) );
  NOR2_X1 U769 ( .A1(n837), .A2(n690), .ZN(n834) );
  NAND2_X1 U770 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U771 ( .A(G166), .ZN(G303) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n793) );
  INV_X1 U774 ( .A(n793), .ZN(n691) );
  NAND2_X1 U775 ( .A1(G8), .A2(n710), .ZN(n771) );
  NOR2_X1 U776 ( .A1(G2084), .A2(n710), .ZN(n747) );
  NOR2_X1 U777 ( .A1(n751), .A2(n747), .ZN(n692) );
  XNOR2_X1 U778 ( .A(n692), .B(KEYINPUT102), .ZN(n693) );
  NAND2_X1 U779 ( .A1(n693), .A2(G8), .ZN(n696) );
  NOR2_X1 U780 ( .A1(G168), .A2(n697), .ZN(n701) );
  XNOR2_X1 U781 ( .A(KEYINPUT25), .B(G2078), .ZN(n986) );
  NOR2_X1 U782 ( .A1(n710), .A2(n986), .ZN(n699) );
  AND2_X1 U783 ( .A1(n710), .A2(G1961), .ZN(n698) );
  NOR2_X1 U784 ( .A1(n699), .A2(n698), .ZN(n704) );
  NOR2_X1 U785 ( .A1(G171), .A2(n704), .ZN(n700) );
  NOR2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n703) );
  XNOR2_X1 U787 ( .A(n703), .B(n702), .ZN(n748) );
  NAND2_X1 U788 ( .A1(G171), .A2(n704), .ZN(n734) );
  INV_X1 U789 ( .A(KEYINPUT101), .ZN(n719) );
  INV_X1 U790 ( .A(G1996), .ZN(n983) );
  NOR2_X1 U791 ( .A1(n710), .A2(n983), .ZN(n705) );
  XOR2_X1 U792 ( .A(n705), .B(KEYINPUT26), .Z(n708) );
  AND2_X1 U793 ( .A1(n710), .A2(G1341), .ZN(n706) );
  NOR2_X1 U794 ( .A1(n706), .A2(n923), .ZN(n707) );
  AND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n709) );
  OR2_X1 U796 ( .A1(n922), .A2(n709), .ZN(n717) );
  NAND2_X1 U797 ( .A1(n709), .A2(n922), .ZN(n715) );
  INV_X1 U798 ( .A(n710), .ZN(n721) );
  AND2_X1 U799 ( .A1(n721), .A2(G2067), .ZN(n711) );
  XOR2_X1 U800 ( .A(n711), .B(KEYINPUT100), .Z(n713) );
  NAND2_X1 U801 ( .A1(n710), .A2(G1348), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U805 ( .A(n719), .B(n718), .ZN(n725) );
  NAND2_X1 U806 ( .A1(n721), .A2(G2072), .ZN(n720) );
  XNOR2_X1 U807 ( .A(n720), .B(KEYINPUT27), .ZN(n723) );
  INV_X1 U808 ( .A(G1956), .ZN(n952) );
  NOR2_X1 U809 ( .A1(n952), .A2(n721), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n727) );
  INV_X1 U811 ( .A(G299), .ZN(n726) );
  NAND2_X1 U812 ( .A1(n727), .A2(n726), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n731) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U815 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U817 ( .A(KEYINPUT29), .B(n732), .Z(n733) );
  NAND2_X1 U818 ( .A1(n734), .A2(n733), .ZN(n749) );
  INV_X1 U819 ( .A(G8), .ZN(n740) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n771), .ZN(n735) );
  XNOR2_X1 U821 ( .A(n735), .B(KEYINPUT104), .ZN(n737) );
  NOR2_X1 U822 ( .A1(n710), .A2(G2090), .ZN(n736) );
  NOR2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U824 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n742) );
  AND2_X1 U826 ( .A1(n749), .A2(n742), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n748), .A2(n741), .ZN(n745) );
  INV_X1 U828 ( .A(n742), .ZN(n743) );
  OR2_X1 U829 ( .A1(n743), .A2(G286), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U831 ( .A(n746), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U832 ( .A1(G8), .A2(n747), .ZN(n753) );
  AND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U834 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U835 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n755), .A2(n754), .ZN(n769) );
  NOR2_X1 U837 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U838 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U839 ( .A1(n769), .A2(n757), .ZN(n758) );
  AND2_X1 U840 ( .A1(n758), .A2(n771), .ZN(n764) );
  NOR2_X1 U841 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U842 ( .A(n759), .B(KEYINPUT98), .Z(n760) );
  XNOR2_X1 U843 ( .A(KEYINPUT24), .B(n760), .ZN(n761) );
  NOR2_X1 U844 ( .A1(n771), .A2(n761), .ZN(n762) );
  XOR2_X1 U845 ( .A(KEYINPUT99), .B(n762), .Z(n763) );
  NOR2_X1 U846 ( .A1(n764), .A2(n763), .ZN(n779) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NOR2_X1 U849 ( .A1(n765), .A2(n932), .ZN(n767) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n766) );
  AND2_X1 U851 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n769), .A2(n768), .ZN(n776) );
  NAND2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n929) );
  INV_X1 U854 ( .A(n929), .ZN(n770) );
  NOR2_X1 U855 ( .A1(KEYINPUT33), .A2(n522), .ZN(n774) );
  NAND2_X1 U856 ( .A1(n932), .A2(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n775) );
  AND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U860 ( .A(G1981), .B(G305), .Z(n941) );
  NAND2_X1 U861 ( .A1(n777), .A2(n941), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n781) );
  INV_X1 U863 ( .A(KEYINPUT105), .ZN(n780) );
  XNOR2_X1 U864 ( .A(n781), .B(n780), .ZN(n813) );
  NAND2_X1 U865 ( .A1(G104), .A2(n883), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G140), .A2(n884), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U868 ( .A(KEYINPUT34), .B(n784), .ZN(n789) );
  NAND2_X1 U869 ( .A1(G116), .A2(n889), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G128), .A2(n887), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U872 ( .A(n787), .B(KEYINPUT35), .Z(n788) );
  NOR2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U874 ( .A(KEYINPUT36), .B(n790), .Z(n791) );
  XNOR2_X1 U875 ( .A(KEYINPUT93), .B(n791), .ZN(n864) );
  XNOR2_X1 U876 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NOR2_X1 U877 ( .A1(n864), .A2(n816), .ZN(n792) );
  XNOR2_X1 U878 ( .A(KEYINPUT94), .B(n792), .ZN(n1020) );
  NOR2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n825) );
  NAND2_X1 U880 ( .A1(n1020), .A2(n825), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT95), .B(n795), .Z(n822) );
  INV_X1 U882 ( .A(n822), .ZN(n812) );
  NAND2_X1 U883 ( .A1(G105), .A2(n883), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n796), .B(KEYINPUT38), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G141), .A2(n884), .ZN(n797) );
  XOR2_X1 U886 ( .A(KEYINPUT97), .B(n797), .Z(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n803) );
  NAND2_X1 U888 ( .A1(G117), .A2(n889), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G129), .A2(n887), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n865) );
  NOR2_X1 U892 ( .A1(n865), .A2(n983), .ZN(n1003) );
  NAND2_X1 U893 ( .A1(G107), .A2(n889), .ZN(n804) );
  XNOR2_X1 U894 ( .A(n804), .B(KEYINPUT96), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n883), .A2(G95), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n810) );
  NAND2_X1 U897 ( .A1(G131), .A2(n884), .ZN(n808) );
  NAND2_X1 U898 ( .A1(G119), .A2(n887), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n878) );
  INV_X1 U901 ( .A(G1991), .ZN(n982) );
  NOR2_X1 U902 ( .A1(n878), .A2(n982), .ZN(n1001) );
  OR2_X1 U903 ( .A1(n1003), .A2(n1001), .ZN(n811) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n925) );
  NAND2_X1 U905 ( .A1(n925), .A2(n825), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n828) );
  NAND2_X1 U907 ( .A1(n864), .A2(n816), .ZN(n1008) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n817) );
  AND2_X1 U909 ( .A1(n982), .A2(n878), .ZN(n1002) );
  NOR2_X1 U910 ( .A1(n817), .A2(n1002), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n523), .A2(n818), .ZN(n820) );
  AND2_X1 U912 ( .A1(n865), .A2(n983), .ZN(n819) );
  XNOR2_X1 U913 ( .A(n819), .B(KEYINPUT106), .ZN(n1011) );
  NOR2_X1 U914 ( .A1(n820), .A2(n1011), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n1008), .A2(n824), .ZN(n826) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U920 ( .A(KEYINPUT40), .B(n829), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U923 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n832) );
  XOR2_X1 U925 ( .A(KEYINPUT109), .B(n832), .Z(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G82), .ZN(G220) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n837), .ZN(G319) );
  XOR2_X1 U936 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U937 ( .A(G2090), .B(G2678), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n840), .B(KEYINPUT42), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U942 ( .A(KEYINPUT110), .B(G2100), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1956), .B(G1971), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1976), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(G1961), .B(G1966), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1981), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U953 ( .A(G2474), .B(KEYINPUT41), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(n855), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n856), .B(n982), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G100), .A2(n883), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G112), .A2(n889), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n887), .A2(G124), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n884), .A2(G136), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U965 ( .A(G160), .B(n864), .ZN(n866) );
  XOR2_X1 U966 ( .A(n866), .B(n865), .Z(n875) );
  NAND2_X1 U967 ( .A1(G118), .A2(n889), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G130), .A2(n887), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G106), .A2(n883), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G142), .A2(n884), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n871), .Z(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U976 ( .A(G162), .B(n1000), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n882) );
  XOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n880) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT114), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(n882), .B(n881), .Z(n897) );
  NAND2_X1 U982 ( .A1(G103), .A2(n883), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U985 ( .A1(G127), .A2(n887), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n888), .B(KEYINPUT112), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G115), .A2(n889), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U991 ( .A(KEYINPUT113), .B(n895), .Z(n1015) );
  XNOR2_X1 U992 ( .A(G164), .B(n1015), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n923), .B(KEYINPUT115), .ZN(n900) );
  XNOR2_X1 U996 ( .A(G171), .B(n922), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n901), .B(G286), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n904), .ZN(G397) );
  XNOR2_X1 U1001 ( .A(G2454), .B(G2446), .ZN(n914) );
  XOR2_X1 U1002 ( .A(G2430), .B(KEYINPUT108), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G2451), .B(G2443), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1005 ( .A(G2427), .B(KEYINPUT107), .Z(n908) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G2435), .B(G2438), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(n915), .A2(G14), .ZN(n921) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  INV_X1 U1021 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1022 ( .A(n922), .B(G1348), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(G1341), .B(n923), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n940) );
  XNOR2_X1 U1026 ( .A(G299), .B(G1956), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(G1971), .B(G166), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(KEYINPUT120), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT121), .B(n933), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(KEYINPUT122), .B(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(G171), .B(G1961), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(G1966), .B(G168), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n943), .B(KEYINPUT57), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n948) );
  XOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .Z(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT119), .B(n946), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n1031) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G19), .B(G1341), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT124), .B(n951), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n952), .B(G20), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT59), .B(G1348), .Z(n955) );
  XNOR2_X1 U1051 ( .A(G4), .B(n955), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT60), .B(n958), .ZN(n972) );
  XOR2_X1 U1054 ( .A(G1966), .B(G21), .Z(n967) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n961) );
  XOR2_X1 U1056 ( .A(G23), .B(KEYINPUT126), .Z(n959) );
  XNOR2_X1 U1057 ( .A(n959), .B(G1976), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1059 ( .A(KEYINPUT125), .B(G1971), .Z(n962) );
  XNOR2_X1 U1060 ( .A(G22), .B(n962), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n970) );
  XOR2_X1 U1064 ( .A(KEYINPUT123), .B(G1961), .Z(n968) );
  XNOR2_X1 U1065 ( .A(G5), .B(n968), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n973), .B(KEYINPUT61), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(KEYINPUT127), .B(n974), .ZN(n976) );
  INV_X1 U1070 ( .A(G16), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n977), .A2(G11), .ZN(n1029) );
  XOR2_X1 U1073 ( .A(G2072), .B(G33), .Z(n978) );
  NAND2_X1 U1074 ( .A1(n978), .A2(G28), .ZN(n981) );
  XOR2_X1 U1075 ( .A(G26), .B(G2067), .Z(n979) );
  XNOR2_X1 U1076 ( .A(KEYINPUT117), .B(n979), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n982), .B(G25), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n983), .B(G32), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1081 ( .A(G27), .B(n986), .Z(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n991), .B(KEYINPUT53), .ZN(n994) );
  XOR2_X1 U1085 ( .A(G2084), .B(G34), .Z(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT54), .B(n992), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G35), .B(G2090), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(KEYINPUT118), .B(n997), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(G29), .A2(n998), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(n999), .B(KEYINPUT55), .ZN(n1027) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(G160), .B(G2084), .Z(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT51), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1023) );
  XNOR2_X1 U1103 ( .A(G2072), .B(n1015), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G164), .B(G2078), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT116), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1019), .B(KEYINPUT50), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT52), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

