

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U325 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n415) );
  XNOR2_X1 U326 ( .A(n304), .B(n303), .ZN(n308) );
  XNOR2_X1 U327 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U328 ( .A(n457), .B(G176GAT), .ZN(n458) );
  XNOR2_X1 U329 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XNOR2_X1 U330 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n292) );
  XNOR2_X1 U331 ( .A(n292), .B(KEYINPUT73), .ZN(n333) );
  XOR2_X1 U332 ( .A(G176GAT), .B(G64GAT), .Z(n407) );
  XNOR2_X1 U333 ( .A(n333), .B(n407), .ZN(n294) );
  AND2_X1 U334 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n304) );
  INV_X1 U336 ( .A(G92GAT), .ZN(n295) );
  NAND2_X1 U337 ( .A1(n295), .A2(G85GAT), .ZN(n298) );
  INV_X1 U338 ( .A(G85GAT), .ZN(n296) );
  NAND2_X1 U339 ( .A1(n296), .A2(G92GAT), .ZN(n297) );
  NAND2_X1 U340 ( .A1(n298), .A2(n297), .ZN(n300) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n354) );
  XNOR2_X1 U343 ( .A(n354), .B(KEYINPUT33), .ZN(n302) );
  INV_X1 U344 ( .A(KEYINPUT75), .ZN(n301) );
  XOR2_X1 U345 ( .A(G204GAT), .B(KEYINPUT74), .Z(n306) );
  XNOR2_X1 U346 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n305) );
  XOR2_X1 U347 ( .A(n306), .B(n305), .Z(n307) );
  XNOR2_X1 U348 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G57GAT), .Z(n311) );
  XOR2_X1 U350 ( .A(G78GAT), .B(G148GAT), .Z(n420) );
  XNOR2_X1 U351 ( .A(n311), .B(n420), .ZN(n309) );
  XNOR2_X1 U352 ( .A(n310), .B(n309), .ZN(n581) );
  XNOR2_X1 U353 ( .A(n581), .B(KEYINPUT41), .ZN(n554) );
  XOR2_X1 U354 ( .A(G162GAT), .B(G85GAT), .Z(n313) );
  XOR2_X1 U355 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n439) );
  XNOR2_X1 U356 ( .A(n439), .B(n311), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n318) );
  XOR2_X1 U358 ( .A(G1GAT), .B(G113GAT), .Z(n379) );
  XNOR2_X1 U359 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n314), .B(KEYINPUT2), .ZN(n425) );
  XOR2_X1 U361 ( .A(n379), .B(n425), .Z(n316) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(n318), .B(n317), .Z(n320) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(G134GAT), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U367 ( .A(KEYINPUT94), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(G127GAT), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U370 ( .A(n324), .B(n323), .Z(n332) );
  XOR2_X1 U371 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n326) );
  XNOR2_X1 U372 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U374 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n328) );
  XNOR2_X1 U375 ( .A(KEYINPUT93), .B(KEYINPUT4), .ZN(n327) );
  XNOR2_X1 U376 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U378 ( .A(n332), .B(n331), .ZN(n520) );
  XOR2_X1 U379 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XOR2_X1 U380 ( .A(n333), .B(n440), .Z(n335) );
  NAND2_X1 U381 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U382 ( .A(n335), .B(n334), .ZN(n351) );
  XOR2_X1 U383 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n337) );
  XNOR2_X1 U384 ( .A(KEYINPUT79), .B(KEYINPUT82), .ZN(n336) );
  XNOR2_X1 U385 ( .A(n337), .B(n336), .ZN(n349) );
  XOR2_X1 U386 ( .A(G211GAT), .B(G78GAT), .Z(n339) );
  XNOR2_X1 U387 ( .A(G8GAT), .B(G22GAT), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n339), .B(n338), .ZN(n347) );
  XOR2_X1 U389 ( .A(G155GAT), .B(G57GAT), .Z(n341) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U392 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n343) );
  XNOR2_X1 U393 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U395 ( .A(n345), .B(n344), .Z(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U397 ( .A(n349), .B(n348), .Z(n350) );
  XNOR2_X1 U398 ( .A(n351), .B(n350), .ZN(n585) );
  XOR2_X1 U399 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n353) );
  XNOR2_X1 U400 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n352) );
  XNOR2_X1 U401 ( .A(n353), .B(n352), .ZN(n361) );
  XOR2_X1 U402 ( .A(G190GAT), .B(G134GAT), .Z(n443) );
  XOR2_X1 U403 ( .A(n354), .B(n443), .Z(n356) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U405 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U406 ( .A(G218GAT), .B(G162GAT), .Z(n424) );
  XOR2_X1 U407 ( .A(n357), .B(n424), .Z(n359) );
  XNOR2_X1 U408 ( .A(KEYINPUT77), .B(KEYINPUT10), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n361), .B(n360), .ZN(n369) );
  XOR2_X1 U411 ( .A(G29GAT), .B(G36GAT), .Z(n363) );
  XNOR2_X1 U412 ( .A(G50GAT), .B(G43GAT), .ZN(n362) );
  XNOR2_X1 U413 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U414 ( .A(KEYINPUT7), .B(KEYINPUT70), .Z(n365) );
  XNOR2_X1 U415 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U417 ( .A(n367), .B(n366), .Z(n376) );
  INV_X1 U418 ( .A(n376), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n369), .B(n368), .ZN(n559) );
  XNOR2_X1 U420 ( .A(KEYINPUT78), .B(n559), .ZN(n569) );
  XNOR2_X1 U421 ( .A(KEYINPUT36), .B(n569), .ZN(n588) );
  NAND2_X1 U422 ( .A1(n585), .A2(n588), .ZN(n371) );
  XOR2_X1 U423 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n372) );
  NOR2_X1 U425 ( .A1(n372), .A2(n581), .ZN(n388) );
  XOR2_X1 U426 ( .A(KEYINPUT66), .B(KEYINPUT71), .Z(n374) );
  XNOR2_X1 U427 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n387) );
  XOR2_X1 U430 ( .A(G197GAT), .B(G15GAT), .Z(n378) );
  XOR2_X1 U431 ( .A(G169GAT), .B(G8GAT), .Z(n408) );
  XOR2_X1 U432 ( .A(G22GAT), .B(G141GAT), .Z(n421) );
  XNOR2_X1 U433 ( .A(n408), .B(n421), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n380) );
  XOR2_X1 U435 ( .A(n380), .B(n379), .Z(n385) );
  XOR2_X1 U436 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n382) );
  NAND2_X1 U437 ( .A1(G229GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U439 ( .A(KEYINPUT67), .B(n383), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n577) );
  XNOR2_X1 U442 ( .A(n577), .B(KEYINPUT72), .ZN(n563) );
  NAND2_X1 U443 ( .A1(n388), .A2(n563), .ZN(n396) );
  NOR2_X1 U444 ( .A1(n577), .A2(n554), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n389), .B(KEYINPUT46), .ZN(n390) );
  NOR2_X1 U446 ( .A1(n390), .A2(n585), .ZN(n392) );
  INV_X1 U447 ( .A(KEYINPUT114), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  NOR2_X1 U449 ( .A1(n393), .A2(n559), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n394), .B(KEYINPUT47), .ZN(n395) );
  NAND2_X1 U451 ( .A1(n396), .A2(n395), .ZN(n398) );
  XNOR2_X1 U452 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n548) );
  XOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n400) );
  XNOR2_X1 U455 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n447) );
  XOR2_X1 U457 ( .A(KEYINPUT96), .B(n447), .Z(n402) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U460 ( .A(G218GAT), .B(G92GAT), .Z(n404) );
  XNOR2_X1 U461 ( .A(G36GAT), .B(G190GAT), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U463 ( .A(n406), .B(n405), .Z(n410) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U466 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n412) );
  XNOR2_X1 U467 ( .A(G197GAT), .B(G211GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U469 ( .A(G204GAT), .B(n413), .ZN(n435) );
  XNOR2_X1 U470 ( .A(n414), .B(n435), .ZN(n522) );
  NAND2_X1 U471 ( .A1(n548), .A2(n522), .ZN(n416) );
  NOR2_X1 U472 ( .A1(n520), .A2(n417), .ZN(n576) );
  XOR2_X1 U473 ( .A(KEYINPUT88), .B(KEYINPUT23), .Z(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT90), .B(KEYINPUT22), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n433) );
  XOR2_X1 U476 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n429) );
  XOR2_X1 U479 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U482 ( .A(n429), .B(n428), .Z(n431) );
  XNOR2_X1 U483 ( .A(G50GAT), .B(G106GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U485 ( .A(n433), .B(n432), .Z(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n465) );
  NAND2_X1 U487 ( .A1(n576), .A2(n465), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n436), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U489 ( .A(G176GAT), .B(G71GAT), .Z(n438) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(G113GAT), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n455) );
  XOR2_X1 U492 ( .A(G99GAT), .B(n439), .Z(n442) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U495 ( .A(n444), .B(n443), .Z(n453) );
  XOR2_X1 U496 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n446) );
  XNOR2_X1 U497 ( .A(G120GAT), .B(KEYINPUT86), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n451) );
  XOR2_X1 U499 ( .A(n447), .B(KEYINPUT85), .Z(n449) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(n526) );
  NAND2_X1 U505 ( .A1(n456), .A2(n526), .ZN(n568) );
  NOR2_X1 U506 ( .A1(n554), .A2(n568), .ZN(n459) );
  XNOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n457) );
  XOR2_X1 U508 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n461) );
  XNOR2_X1 U509 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n460) );
  XNOR2_X1 U510 ( .A(n461), .B(n460), .ZN(n477) );
  INV_X1 U511 ( .A(n520), .ZN(n506) );
  NOR2_X1 U512 ( .A1(n581), .A2(n563), .ZN(n491) );
  XOR2_X1 U513 ( .A(n522), .B(KEYINPUT27), .Z(n467) );
  NOR2_X1 U514 ( .A1(n467), .A2(n506), .ZN(n547) );
  XNOR2_X1 U515 ( .A(n465), .B(KEYINPUT28), .ZN(n528) );
  NAND2_X1 U516 ( .A1(n547), .A2(n528), .ZN(n533) );
  XOR2_X1 U517 ( .A(KEYINPUT97), .B(n533), .Z(n462) );
  NOR2_X1 U518 ( .A1(n526), .A2(n462), .ZN(n473) );
  NAND2_X1 U519 ( .A1(n522), .A2(n526), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n465), .A2(n463), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT25), .ZN(n470) );
  NOR2_X1 U522 ( .A1(n526), .A2(n465), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT26), .ZN(n575) );
  INV_X1 U524 ( .A(n575), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n470), .A2(n469), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n520), .A2(n471), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n488) );
  INV_X1 U529 ( .A(n585), .ZN(n566) );
  NOR2_X1 U530 ( .A1(n569), .A2(n566), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n474), .Z(n475) );
  NOR2_X1 U532 ( .A1(n488), .A2(n475), .ZN(n505) );
  NAND2_X1 U533 ( .A1(n491), .A2(n505), .ZN(n484) );
  NOR2_X1 U534 ( .A1(n506), .A2(n484), .ZN(n476) );
  XOR2_X1 U535 ( .A(n477), .B(n476), .Z(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT98), .B(n478), .ZN(G1324GAT) );
  INV_X1 U537 ( .A(n522), .ZN(n509) );
  NOR2_X1 U538 ( .A1(n509), .A2(n484), .ZN(n479) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  INV_X1 U540 ( .A(n526), .ZN(n534) );
  NOR2_X1 U541 ( .A1(n484), .A2(n534), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n481) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n528), .A2(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1327GAT) );
  NAND2_X1 U549 ( .A1(n588), .A2(n566), .ZN(n487) );
  NOR2_X1 U550 ( .A1(n488), .A2(n487), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT104), .B(KEYINPUT37), .Z(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n517) );
  NAND2_X1 U553 ( .A1(n517), .A2(n491), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(KEYINPUT38), .ZN(n501) );
  NOR2_X1 U555 ( .A1(n506), .A2(n501), .ZN(n496) );
  XOR2_X1 U556 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n494) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n501), .A2(n509), .ZN(n497) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n497), .Z(G1329GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n499) );
  NOR2_X1 U563 ( .A1(n534), .A2(n501), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n501), .A2(n528), .ZN(n502) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  INV_X1 U568 ( .A(n577), .ZN(n503) );
  NOR2_X1 U569 ( .A1(n554), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT108), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n505), .A2(n518), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n506), .A2(n514), .ZN(n507) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n507), .Z(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n514), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n534), .A2(n514), .ZN(n512) );
  XOR2_X1 U579 ( .A(KEYINPUT110), .B(n512), .Z(n513) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n528), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(KEYINPUT111), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n520), .A2(n530), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n524) );
  NAND2_X1 U589 ( .A1(n530), .A2(n522), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n525), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n530), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  INV_X1 U594 ( .A(n528), .ZN(n529) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n535), .A2(n548), .ZN(n543) );
  NOR2_X1 U600 ( .A1(n563), .A2(n543), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  NOR2_X1 U603 ( .A1(n554), .A2(n543), .ZN(n539) );
  XNOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n566), .A2(n543), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n541), .Z(n542) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  INV_X1 U611 ( .A(n543), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n544), .A2(n569), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  AND2_X1 U614 ( .A1(n547), .A2(n575), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n577), .A2(n558), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n553) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n554), .A2(n558), .ZN(n555) );
  XOR2_X1 U623 ( .A(n556), .B(n555), .Z(G1345GAT) );
  NOR2_X1 U624 ( .A1(n566), .A2(n558), .ZN(n557) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  XOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT121), .Z(n562) );
  INV_X1 U627 ( .A(n558), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n568), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n568), .ZN(n567) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  INV_X1 U635 ( .A(n568), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n574) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n580) );
  NOR2_X1 U643 ( .A1(n577), .A2(n580), .ZN(n578) );
  XOR2_X1 U644 ( .A(n579), .B(n578), .Z(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U646 ( .A(n580), .ZN(n589) );
  NAND2_X1 U647 ( .A1(n589), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NAND2_X1 U650 ( .A1(n589), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT126), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

