//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999, new_n1000;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  AND3_X1   g006(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n217), .A2(KEYINPUT67), .A3(new_n205), .A4(new_n207), .ZN(new_n218));
  NAND3_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g020(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n221), .A2(new_n222), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n218), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n203), .A3(new_n204), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT69), .B1(G169gat), .B2(G176gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n206), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT68), .B1(new_n215), .B2(new_n216), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n233), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n207), .A2(KEYINPUT25), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n225), .A2(new_n228), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n219), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n232), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n227), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(KEYINPUT70), .B2(KEYINPUT28), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT27), .B(G183gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n227), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(new_n251), .A3(new_n223), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(KEYINPUT71), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n256), .A2(new_n257), .B1(new_n215), .B2(new_n216), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n235), .A2(new_n236), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n258), .A2(new_n259), .B1(new_n260), .B2(KEYINPUT26), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n259), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n202), .B1(new_n244), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n230), .A2(new_n231), .B1(new_n239), .B2(new_n242), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT26), .B1(new_n235), .B2(new_n236), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n256), .A2(new_n257), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n217), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n271), .B2(KEYINPUT72), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n252), .B1(new_n272), .B2(new_n262), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n267), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n265), .B1(new_n202), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G211gat), .B(G218gat), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT77), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n278), .ZN(new_n282));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT22), .ZN(new_n284));
  INV_X1    g083(.A(G211gat), .ZN(new_n285));
  INV_X1    g084(.A(G218gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n281), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n288), .A4(new_n278), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT79), .B1(new_n275), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT37), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT79), .ZN(new_n296));
  INV_X1    g095(.A(new_n202), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n244), .A2(new_n264), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(new_n267), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n296), .B(new_n292), .C1(new_n299), .C2(new_n265), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n268), .B2(new_n273), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n202), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n297), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n293), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n294), .A2(new_n295), .A3(new_n300), .A4(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G64gat), .B(G92gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT80), .ZN(new_n308));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n292), .B1(new_n299), .B2(new_n265), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n265), .B1(new_n202), .B2(new_n302), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n313), .A2(KEYINPUT79), .B1(new_n293), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n295), .B1(new_n315), .B2(new_n300), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT38), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n310), .B(KEYINPUT81), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT38), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n275), .A2(new_n292), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(new_n295), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n292), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n306), .ZN(new_n324));
  OR2_X1    g123(.A1(G127gat), .A2(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(G113gat), .B2(G120gat), .ZN(new_n328));
  AND2_X1   g127(.A1(G113gat), .A2(G120gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n325), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT1), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n337), .A2(new_n338), .A3(new_n332), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n330), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT83), .ZN(new_n341));
  OR2_X1    g140(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(G113gat), .A3(new_n336), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(new_n334), .A3(new_n331), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n330), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347));
  AND2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351));
  INV_X1    g150(.A(G141gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(G148gat), .ZN(new_n353));
  INV_X1    g152(.A(G148gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(G141gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n351), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT82), .B1(new_n352), .B2(G148gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(new_n354), .A3(G141gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n352), .A2(G148gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  INV_X1    g161(.A(G155gat), .ZN(new_n363));
  INV_X1    g162(.A(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n365), .B2(KEYINPUT2), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n350), .A2(new_n356), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n341), .A2(new_n346), .B1(new_n347), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT86), .B(KEYINPUT5), .Z(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n366), .ZN(new_n377));
  XNOR2_X1  g176(.A(G141gat), .B(G148gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n350), .B1(new_n378), .B2(KEYINPUT2), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n377), .A2(new_n344), .A3(new_n379), .A4(new_n330), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n328), .B1(new_n325), .B2(new_n326), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n334), .B1(new_n332), .B2(new_n333), .ZN(new_n384));
  INV_X1    g183(.A(new_n331), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n343), .A2(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n367), .A3(KEYINPUT85), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n376), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT87), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  INV_X1    g190(.A(new_n389), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n386), .A2(new_n367), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n371), .B(new_n375), .C1(new_n388), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n382), .A2(new_n387), .A3(new_n376), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n389), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n374), .B1(new_n368), .B2(new_n370), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n341), .A2(new_n346), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n369), .A2(new_n401), .B1(new_n382), .B2(new_n387), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n372), .B1(new_n402), .B2(new_n373), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n395), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405));
  INV_X1    g204(.A(G85gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT0), .B(G57gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  INV_X1    g210(.A(new_n409), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n412), .B(new_n395), .C1(new_n400), .C2(new_n403), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n294), .A2(new_n300), .A3(new_n305), .A4(new_n310), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n317), .A2(new_n324), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n290), .A2(new_n301), .A3(new_n291), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n347), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n369), .ZN(new_n421));
  INV_X1    g220(.A(G228gat), .ZN(new_n422));
  INV_X1    g221(.A(G233gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n367), .A2(new_n347), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n267), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n292), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n290), .A2(new_n267), .A3(new_n291), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n367), .B1(new_n429), .B2(new_n347), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n292), .A2(new_n426), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n430), .A2(new_n431), .B1(new_n422), .B2(new_n423), .ZN(new_n432));
  NAND2_X1  g231(.A1(KEYINPUT89), .A2(G22gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT31), .B(G50gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(G106gat), .ZN(new_n435));
  XOR2_X1   g234(.A(KEYINPUT88), .B(G78gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  MUX2_X1   g236(.A(new_n433), .B(G22gat), .S(new_n437), .Z(new_n438));
  AND3_X1   g237(.A1(new_n428), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n428), .B2(new_n432), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n371), .B1(new_n388), .B2(new_n394), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT90), .B(KEYINPUT39), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n374), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n412), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n442), .A2(new_n374), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n402), .A2(new_n373), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT39), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n444), .B2(new_n412), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT40), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n444), .A2(new_n412), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT91), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n457), .B(new_n446), .C1(new_n448), .C2(new_n450), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(KEYINPUT92), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n460), .A3(new_n410), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT30), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n315), .A2(new_n462), .A3(new_n300), .A4(new_n310), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n416), .A2(KEYINPUT30), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n318), .B1(new_n315), .B2(new_n300), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n418), .B(new_n441), .C1(new_n461), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n414), .A2(new_n415), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n441), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT74), .B(G71gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G99gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G43gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n386), .B1(new_n268), .B2(new_n273), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n244), .A2(new_n264), .A3(new_n340), .ZN(new_n476));
  NAND2_X1  g275(.A1(G227gat), .A2(G233gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n476), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n477), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(new_n477), .C1(new_n480), .C2(new_n474), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n479), .A2(KEYINPUT32), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n477), .B2(KEYINPUT75), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n489), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n479), .A2(KEYINPUT32), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n484), .A2(new_n490), .A3(new_n492), .A4(new_n485), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT36), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n486), .A2(new_n493), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n484), .A2(new_n485), .B1(new_n490), .B2(new_n492), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n469), .A2(new_n470), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n498), .A2(new_n499), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n441), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT35), .B1(new_n469), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n318), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n274), .A2(new_n202), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n293), .B1(new_n507), .B2(new_n304), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n305), .B1(new_n508), .B2(new_n296), .ZN(new_n509));
  INV_X1    g308(.A(new_n300), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(KEYINPUT30), .A3(new_n416), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n512), .A2(new_n463), .B1(new_n415), .B2(new_n414), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n441), .A2(new_n494), .A3(new_n495), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G1gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT16), .ZN(new_n520));
  INV_X1    g319(.A(G15gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(G22gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G15gat), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(G1gat), .B1(new_n522), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g325(.A(G8gat), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n528), .B(new_n529), .C1(G1gat), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  OR2_X1    g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G57gat), .ZN(new_n537));
  INV_X1    g336(.A(G64gat), .ZN(new_n538));
  OR3_X1    g337(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT97), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n537), .B2(KEYINPUT97), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n537), .A2(new_n538), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n533), .B(new_n534), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n532), .B1(KEYINPUT21), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT100), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n545), .A2(KEYINPUT21), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  XOR2_X1   g350(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n552));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G127gat), .B(G155gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n549), .B(new_n550), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n558), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n563), .B1(new_n406), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT7), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n406), .B2(new_n564), .ZN(new_n567));
  NAND3_X1  g366(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G99gat), .B(G106gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G43gat), .B(G50gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n576));
  INV_X1    g375(.A(G29gat), .ZN(new_n577));
  INV_X1    g376(.A(G36gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT93), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G29gat), .A2(G36gat), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n581), .ZN(new_n587));
  NOR3_X1   g386(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G50gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT94), .B1(new_n590), .B2(G43gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT15), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(G43gat), .ZN(new_n594));
  INV_X1    g393(.A(G43gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(G50gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n574), .A2(new_n592), .A3(new_n591), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n589), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n586), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n573), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT41), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n606), .B2(new_n602), .ZN(new_n609));
  XOR2_X1   g408(.A(G134gat), .B(G162gat), .Z(new_n610));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n609), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n541), .A2(new_n544), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n571), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n569), .A2(new_n570), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n569), .A2(new_n570), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n545), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT101), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n615), .A2(new_n624), .A3(new_n618), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n545), .A2(new_n616), .A3(KEYINPUT10), .A4(new_n617), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n622), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT102), .B(G176gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n623), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n622), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n560), .A2(new_n562), .A3(new_n613), .A4(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n572), .B1(new_n586), .B2(new_n600), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n583), .A2(new_n581), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n588), .A2(new_n582), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n585), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n575), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n579), .A2(new_n581), .B1(G29gat), .B2(G36gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n593), .A2(new_n597), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n650), .A3(KEYINPUT17), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n527), .A2(new_n531), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n641), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n532), .B1(new_n586), .B2(new_n600), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n653), .A2(KEYINPUT18), .A3(new_n654), .A4(new_n655), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n532), .A2(new_n586), .A3(new_n600), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n646), .A2(new_n650), .B1(new_n527), .B2(new_n531), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n654), .B(KEYINPUT13), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT95), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n652), .A2(new_n650), .A3(new_n646), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n655), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n667));
  INV_X1    g466(.A(new_n663), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n658), .A2(new_n659), .A3(new_n664), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671));
  INV_X1    g470(.A(G197gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT11), .B(G169gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT12), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT96), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT95), .B(new_n663), .C1(new_n665), .C2(new_n655), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n682), .A2(new_n659), .A3(new_n658), .A4(new_n676), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n670), .A2(KEYINPUT96), .A3(new_n677), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n640), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n518), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n468), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n519), .ZN(G1324gat));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n466), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n529), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT103), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(G1325gat));
  INV_X1    g496(.A(new_n688), .ZN(new_n698));
  AOI21_X1  g497(.A(G15gat), .B1(new_n698), .B2(new_n503), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n500), .A2(new_n496), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n521), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT104), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n698), .B2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n441), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  AOI22_X1  g505(.A1(new_n467), .A2(new_n501), .B1(new_n505), .B2(new_n516), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n613), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n561), .B(new_n559), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n638), .A3(new_n686), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n468), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n577), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT44), .B1(new_n707), .B2(new_n613), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  INV_X1    g515(.A(new_n613), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n700), .B1(new_n513), .B2(new_n441), .ZN(new_n718));
  INV_X1    g517(.A(new_n466), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n719), .A2(new_n410), .A3(new_n460), .A4(new_n455), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n306), .B2(new_n323), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n470), .B1(new_n722), .B2(new_n317), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n718), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  AND4_X1   g523(.A1(new_n514), .A2(new_n515), .A3(new_n466), .A4(new_n468), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n716), .B(new_n717), .C1(new_n724), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n715), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n709), .A2(new_n638), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n686), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n685), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n729), .A2(KEYINPUT106), .A3(new_n737), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n468), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n714), .B1(new_n741), .B2(new_n577), .ZN(G1328gat));
  NAND2_X1  g541(.A1(new_n719), .A2(new_n578), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n708), .A2(new_n710), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT46), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n740), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT108), .B1(new_n751), .B2(new_n719), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n753), .B(new_n736), .C1(new_n715), .C2(new_n728), .ZN(new_n754));
  OAI211_X1 g553(.A(KEYINPUT108), .B(new_n719), .C1(new_n738), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G36gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n752), .B2(new_n756), .ZN(G1329gat));
  NAND2_X1  g556(.A1(new_n729), .A2(new_n737), .ZN(new_n758));
  OAI21_X1  g557(.A(G43gat), .B1(new_n758), .B2(new_n700), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n711), .A2(new_n595), .A3(new_n503), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(KEYINPUT47), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n760), .ZN(new_n762));
  INV_X1    g561(.A(new_n700), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n738), .B2(new_n754), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(G43gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n765), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g565(.A(G50gat), .B1(new_n758), .B2(new_n441), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n711), .A2(new_n590), .A3(new_n470), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(KEYINPUT48), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n768), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n470), .B1(new_n738), .B2(new_n754), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(G50gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n772), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g572(.A1(new_n709), .A2(new_n613), .A3(new_n638), .A4(new_n734), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT109), .Z(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n518), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n468), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n537), .ZN(G1332gat));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n466), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  AND2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n779), .B2(new_n780), .ZN(G1333gat));
  INV_X1    g582(.A(new_n776), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(G71gat), .A3(new_n763), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n776), .A2(new_n498), .A3(new_n499), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(G71gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n470), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g589(.A1(new_n735), .A2(new_n709), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n638), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n715), .B2(new_n728), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n712), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G85gat), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n793), .B2(new_n712), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n717), .B(new_n791), .C1(new_n724), .C2(new_n727), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n518), .A2(KEYINPUT51), .A3(new_n717), .A4(new_n791), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT111), .B1(new_n799), .B2(new_n800), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n712), .A2(new_n406), .A3(new_n638), .ZN(new_n806));
  OAI22_X1  g605(.A1(new_n796), .A2(new_n797), .B1(new_n805), .B2(new_n806), .ZN(G1336gat));
  AOI21_X1  g606(.A(new_n564), .B1(new_n793), .B2(new_n719), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n719), .A2(new_n564), .A3(new_n638), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n801), .B2(new_n802), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT52), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n812));
  AND2_X1   g611(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n808), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n805), .A2(new_n809), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(G1337gat));
  INV_X1    g615(.A(G99gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n503), .A2(new_n817), .A3(new_n638), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n793), .A2(new_n763), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n805), .A2(new_n818), .B1(new_n819), .B2(new_n817), .ZN(G1338gat));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  INV_X1    g620(.A(new_n792), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n716), .B1(new_n518), .B2(new_n717), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n707), .A2(KEYINPUT44), .A3(new_n613), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n470), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n793), .A2(KEYINPUT115), .A3(new_n470), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(G106gat), .A3(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n441), .A2(G106gat), .A3(new_n639), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n803), .B2(new_n804), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n825), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT113), .B1(new_n825), .B2(G106gat), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n830), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n801), .B2(new_n802), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT53), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT114), .B(new_n836), .C1(new_n801), .C2(new_n802), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n821), .A2(new_n832), .B1(new_n835), .B2(new_n841), .ZN(G1339gat));
  INV_X1    g641(.A(new_n709), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n625), .A2(new_n626), .A3(new_n621), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n628), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n632), .B1(new_n636), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n847), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n633), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n732), .A2(new_n733), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n666), .A2(new_n668), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n675), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n638), .A2(new_n683), .A3(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT116), .Z(new_n859));
  AOI21_X1  g658(.A(new_n717), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n717), .A2(new_n853), .A3(new_n683), .A4(new_n857), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n843), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n640), .A2(new_n735), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n712), .A3(new_n515), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n719), .B1(new_n867), .B2(KEYINPUT117), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n504), .B1(new_n863), .B2(new_n865), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n712), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n332), .A3(new_n735), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n719), .A2(new_n468), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n686), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1340gat));
  OAI211_X1 g676(.A(new_n872), .B(new_n638), .C1(new_n338), .C2(new_n337), .ZN(new_n878));
  OAI21_X1  g677(.A(G120gat), .B1(new_n875), .B2(new_n639), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1341gat));
  AOI21_X1  g679(.A(G127gat), .B1(new_n872), .B2(new_n709), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n709), .A2(G127gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT118), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n881), .A2(new_n884), .ZN(G1342gat));
  NAND2_X1  g684(.A1(new_n867), .A2(KEYINPUT117), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n613), .A2(G134gat), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n466), .A3(new_n871), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT119), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n868), .A2(new_n890), .A3(new_n871), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G134gat), .B1(new_n875), .B2(new_n613), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n889), .A2(KEYINPUT56), .A3(new_n891), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n866), .A2(new_n898), .A3(new_n470), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n874), .A2(new_n700), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n858), .B1(new_n686), .B2(new_n852), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n613), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n709), .B1(new_n861), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n470), .B1(new_n903), .B2(new_n864), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n900), .B1(new_n904), .B2(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G141gat), .B1(new_n906), .B2(new_n686), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n685), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT105), .B1(new_n684), .B2(new_n685), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n852), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n858), .B(KEYINPUT116), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n613), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n709), .B1(new_n912), .B2(new_n861), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n470), .B1(new_n913), .B2(new_n864), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n900), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n686), .A2(G141gat), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT58), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n899), .B2(new_n905), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n735), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n922), .A2(G141gat), .B1(new_n915), .B2(new_n916), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT58), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(G1344gat));
  NAND3_X1  g724(.A1(new_n915), .A2(new_n354), .A3(new_n638), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G148gat), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n906), .B(KEYINPUT120), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n638), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n470), .A2(new_n898), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n902), .A2(new_n861), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n843), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n709), .A2(new_n613), .A3(new_n639), .A4(new_n686), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n441), .B1(new_n863), .B2(new_n865), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n936), .B(new_n638), .C1(new_n937), .C2(new_n898), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n938), .A2(new_n900), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n927), .B1(new_n939), .B2(G148gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n926), .B1(new_n930), .B2(new_n940), .ZN(G1345gat));
  AOI21_X1  g740(.A(G155gat), .B1(new_n915), .B2(new_n709), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n843), .A2(new_n363), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n929), .B2(new_n943), .ZN(G1346gat));
  AOI21_X1  g743(.A(G162gat), .B1(new_n915), .B2(new_n717), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n613), .A2(new_n364), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n929), .B2(new_n946), .ZN(G1347gat));
  NOR2_X1   g746(.A1(new_n466), .A2(new_n712), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n869), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n686), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n735), .A2(new_n203), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(G1348gat));
  NOR2_X1   g751(.A1(new_n949), .A2(new_n639), .ZN(new_n953));
  XOR2_X1   g752(.A(KEYINPUT121), .B(G176gat), .Z(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(G1349gat));
  NOR2_X1   g754(.A1(new_n949), .A2(new_n843), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n249), .B1(KEYINPUT122), .B2(G183gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n226), .A2(KEYINPUT122), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n960), .B(new_n961), .ZN(G1350gat));
  XNOR2_X1  g761(.A(KEYINPUT61), .B(G190gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n613), .ZN(new_n965));
  MUX2_X1   g764(.A(new_n963), .B(new_n964), .S(new_n965), .Z(G1351gat));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n700), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n936), .B(new_n968), .C1(new_n937), .C2(new_n898), .ZN(new_n969));
  OAI21_X1  g768(.A(G197gat), .B1(new_n969), .B2(new_n686), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n914), .A2(new_n967), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n672), .A3(new_n735), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1352gat));
  OAI21_X1  g772(.A(KEYINPUT123), .B1(new_n938), .B2(new_n967), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n935), .B1(new_n914), .B2(KEYINPUT57), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n975), .A2(new_n976), .A3(new_n638), .A4(new_n968), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n977), .A3(G204gat), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n639), .A2(G204gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n937), .A2(new_n968), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT62), .Z(new_n981));
  NAND2_X1  g780(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n978), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1353gat));
  OAI211_X1 g785(.A(KEYINPUT63), .B(G211gat), .C1(new_n969), .C2(new_n843), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(KEYINPUT126), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(KEYINPUT126), .ZN(new_n989));
  OAI21_X1  g788(.A(G211gat), .B1(new_n969), .B2(new_n843), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT63), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n988), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n971), .A2(new_n285), .A3(new_n709), .ZN(new_n994));
  XOR2_X1   g793(.A(new_n994), .B(KEYINPUT125), .Z(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(G1354gat));
  AND2_X1   g795(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n717), .B1(new_n969), .B2(KEYINPUT127), .ZN(new_n998));
  OAI21_X1  g797(.A(G218gat), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n971), .A2(new_n286), .A3(new_n717), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1355gat));
endmodule


