//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(G237), .A2(G953), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(G143), .A3(G214), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT92), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT18), .A2(G131), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n199), .B(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n206), .A2(KEYINPUT76), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(KEYINPUT76), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(G146), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n201), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AND4_X1   g028(.A1(G143), .A2(new_n190), .A3(new_n191), .A4(G214), .ZN(new_n215));
  AOI21_X1  g029(.A(G143), .B1(new_n195), .B2(G214), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT93), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n197), .A2(KEYINPUT93), .A3(G131), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(new_n220), .C1(G131), .C2(new_n197), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT16), .ZN(new_n222));
  OR3_X1    g036(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G146), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT19), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n207), .A2(new_n225), .A3(new_n209), .ZN(new_n226));
  INV_X1    g040(.A(new_n206), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n221), .B(new_n224), .C1(new_n228), .C2(G146), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n189), .B1(new_n214), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n223), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n208), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n224), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n219), .A2(new_n220), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT94), .B1(new_n236), .B2(KEYINPUT17), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT94), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT17), .ZN(new_n239));
  AOI211_X1 g053(.A(new_n238), .B(new_n239), .C1(new_n219), .C2(new_n220), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n235), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n231), .B1(new_n241), .B2(KEYINPUT95), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT93), .B1(new_n197), .B2(G131), .ZN(new_n243));
  INV_X1    g057(.A(G131), .ZN(new_n244));
  AOI211_X1 g058(.A(new_n218), .B(new_n244), .C1(new_n194), .C2(new_n196), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT17), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n238), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n236), .A2(KEYINPUT94), .A3(KEYINPUT17), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n234), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT95), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n213), .B1(new_n242), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n230), .B1(new_n252), .B2(new_n189), .ZN(new_n253));
  NOR2_X1   g067(.A1(G475), .A2(G902), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT20), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n231), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n249), .B2(new_n250), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n241), .A2(KEYINPUT95), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n189), .B(new_n214), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n230), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT20), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n254), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(G234), .A2(G237), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(G952), .A3(new_n191), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT99), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT72), .B(G902), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n271), .A2(G953), .A3(new_n266), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT21), .B(G898), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT96), .ZN(new_n276));
  INV_X1    g090(.A(G122), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G116), .ZN(new_n278));
  INV_X1    g092(.A(G116), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT96), .A3(G122), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G107), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n279), .A2(G122), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n193), .A2(G128), .ZN(new_n286));
  INV_X1    g100(.A(G128), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G143), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n288), .A3(G134), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n288), .ZN(new_n290));
  INV_X1    g104(.A(G134), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT97), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n284), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT14), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n278), .B2(new_n280), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT97), .B1(new_n298), .B2(new_n283), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n296), .B(new_n299), .C1(KEYINPUT14), .C2(new_n281), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n293), .B1(new_n300), .B2(G107), .ZN(new_n301));
  INV_X1    g115(.A(new_n285), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n282), .B1(new_n281), .B2(new_n284), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT13), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n288), .A2(new_n305), .A3(G134), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n292), .A2(new_n289), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n292), .B2(new_n289), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  INV_X1    g124(.A(G217), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n310), .A2(new_n311), .A3(G953), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n301), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT98), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n313), .B1(new_n301), .B2(new_n309), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n314), .B2(new_n315), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n270), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G478), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(KEYINPUT15), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n319), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n242), .A2(new_n251), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n189), .B1(new_n325), .B2(new_n214), .ZN(new_n326));
  INV_X1    g140(.A(new_n189), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n327), .B(new_n213), .C1(new_n242), .C2(new_n251), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G475), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n265), .A2(new_n275), .A3(new_n323), .A4(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G214), .B1(G237), .B2(G902), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G210), .B1(G237), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n282), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n188), .A2(KEYINPUT80), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G104), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n282), .A3(G104), .ZN(new_n343));
  NAND2_X1  g157(.A1(KEYINPUT3), .A2(G107), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(G107), .B1(new_n338), .B2(new_n340), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT81), .B1(new_n282), .B2(G104), .ZN(new_n347));
  OAI21_X1  g161(.A(G101), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n339), .A2(G104), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n188), .A2(KEYINPUT80), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n282), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n345), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n355));
  INV_X1    g169(.A(G113), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n279), .A2(G119), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT5), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G119), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G116), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n279), .A2(G119), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT5), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n356), .A2(KEYINPUT2), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G113), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n359), .A2(new_n363), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n354), .A2(new_n355), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G122), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT8), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n352), .B(G101), .C1(new_n346), .C2(new_n347), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n345), .A3(new_n369), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT89), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n369), .B1(new_n374), .B2(new_n345), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n371), .B(new_n373), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n344), .B1(new_n337), .B2(new_n188), .ZN(new_n381));
  OAI21_X1  g195(.A(G101), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n345), .A3(KEYINPUT4), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(G101), .C1(new_n380), .C2(new_n381), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n364), .A2(new_n368), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n364), .A2(new_n368), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n375), .A3(new_n372), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT64), .B1(new_n193), .B2(G146), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n208), .A3(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n193), .A2(G146), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n193), .A2(G146), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n397));
  OAI21_X1  g211(.A(G128), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G143), .B(G146), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n287), .A2(KEYINPUT1), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n395), .A2(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n204), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n191), .A2(G224), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n405), .A2(KEYINPUT90), .ZN(new_n406));
  AND2_X1   g220(.A1(KEYINPUT0), .A2(G128), .ZN(new_n407));
  NOR2_X1   g221(.A1(KEYINPUT0), .A2(G128), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n395), .A2(new_n409), .B1(new_n399), .B2(new_n407), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n402), .B(new_n406), .C1(new_n204), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(KEYINPUT90), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n410), .A2(new_n204), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n414), .A2(KEYINPUT90), .A3(new_n402), .A4(new_n405), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n390), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n324), .B1(new_n379), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n378), .A2(new_n390), .A3(new_n413), .A4(new_n415), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT91), .A3(new_n324), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n402), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n403), .B(KEYINPUT88), .Z(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n389), .A2(new_n375), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT87), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n389), .A2(new_n429), .A3(new_n375), .ZN(new_n430));
  INV_X1    g244(.A(new_n372), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  INV_X1    g247(.A(new_n390), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n372), .B1(new_n427), .B2(KEYINPUT87), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n426), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n335), .B1(new_n422), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n437), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n436), .A2(new_n430), .B1(KEYINPUT6), .B2(new_n390), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n425), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n442), .A2(new_n334), .A3(new_n421), .A4(new_n419), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n333), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n331), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n360), .A2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n287), .A2(G119), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT73), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT24), .B(G110), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT23), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n287), .A2(KEYINPUT23), .A3(G119), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n447), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G110), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n222), .A2(G146), .A3(new_n223), .ZN(new_n460));
  AOI21_X1  g274(.A(G146), .B1(new_n222), .B2(new_n223), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n454), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n234), .A2(KEYINPUT74), .A3(new_n454), .A4(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n456), .A2(new_n447), .ZN(new_n467));
  INV_X1    g281(.A(G110), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(KEYINPUT75), .A3(new_n468), .A4(new_n457), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT75), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n458), .B2(G110), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n450), .A2(new_n452), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n469), .B(new_n471), .C1(new_n472), .C2(new_n453), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n210), .A2(new_n224), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT22), .B(G137), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n466), .A2(new_n475), .A3(new_n479), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n270), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n481), .A2(KEYINPUT25), .A3(new_n270), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n311), .B1(new_n270), .B2(G234), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT77), .ZN(new_n490));
  INV_X1    g304(.A(new_n482), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n479), .B1(new_n466), .B2(new_n475), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n488), .A2(G902), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n488), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n485), .B2(new_n486), .ZN(new_n498));
  INV_X1    g312(.A(new_n495), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT77), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n395), .A2(new_n398), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n399), .A2(new_n400), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT11), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n291), .B2(G137), .ZN(new_n506));
  INV_X1    g320(.A(G137), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT11), .A3(G134), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n291), .A2(G137), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n506), .A2(new_n508), .A3(new_n244), .A4(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n291), .A2(G137), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n507), .A2(G134), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n504), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT67), .B1(new_n401), .B2(new_n514), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n510), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n410), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT30), .A4(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT65), .B1(new_n521), .B2(new_n410), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(KEYINPUT65), .A3(new_n410), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n401), .B1(new_n527), .B2(new_n514), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n515), .A2(KEYINPUT66), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n525), .A2(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n388), .B(new_n523), .C1(new_n530), .C2(KEYINPUT30), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n518), .A2(new_n522), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n386), .A2(new_n387), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n517), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n517), .A2(new_n518), .A3(new_n534), .A4(new_n522), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT68), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n195), .A2(G210), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT27), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(G101), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n531), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n531), .A2(new_n538), .A3(KEYINPUT31), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n504), .A2(new_n515), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n534), .A3(new_n522), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n514), .A2(new_n527), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n529), .A2(new_n504), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n526), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n524), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n535), .A2(new_n537), .B1(new_n388), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n560), .B2(new_n551), .ZN(new_n561));
  INV_X1    g375(.A(new_n542), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n547), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  NOR2_X1   g379(.A1(G472), .A2(G902), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n545), .A2(new_n546), .B1(new_n561), .B2(new_n562), .ZN(new_n568));
  INV_X1    g382(.A(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT32), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n531), .A2(new_n538), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n562), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT29), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n573), .B(new_n574), .C1(new_n561), .C2(new_n562), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n532), .A2(new_n517), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n388), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n538), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT70), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n535), .A2(new_n537), .B1(new_n576), .B2(new_n388), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n551), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n553), .B2(new_n554), .ZN(new_n584));
  INV_X1    g398(.A(new_n554), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT71), .A3(new_n552), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n562), .A2(new_n574), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n579), .A2(new_n582), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n575), .A2(new_n589), .A3(new_n270), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n501), .B1(new_n571), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT86), .ZN(new_n593));
  XOR2_X1   g407(.A(G110), .B(G140), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT79), .ZN(new_n595));
  INV_X1    g409(.A(G227), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(G953), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n595), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n208), .A2(G143), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n287), .B1(new_n600), .B2(KEYINPUT1), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n503), .B1(new_n601), .B2(new_n399), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n374), .A2(new_n345), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n383), .A2(new_n385), .A3(new_n410), .ZN(new_n606));
  INV_X1    g420(.A(new_n521), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n374), .A2(new_n504), .A3(KEYINPUT10), .A4(new_n345), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT82), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT12), .B1(new_n521), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n354), .A2(new_n401), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n603), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n614), .B2(new_n521), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n607), .B(new_n611), .C1(new_n613), .C2(new_n603), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT83), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT83), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n619), .B(new_n609), .C1(new_n615), .C2(new_n616), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n599), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n609), .A2(new_n599), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n521), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(KEYINPUT84), .A3(new_n521), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n324), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n614), .A2(new_n521), .A3(new_n612), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n374), .A2(new_n345), .A3(new_n602), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n504), .B1(new_n345), .B2(new_n374), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n521), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n611), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n622), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n623), .A2(KEYINPUT84), .A3(new_n521), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT84), .B1(new_n623), .B2(new_n521), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n609), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n638), .B2(new_n598), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n271), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT85), .B(G469), .Z(new_n641));
  AOI22_X1  g455(.A1(new_n629), .A2(G469), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(G221), .B1(new_n310), .B2(G902), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT78), .Z(new_n644));
  OAI21_X1  g458(.A(new_n593), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n626), .A2(new_n627), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n599), .B1(new_n646), .B2(new_n609), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n270), .B(new_n641), .C1(new_n647), .C2(new_n635), .ZN(new_n648));
  INV_X1    g462(.A(new_n620), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n634), .A2(new_n630), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n619), .B1(new_n650), .B2(new_n609), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n598), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n628), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(G469), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n644), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(KEYINPUT86), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n446), .A2(new_n592), .A3(new_n645), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G101), .ZN(G3));
  NOR3_X1   g474(.A1(new_n642), .A2(new_n593), .A3(new_n644), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT86), .B1(new_n656), .B2(new_n657), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n271), .B1(new_n547), .B2(new_n563), .ZN(new_n664));
  INV_X1    g478(.A(G472), .ZN(new_n665));
  OAI22_X1  g479(.A1(new_n664), .A2(new_n665), .B1(new_n569), .B2(new_n568), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n501), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n263), .B1(new_n262), .B2(new_n254), .ZN(new_n668));
  AOI211_X1 g482(.A(KEYINPUT20), .B(new_n255), .C1(new_n260), .C2(new_n261), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n214), .B1(new_n258), .B2(new_n259), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n327), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n671), .B2(new_n260), .ZN(new_n672));
  INV_X1    g486(.A(G475), .ZN(new_n673));
  OAI22_X1  g487(.A1(new_n668), .A2(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n319), .A2(new_n320), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT101), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n319), .A2(new_n677), .A3(new_n320), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT33), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n316), .B2(new_n318), .ZN(new_n680));
  INV_X1    g494(.A(new_n314), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n317), .A3(KEYINPUT100), .A4(KEYINPUT33), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n317), .A2(KEYINPUT33), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n683), .B1(new_n684), .B2(new_n314), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n271), .A2(new_n320), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n680), .A2(new_n682), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n676), .A2(new_n678), .A3(new_n687), .ZN(new_n688));
  AND4_X1   g502(.A1(new_n444), .A2(new_n674), .A3(new_n275), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n663), .A2(new_n667), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT34), .B(G104), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G6));
  XNOR2_X1  g506(.A(new_n274), .B(KEYINPUT102), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n422), .A2(new_n438), .A3(new_n335), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n420), .A2(KEYINPUT91), .A3(new_n324), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT91), .B1(new_n420), .B2(new_n324), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n334), .B1(new_n697), .B2(new_n442), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n332), .B(new_n693), .C1(new_n694), .C2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n699), .A2(new_n323), .A3(new_n674), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n645), .A3(new_n658), .A4(new_n667), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT35), .B(G107), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G9));
  NOR2_X1   g517(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n476), .B(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n494), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n498), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n666), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n446), .A2(new_n645), .A3(new_n658), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT37), .B(G110), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G12));
  AOI22_X1  g525(.A1(new_n567), .A2(new_n570), .B1(G472), .B2(new_n590), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n712), .A2(new_n445), .A3(new_n707), .ZN(new_n713));
  INV_X1    g527(.A(G900), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n269), .B1(new_n272), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n674), .A2(new_n323), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n663), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT103), .B(G128), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G30));
  NOR2_X1   g533(.A1(new_n694), .A2(new_n698), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT38), .Z(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n332), .A3(new_n707), .ZN(new_n722));
  INV_X1    g536(.A(new_n674), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n323), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n715), .B(KEYINPUT39), .Z(new_n725));
  NAND2_X1  g539(.A1(new_n663), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n726), .A2(KEYINPUT40), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(KEYINPUT40), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n572), .A2(new_n542), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n729), .B(new_n324), .C1(new_n578), .C2(new_n542), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n571), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n724), .A2(new_n727), .A3(new_n728), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G143), .ZN(G45));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  INV_X1    g549(.A(new_n715), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n674), .A2(new_n688), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n674), .A2(new_n688), .A3(new_n736), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT104), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n663), .A2(new_n713), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n639), .B2(new_n271), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n648), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n742), .B1(new_n744), .B2(new_n644), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n743), .A2(new_n648), .A3(KEYINPUT105), .A4(new_n657), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n689), .A3(new_n592), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n592), .A3(new_n700), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  NOR2_X1   g567(.A1(new_n747), .A2(new_n331), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n713), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  AND3_X1   g570(.A1(new_n745), .A2(new_n693), .A3(new_n746), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n319), .B(new_n321), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n674), .A2(new_n444), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(G472), .B1(new_n568), .B2(new_n271), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n498), .A2(new_n499), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n579), .A2(new_n582), .A3(new_n587), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n762), .A2(new_n562), .B1(new_n545), .B2(new_n546), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n760), .B(new_n761), .C1(new_n569), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT106), .B(G122), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G24));
  AND3_X1   g582(.A1(new_n745), .A2(new_n444), .A3(new_n746), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n763), .A2(new_n569), .ZN(new_n770));
  INV_X1    g584(.A(new_n707), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n770), .A2(new_n760), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n772), .A3(new_n739), .A4(new_n737), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  AND2_X1   g588(.A1(new_n739), .A2(new_n737), .ZN(new_n775));
  INV_X1    g589(.A(new_n761), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n712), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n439), .A2(new_n332), .A3(new_n443), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n642), .A2(new_n778), .A3(new_n779), .A4(new_n644), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n642), .A2(new_n778), .A3(new_n644), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n739), .A2(new_n592), .A3(new_n737), .A4(new_n782), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n775), .A2(new_n781), .B1(new_n783), .B2(new_n779), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT107), .B(G131), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G33));
  NAND3_X1  g600(.A1(new_n592), .A2(new_n782), .A3(new_n716), .ZN(new_n787));
  XOR2_X1   g601(.A(KEYINPUT108), .B(G134), .Z(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G36));
  NAND2_X1  g603(.A1(new_n723), .A2(new_n688), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n666), .A2(new_n771), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT110), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT112), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n621), .A2(new_n628), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT45), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(KEYINPUT45), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(G469), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(G469), .A2(G902), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT46), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n640), .B2(new_n641), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n804), .A2(KEYINPUT46), .A3(new_n805), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n644), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n725), .ZN(new_n810));
  INV_X1    g624(.A(new_n778), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n797), .B2(new_n798), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n800), .B(new_n814), .C1(new_n813), .C2(new_n812), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  XNOR2_X1  g630(.A(new_n809), .B(KEYINPUT47), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n775), .A2(new_n712), .A3(new_n501), .A4(new_n811), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT113), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NOR2_X1   g635(.A1(G952), .A2(G953), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT121), .Z(new_n823));
  NOR4_X1   g637(.A1(new_n794), .A2(new_n268), .A3(new_n747), .A4(new_n778), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n777), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT48), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n732), .A2(new_n501), .A3(new_n268), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n748), .A3(new_n811), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n674), .A2(new_n688), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(G952), .B(new_n191), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n794), .A2(new_n268), .A3(new_n764), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(new_n769), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n748), .A2(KEYINPUT119), .A3(new_n333), .ZN(new_n835));
  INV_X1    g649(.A(new_n721), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n747), .B2(new_n332), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n828), .A2(new_n674), .A3(new_n688), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n824), .B2(new_n772), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n744), .A2(new_n657), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n811), .B(new_n832), .C1(new_n817), .C2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(KEYINPUT120), .A3(new_n845), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(KEYINPUT51), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT120), .B1(new_n843), .B2(new_n845), .ZN(new_n851));
  OAI221_X1 g665(.A(new_n834), .B1(new_n848), .B2(KEYINPUT51), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n759), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n642), .A2(new_n644), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n771), .A2(new_n715), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n732), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n740), .A2(new_n717), .A3(new_n773), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT115), .B1(new_n857), .B2(new_n858), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT52), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n857), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n659), .A2(new_n709), .A3(new_n701), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n674), .A2(new_n444), .A3(new_n688), .A4(new_n693), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT114), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n645), .A2(new_n667), .A3(new_n658), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n787), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n783), .A2(new_n779), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n777), .A2(new_n780), .A3(new_n739), .A4(new_n737), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n748), .B(new_n592), .C1(new_n689), .C2(new_n700), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n880), .A2(new_n755), .A3(new_n766), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n712), .A2(new_n707), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n674), .A2(new_n778), .A3(new_n758), .A4(new_n715), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n645), .A4(new_n658), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n772), .A2(new_n739), .A3(new_n737), .A4(new_n782), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n875), .A2(new_n879), .A3(new_n881), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT53), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n784), .A2(new_n876), .A3(new_n886), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n880), .A2(new_n755), .A3(new_n766), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n868), .A3(new_n874), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n571), .A2(new_n591), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n444), .A3(new_n771), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n645), .A2(new_n658), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n775), .B2(new_n716), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n862), .A3(new_n773), .A4(new_n856), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n857), .A2(KEYINPUT52), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n890), .A2(new_n892), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n867), .A2(new_n889), .B1(KEYINPUT53), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n754), .A2(new_n713), .B1(new_n757), .B2(new_n765), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n903), .A2(KEYINPUT118), .A3(new_n880), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT118), .B1(new_n903), .B2(new_n880), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n879), .A2(new_n887), .ZN(new_n907));
  INV_X1    g721(.A(new_n874), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n659), .A2(new_n701), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT53), .A4(new_n709), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n865), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n866), .B1(new_n864), .B2(KEYINPUT52), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n899), .A2(new_n898), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n888), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n916), .B1(new_n900), .B2(new_n917), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n914), .B(new_n915), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n902), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n823), .B1(new_n852), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n836), .A2(new_n761), .A3(new_n657), .A4(new_n332), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n744), .B(KEYINPUT49), .ZN(new_n926));
  OR4_X1    g740(.A1(new_n732), .A2(new_n925), .A3(new_n790), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(G75));
  NOR2_X1   g742(.A1(new_n440), .A2(new_n441), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n426), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n442), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n917), .B1(new_n918), .B2(new_n888), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT117), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n934), .A2(new_n919), .B1(new_n867), .B2(new_n911), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n935), .A2(new_n270), .A3(new_n334), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n932), .B1(new_n936), .B2(KEYINPUT56), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n191), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n935), .A2(new_n941), .A3(new_n270), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT122), .B1(new_n943), .B2(new_n271), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n335), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n932), .A2(KEYINPUT56), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(G51));
  NAND2_X1  g762(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n922), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n805), .B(KEYINPUT57), .Z(new_n951));
  AOI21_X1  g765(.A(new_n639), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n953));
  INV_X1    g767(.A(new_n804), .ZN(new_n954));
  AOI22_X1  g768(.A1(new_n952), .A2(new_n953), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n951), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n949), .B2(new_n922), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT123), .B1(new_n957), .B2(new_n639), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n938), .B1(new_n955), .B2(new_n958), .ZN(G54));
  OAI21_X1  g773(.A(new_n941), .B1(new_n935), .B2(new_n270), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n943), .A2(KEYINPUT122), .A3(new_n271), .ZN(new_n961));
  AND2_X1   g775(.A1(KEYINPUT58), .A2(G475), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n253), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n939), .B1(new_n963), .B2(new_n253), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n963), .B2(new_n253), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(G60));
  AND3_X1   g782(.A1(new_n680), .A2(new_n682), .A3(new_n685), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT59), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n950), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n923), .B2(new_n971), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n972), .A2(new_n938), .A3(new_n973), .ZN(G63));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n943), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n979), .B2(new_n705), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(KEYINPUT61), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n938), .B1(new_n979), .B2(new_n705), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n978), .B1(new_n491), .B2(new_n492), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n983), .B(new_n982), .C1(new_n980), .C2(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G66));
  INV_X1    g801(.A(G224), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n273), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n892), .B2(G953), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n929), .B1(G898), .B2(new_n191), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G69));
  OAI21_X1  g806(.A(new_n523), .B1(new_n530), .B2(KEYINPUT30), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(new_n228), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(G953), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n815), .A2(new_n820), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n829), .B1(new_n758), .B2(new_n723), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n592), .A2(new_n811), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n726), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n897), .A2(new_n773), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n733), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n1001), .A2(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(KEYINPUT62), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n995), .B1(new_n996), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n714), .A2(G953), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n809), .A2(new_n725), .A3(new_n853), .A4(new_n777), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1009), .A2(new_n879), .A3(new_n1000), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n815), .A2(new_n820), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1008), .B1(new_n1011), .B2(new_n191), .ZN(new_n1012));
  OAI21_X1  g826(.A(G953), .B1(new_n596), .B2(new_n714), .ZN(new_n1013));
  OR3_X1    g827(.A1(new_n1005), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1013), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(G72));
  NAND3_X1  g830(.A1(new_n996), .A2(new_n892), .A3(new_n1004), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  AOI21_X1  g833(.A(new_n729), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n531), .A2(new_n538), .A3(new_n562), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n815), .A2(new_n820), .A3(new_n1010), .A4(new_n892), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1021), .B1(new_n1022), .B2(new_n1019), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n573), .B(KEYINPUT127), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n543), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n901), .A2(new_n1019), .A3(new_n1025), .ZN(new_n1026));
  NOR4_X1   g840(.A1(new_n1020), .A2(new_n1023), .A3(new_n938), .A4(new_n1026), .ZN(G57));
endmodule


