//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT64), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT64), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g027(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n453));
  NAND3_X1  g028(.A1(new_n437), .A2(new_n438), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(KEYINPUT65), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(new_n464), .A3(G125), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n460), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n460), .A2(G137), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n477));
  XOR2_X1   g052(.A(KEYINPUT3), .B(G2104), .Z(new_n478));
  OAI211_X1 g053(.A(new_n477), .B(new_n470), .C1(new_n478), .C2(new_n472), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n467), .A2(new_n476), .A3(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n481));
  OR3_X1    g056(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n460), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n478), .A2(G2105), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n484), .B(new_n487), .C1(G136), .C2(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(G114), .B2(new_n460), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n460), .A2(G138), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n461), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n461), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT68), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n501), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n503), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G166));
  NAND2_X1  g094(.A1(new_n504), .A2(new_n506), .ZN(new_n520));
  INV_X1    g095(.A(new_n502), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n520), .A2(new_n521), .A3(new_n515), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n513), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(new_n513), .A2(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n530), .B1(new_n516), .B2(new_n531), .C1(new_n532), .C2(new_n509), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  AND3_X1   g109(.A1(new_n520), .A2(G56), .A3(new_n521), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(G651), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n520), .A2(G81), .A3(new_n521), .A4(new_n515), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n513), .A2(G43), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(new_n512), .ZN(new_n549));
  NOR2_X1   g124(.A1(KEYINPUT6), .A2(G651), .ZN(new_n550));
  OAI211_X1 g125(.A(G53), .B(G543), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n515), .A2(new_n553), .A3(G53), .A4(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n507), .A2(G91), .A3(new_n515), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT69), .A2(G65), .ZN(new_n558));
  NOR2_X1   g133(.A1(KEYINPUT69), .A2(G65), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n520), .A2(new_n521), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n509), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n557), .A2(new_n563), .A3(KEYINPUT70), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n522), .A2(G91), .B1(new_n552), .B2(new_n554), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n562), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n564), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  OR2_X1    g146(.A1(new_n510), .A2(new_n518), .ZN(G303));
  AOI22_X1  g147(.A1(new_n522), .A2(G87), .B1(G49), .B2(new_n513), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n509), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n522), .A2(G86), .B1(G48), .B2(new_n513), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n509), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n513), .A2(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n516), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n513), .A2(G54), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n516), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n507), .A2(KEYINPUT10), .A3(G92), .A4(new_n515), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  AOI211_X1 g174(.A(new_n599), .B(new_n502), .C1(new_n504), .C2(new_n506), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT72), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT73), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n507), .A2(G66), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n605), .A2(new_n606), .A3(new_n602), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(G651), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n598), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n591), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n591), .B1(new_n610), .B2(G868), .ZN(G321));
  MUX2_X1   g187(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g188(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g189(.A(KEYINPUT74), .B(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n610), .B1(G860), .B2(new_n615), .ZN(G148));
  NAND2_X1  g191(.A1(new_n610), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n461), .A2(new_n469), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n488), .A2(G135), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n460), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT75), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n485), .A2(new_n629), .A3(G123), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n485), .B2(G123), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n626), .B1(new_n627), .B2(new_n628), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n623), .A2(new_n624), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(G2096), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n625), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT77), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n638), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT78), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT79), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n624), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(new_n685), .B(new_n684), .S(new_n677), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT80), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n687), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n674), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n690), .A2(new_n694), .A3(new_n674), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n697), .ZN(new_n700));
  INV_X1    g275(.A(new_n698), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n695), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G29), .B2(G32), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n488), .A2(G141), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT90), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n485), .A2(G129), .B1(G105), .B2(new_n469), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT92), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n706), .B1(new_n714), .B2(G29), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n713), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n715), .B1(KEYINPUT93), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n724), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT94), .Z(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G1966), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT31), .B(G11), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G28), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n718), .B1(new_n731), .B2(G28), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n730), .B1(new_n732), .B2(new_n733), .C1(new_n632), .C2(new_n718), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n724), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n724), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n734), .B1(new_n736), .B2(G1961), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n728), .A2(new_n729), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT95), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n718), .B1(new_n742), .B2(G34), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT88), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(KEYINPUT88), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n742), .B2(G34), .ZN(new_n746));
  AOI22_X1  g321(.A1(G160), .A2(G29), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G2084), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT89), .Z(new_n749));
  OR2_X1    g324(.A1(new_n747), .A2(G2084), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n718), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n718), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT29), .Z(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n750), .B1(G1961), .B2(new_n736), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n723), .A2(new_n740), .A3(new_n741), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n718), .A2(G26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G116), .B2(new_n460), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT85), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n488), .A2(G140), .B1(G128), .B2(new_n485), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n759), .B1(new_n765), .B2(new_n718), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT86), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n718), .A2(G33), .ZN(new_n769));
  NAND2_X1  g344(.A1(G115), .A2(G2104), .ZN(new_n770));
  INV_X1    g345(.A(G127), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n478), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n460), .B1(new_n772), .B2(KEYINPUT87), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(KEYINPUT87), .B2(new_n772), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n775));
  NAND2_X1  g350(.A1(G103), .A2(G2104), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G2105), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n488), .A2(G139), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n769), .B1(new_n780), .B2(new_n718), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n753), .A2(new_n754), .B1(G2072), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n724), .A2(G19), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n543), .B2(new_n724), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1341), .Z(new_n785));
  NOR2_X1   g360(.A1(new_n781), .A2(G2072), .ZN(new_n786));
  NOR2_X1   g361(.A1(G164), .A2(new_n718), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G27), .B2(new_n718), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n786), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AND4_X1   g367(.A1(new_n768), .A2(new_n782), .A3(new_n785), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G4), .A2(G16), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT84), .Z(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n609), .B2(new_n724), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1348), .ZN(new_n797));
  NAND2_X1  g372(.A1(G299), .A2(G16), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n724), .A2(G20), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT23), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G1956), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n793), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n757), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT83), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT34), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT83), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n810), .A2(new_n815), .A3(new_n811), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n724), .A2(G23), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n573), .A2(new_n574), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n724), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT33), .B(G1976), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n724), .A2(G22), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G166), .B2(new_n724), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1971), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n488), .A2(G131), .B1(G119), .B2(new_n485), .ZN(new_n827));
  OAI21_X1  g402(.A(KEYINPUT81), .B1(G95), .B2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NOR3_X1   g404(.A1(KEYINPUT81), .A2(G95), .A3(G2105), .ZN(new_n830));
  OAI221_X1 g405(.A(G2104), .B1(G107), .B2(new_n460), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  MUX2_X1   g407(.A(G25), .B(new_n832), .S(G29), .Z(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n724), .A2(G24), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n589), .B2(new_n724), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT82), .B(G1986), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  AND3_X1   g414(.A1(new_n826), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n813), .A2(new_n816), .A3(new_n825), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT34), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n845), .A3(new_n842), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n806), .B1(new_n844), .B2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n805), .ZN(G150));
  NAND2_X1  g424(.A1(new_n610), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  AOI211_X1 g427(.A(new_n852), .B(new_n502), .C1(new_n504), .C2(new_n506), .ZN(new_n853));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(G651), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n520), .A2(G93), .A3(new_n521), .A4(new_n515), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n513), .A2(G55), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n538), .A2(new_n856), .A3(new_n541), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n507), .A2(G56), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n509), .B1(new_n861), .B2(new_n536), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n539), .A2(new_n540), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n520), .A2(G67), .A3(new_n521), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n509), .B1(new_n864), .B2(new_n854), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(new_n858), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n862), .A2(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n851), .B(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n865), .A2(new_n866), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(new_n872), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(G145));
  NAND2_X1  g453(.A1(new_n497), .A2(new_n499), .ZN(new_n879));
  INV_X1    g454(.A(G114), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n491), .B1(new_n880), .B2(G2105), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(G126), .B2(new_n485), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n780), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(new_n765), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n765), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n717), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n717), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n485), .A2(G130), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n460), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(G142), .B2(new_n488), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n622), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n832), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n886), .A2(new_n887), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n714), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(G164), .A3(new_n888), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n891), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n898), .B1(new_n891), .B2(new_n901), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n903), .A3(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G160), .B(new_n632), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(G162), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  INV_X1    g488(.A(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n915), .B2(new_n905), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT40), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n907), .B2(new_n908), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n919), .A2(new_n920), .A3(new_n916), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n918), .A2(new_n921), .ZN(G395));
  XNOR2_X1  g497(.A(new_n818), .B(G166), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n589), .B1(new_n581), .B2(new_n582), .ZN(new_n924));
  INV_X1    g499(.A(new_n582), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n580), .A3(G290), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n923), .B1(new_n926), .B2(new_n924), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n929), .B(KEYINPUT42), .Z(new_n930));
  XNOR2_X1  g505(.A(new_n617), .B(new_n869), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT70), .B1(new_n557), .B2(new_n563), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n566), .A2(new_n568), .A3(new_n565), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n933), .A2(new_n934), .A3(new_n608), .A4(new_n598), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n933), .A2(new_n934), .B1(new_n598), .B2(new_n608), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n609), .B1(new_n569), .B2(new_n564), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n933), .A2(new_n934), .A3(new_n608), .A4(new_n598), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(KEYINPUT41), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(KEYINPUT98), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT98), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n932), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n931), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n942), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n931), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n930), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n930), .A2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(G868), .B2(new_n875), .ZN(G295));
  OAI21_X1  g526(.A(new_n950), .B1(G868), .B2(new_n875), .ZN(G331));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n860), .A2(new_n867), .A3(G301), .ZN(new_n954));
  AOI21_X1  g529(.A(G301), .B1(new_n860), .B2(new_n867), .ZN(new_n955));
  OAI21_X1  g530(.A(G286), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n868), .A2(G171), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n860), .A2(new_n867), .A3(G301), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(G168), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n953), .B1(new_n960), .B2(new_n946), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n941), .A3(new_n944), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(KEYINPUT100), .A3(new_n942), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n961), .A2(new_n962), .A3(new_n929), .A4(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI221_X4 g542(.A(new_n953), .B1(new_n939), .B2(new_n938), .C1(new_n956), .C2(new_n959), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT100), .B1(new_n963), .B2(new_n942), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n970), .A2(KEYINPUT101), .A3(new_n929), .A4(new_n962), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n974));
  INV_X1    g549(.A(new_n929), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT44), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n937), .A2(new_n940), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n960), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n946), .B2(new_n960), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n975), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n973), .B1(new_n972), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT102), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n972), .A2(new_n982), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n987), .A3(KEYINPUT44), .A4(new_n977), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n972), .A2(new_n976), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n972), .A2(new_n973), .A3(new_n982), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT99), .B(KEYINPUT44), .Z(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n995), .ZN(G397));
  XNOR2_X1  g571(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G164), .B2(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n476), .A2(new_n479), .A3(G40), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n998), .A2(new_n466), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT105), .ZN(new_n1001));
  INV_X1    g576(.A(G2067), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n765), .B(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n717), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n717), .A2(new_n1006), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n714), .A2(new_n1005), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(new_n1003), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1012), .B2(new_n1001), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n832), .B(new_n834), .Z(new_n1014));
  NAND2_X1  g589(.A1(new_n1001), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G290), .A2(G1986), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1000), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT48), .Z(new_n1019));
  OAI21_X1  g594(.A(new_n1009), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1013), .A2(new_n834), .A3(new_n831), .A4(new_n827), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n765), .A2(new_n1002), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1001), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT55), .ZN(new_n1026));
  NOR2_X1   g601(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT110), .B1(G164), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n883), .A2(new_n1030), .A3(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n466), .A2(new_n999), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1032), .A2(new_n754), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n879), .B2(new_n882), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT45), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n998), .A2(new_n1037), .A3(new_n1033), .ZN(new_n1038));
  INV_X1    g613(.A(G1971), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT111), .B(new_n1026), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1025), .B(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1042), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n577), .A2(new_n579), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n576), .A2(new_n509), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT108), .ZN(new_n1054));
  OAI21_X1  g629(.A(G1981), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n577), .A2(new_n1054), .A3(G1981), .A4(new_n579), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1051), .B1(new_n1059), .B2(KEYINPUT49), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1056), .A2(new_n1057), .A3(new_n1061), .A4(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(new_n999), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n467), .A2(new_n1063), .A3(new_n1036), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n573), .A2(G1976), .A3(new_n574), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(G8), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT107), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1066), .A2(new_n1070), .B1(G288), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1050), .A2(new_n1065), .A3(new_n1069), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1060), .A2(new_n1062), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT106), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n883), .B2(new_n1027), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT106), .B(new_n1028), .C1(new_n879), .C2(new_n882), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1033), .B(new_n1034), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1040), .B1(G2090), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n1047), .A3(G8), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n997), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1036), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(new_n1033), .C1(KEYINPUT45), .C2(new_n1036), .ZN(new_n1084));
  INV_X1    g659(.A(G1966), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT106), .B1(G164), .B2(new_n1028), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n883), .A2(new_n1075), .A3(new_n1027), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G2084), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G286), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1049), .A2(new_n1081), .A3(KEYINPUT112), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1043), .A2(new_n1074), .A3(new_n1048), .A4(new_n1080), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1094), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT63), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1079), .A2(G8), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1026), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1081), .A2(KEYINPUT63), .A3(new_n1094), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g680(.A(G1976), .B(G288), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1052), .A2(G1981), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1080), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1108), .A2(new_n1050), .B1(new_n1109), .B2(new_n1074), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G168), .A2(new_n1042), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1092), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n1084), .A2(new_n1114), .A3(G2078), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1038), .B2(G2078), .ZN(new_n1116));
  INV_X1    g691(.A(G1961), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1078), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1119), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1042), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1112), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1093), .A2(KEYINPUT118), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1122), .A2(KEYINPUT51), .A3(new_n1112), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1113), .B(new_n1120), .C1(new_n1129), .C2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1119), .A2(G171), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT62), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1034), .A2(new_n1033), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n802), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n566), .A2(new_n568), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n1139), .B(KEYINPUT57), .Z(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT56), .B(G2072), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n998), .A2(new_n1037), .A3(new_n1033), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1138), .A2(KEYINPUT113), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1140), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AND4_X1   g725(.A1(new_n1002), .A2(new_n467), .A3(new_n1063), .A4(new_n1036), .ZN(new_n1151));
  INV_X1    g726(.A(G1348), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1078), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT114), .B1(new_n1153), .B2(new_n609), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1153), .A2(KEYINPUT114), .A3(new_n609), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1147), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n609), .B1(new_n1153), .B2(KEYINPUT60), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1158), .A2(new_n1159), .B1(KEYINPUT60), .B2(new_n1153), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n543), .A2(KEYINPUT117), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT115), .B(G1996), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n998), .A2(new_n1037), .A3(new_n1033), .A4(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT58), .B(G1341), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1165), .B2(KEYINPUT116), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1165), .A2(KEYINPUT116), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1161), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1170), .B(new_n1161), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1150), .A2(KEYINPUT61), .A3(new_n1143), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1160), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT61), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1157), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1114), .B(G2078), .C1(new_n1036), .C2(KEYINPUT45), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n998), .A2(new_n1033), .A3(KEYINPUT122), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT122), .B1(new_n998), .B2(new_n1033), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT123), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1180), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n1178), .A4(new_n1177), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1118), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1078), .A2(KEYINPUT121), .A3(new_n1117), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1189), .A3(new_n1116), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1134), .B1(new_n1190), .B2(G171), .ZN(new_n1191));
  XOR2_X1   g766(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(G171), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT54), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(G301), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1191), .A2(new_n1192), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1135), .B1(new_n1176), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1113), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT51), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1130), .B1(new_n1201), .B2(KEYINPUT119), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1199), .B1(new_n1202), .B2(new_n1128), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1133), .B1(new_n1198), .B2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1097), .B(KEYINPUT124), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1111), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1017), .ZN(new_n1207));
  NAND2_X1  g782(.A1(G290), .A2(G1986), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1207), .A2(KEYINPUT104), .A3(new_n1208), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1209), .B(new_n1000), .C1(KEYINPUT104), .C2(new_n1208), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1013), .A2(new_n1015), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1024), .B1(new_n1206), .B2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g787(.A1(new_n670), .A2(G319), .A3(new_n671), .ZN(new_n1214));
  XNOR2_X1  g788(.A(new_n1214), .B(KEYINPUT125), .ZN(new_n1215));
  OR3_X1    g789(.A1(new_n1215), .A2(G401), .A3(KEYINPUT126), .ZN(new_n1216));
  OAI21_X1  g790(.A(KEYINPUT126), .B1(new_n1215), .B2(G401), .ZN(new_n1217));
  AND3_X1   g791(.A1(new_n1216), .A2(new_n703), .A3(new_n1217), .ZN(new_n1218));
  OAI211_X1 g792(.A(new_n993), .B(new_n1218), .C1(new_n919), .C2(new_n916), .ZN(G225));
  INV_X1    g793(.A(G225), .ZN(G308));
endmodule


