//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  MUX2_X1   g003(.A(G1gat), .B(new_n203), .S(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G43gat), .B(G50gat), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OR3_X1    g012(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(KEYINPUT91), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT91), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n215), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n214), .A2(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n213), .A2(new_n219), .B1(new_n220), .B2(new_n210), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT92), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT17), .Z(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n224), .B2(new_n206), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT18), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n206), .B(new_n221), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n226), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT93), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT11), .ZN(new_n238));
  INV_X1    g037(.A(G169gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT89), .B(G197gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n243));
  XOR2_X1   g042(.A(new_n242), .B(new_n243), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n236), .A2(new_n245), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250));
  NOR3_X1   g049(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n251), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n250), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(new_n252), .ZN(new_n262));
  OAI211_X1 g061(.A(KEYINPUT64), .B(new_n258), .C1(new_n262), .C2(new_n251), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  INV_X1    g063(.A(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT28), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n260), .A2(new_n263), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n265), .A2(new_n271), .B1(new_n252), .B2(KEYINPUT23), .ZN(new_n272));
  OR2_X1    g071(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(G190gat), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n254), .A2(KEYINPUT23), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT25), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n272), .A2(new_n277), .A3(new_n275), .A4(KEYINPUT25), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n270), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G127gat), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n284), .A2(KEYINPUT65), .A3(G134gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G134gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G127gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(G134gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT65), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G113gat), .ZN(new_n293));
  INV_X1    g092(.A(G113gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G120gat), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT1), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT66), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n285), .B1(new_n298), .B2(KEYINPUT65), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n295), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n297), .A2(new_n304), .B1(new_n296), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n296), .A2(new_n298), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n291), .A2(KEYINPUT66), .A3(new_n296), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n300), .B1(new_n299), .B2(new_n303), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n282), .A3(new_n270), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G227gat), .ZN(new_n313));
  INV_X1    g112(.A(G233gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G15gat), .B(G43gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(G71gat), .B(G99gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n313), .A2(new_n314), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n311), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n323), .B2(KEYINPUT32), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT33), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n325), .B1(new_n323), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(KEYINPUT68), .B(new_n324), .C1(new_n327), .C2(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n323), .A2(KEYINPUT32), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n321), .A2(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n318), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n336), .ZN(new_n338));
  AOI211_X1 g137(.A(new_n338), .B(new_n317), .C1(new_n331), .C2(new_n332), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT86), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n326), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT68), .B1(new_n344), .B2(new_n324), .ZN(new_n345));
  INV_X1    g144(.A(new_n332), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n336), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n317), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT86), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n336), .A3(new_n318), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n340), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT35), .ZN(new_n354));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT72), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n356), .B(KEYINPUT73), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n267), .A2(new_n263), .A3(new_n269), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n359), .A2(new_n260), .B1(new_n280), .B2(new_n281), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(KEYINPUT75), .B(new_n358), .C1(new_n360), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n270), .B2(new_n282), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(new_n357), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n283), .A2(new_n356), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G204gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G197gat), .ZN(new_n370));
  INV_X1    g169(.A(G197gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G204gat), .ZN(new_n372));
  INV_X1    g171(.A(G211gat), .ZN(new_n373));
  INV_X1    g172(.A(G218gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n370), .B(new_n372), .C1(new_n375), .C2(KEYINPUT22), .ZN(new_n376));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(KEYINPUT71), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n376), .B2(KEYINPUT71), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n368), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n360), .A2(new_n358), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n356), .B1(new_n283), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n383), .A2(new_n385), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n389), .A2(new_n380), .ZN(new_n397));
  INV_X1    g196(.A(new_n385), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n384), .B1(new_n368), .B2(new_n381), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n395), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT30), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n385), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n395), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n396), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  XOR2_X1   g209(.A(G155gat), .B(G162gat), .Z(new_n411));
  NAND2_X1  g210(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n414));
  OAI21_X1  g213(.A(G155gat), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(KEYINPUT2), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  INV_X1    g216(.A(G141gat), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT77), .B1(new_n418), .B2(G148gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(G148gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT77), .ZN(new_n424));
  INV_X1    g223(.A(G148gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(G141gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(G141gat), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(new_n422), .A3(new_n417), .A4(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n416), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G155gat), .B(G162gat), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n418), .A2(G148gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n427), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT3), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n430), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n440), .A3(new_n310), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n422), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n428), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n435), .B1(new_n445), .B2(new_n416), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n305), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(KEYINPUT4), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n305), .B2(new_n446), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n441), .B(new_n442), .C1(new_n448), .C2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n310), .A2(new_n437), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n447), .ZN(new_n454));
  INV_X1    g253(.A(new_n442), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n456), .A3(KEYINPUT80), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT81), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n447), .B2(KEYINPUT4), .ZN(new_n463));
  INV_X1    g262(.A(new_n450), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n455), .A2(KEYINPUT5), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n441), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n410), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n451), .A2(new_n456), .A3(KEYINPUT80), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT80), .B1(new_n451), .B2(new_n456), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n469), .B(new_n410), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n406), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(new_n410), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n405), .ZN(new_n479));
  AND4_X1   g278(.A1(new_n354), .A2(new_n404), .A3(new_n475), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT3), .B1(new_n380), .B2(new_n387), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n362), .B1(new_n446), .B2(new_n439), .ZN(new_n484));
  OAI221_X1 g283(.A(new_n482), .B1(new_n483), .B2(new_n446), .C1(new_n380), .C2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n362), .B1(new_n376), .B2(new_n377), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n377), .B2(new_n376), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n446), .B1(new_n439), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT83), .B1(new_n484), .B2(new_n380), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n490));
  AOI211_X1 g289(.A(KEYINPUT3), .B(new_n435), .C1(new_n445), .C2(new_n416), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n381), .B(new_n490), .C1(new_n491), .C2(new_n362), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n485), .B1(new_n493), .B2(new_n482), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(G22gat), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n485), .C1(new_n493), .C2(new_n482), .ZN(new_n497));
  XNOR2_X1  g296(.A(G78gat), .B(G106gat), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n495), .B2(new_n497), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT31), .B(G50gat), .Z(new_n501));
  NOR3_X1   g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  INV_X1    g302(.A(new_n498), .ZN(new_n504));
  INV_X1    g303(.A(new_n488), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n440), .A2(new_n361), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n490), .B1(new_n506), .B2(new_n381), .ZN(new_n507));
  AOI211_X1 g306(.A(KEYINPUT83), .B(new_n380), .C1(new_n440), .C2(new_n361), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n481), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n496), .B1(new_n510), .B2(new_n485), .ZN(new_n511));
  INV_X1    g310(.A(new_n497), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n502), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n352), .A2(new_n353), .A3(new_n480), .A4(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n340), .A3(new_n351), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n404), .A2(new_n475), .A3(new_n354), .A4(new_n479), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT87), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n337), .A2(new_n339), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n404), .A2(new_n475), .A3(new_n479), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT35), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n441), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n465), .B2(new_n466), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n455), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n453), .A2(new_n447), .A3(new_n442), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT39), .B(new_n531), .C1(new_n527), .C2(new_n442), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n532), .A3(new_n410), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT40), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(KEYINPUT84), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(KEYINPUT84), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n530), .A2(new_n532), .A3(new_n410), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(new_n478), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n405), .B1(new_n478), .B2(new_n473), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n470), .A2(new_n406), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n400), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT38), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n402), .A2(new_n397), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT37), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n395), .B1(new_n390), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n368), .B2(new_n381), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n381), .B1(new_n386), .B2(new_n388), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n368), .A2(new_n547), .A3(new_n381), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT37), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n545), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n394), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n544), .A2(new_n546), .B1(new_n554), .B2(new_n542), .ZN(new_n555));
  OAI221_X1 g354(.A(new_n516), .B1(new_n538), .B2(new_n404), .C1(new_n541), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT70), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n337), .B2(new_n339), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  INV_X1    g360(.A(new_n516), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n523), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n556), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n525), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT88), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n525), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n249), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G183gat), .B(G211gat), .Z(new_n570));
  OR2_X1    g369(.A1(G57gat), .A2(G64gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G57gat), .A2(G64gat), .ZN(new_n572));
  AND2_X1   g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(KEYINPUT9), .ZN(new_n574));
  XNOR2_X1  g373(.A(G71gat), .B(G78gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT94), .Z(new_n577));
  XOR2_X1   g376(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT20), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n577), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n207), .B1(new_n590), .B2(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n589), .A2(new_n591), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n570), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  INV_X1    g395(.A(new_n570), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G134gat), .B(G162gat), .Z(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT7), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(KEYINPUT98), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  INV_X1    g408(.A(G92gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(KEYINPUT8), .A2(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G99gat), .B(G106gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT99), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n615), .A2(new_n221), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT102), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n614), .A2(KEYINPUT99), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n614), .A2(KEYINPUT99), .ZN(new_n620));
  OR3_X1    g419(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n615), .A2(KEYINPUT100), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n622), .A3(new_n224), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n623), .A2(KEYINPUT101), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(KEYINPUT101), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT97), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n627), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n618), .A2(new_n624), .A3(new_n625), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n631), .B1(new_n628), .B2(new_n633), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n600), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  INV_X1    g437(.A(new_n600), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n577), .A2(new_n614), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n612), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n613), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n613), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n576), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT105), .Z(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n648), .A2(KEYINPUT10), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n590), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n649), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n658), .A2(new_n660), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n649), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n655), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n569), .A2(new_n599), .A3(new_n641), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n475), .A2(new_n479), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g475(.A1(new_n672), .A2(new_n404), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(KEYINPUT42), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n677), .B(KEYINPUT106), .Z(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(G8gat), .ZN(new_n682));
  OAI221_X1 g481(.A(new_n679), .B1(KEYINPUT42), .B2(new_n678), .C1(new_n680), .C2(new_n682), .ZN(G1325gat));
  AOI21_X1  g482(.A(G15gat), .B1(new_n673), .B2(new_n352), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n560), .A2(new_n561), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G15gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT107), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n673), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n516), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NOR3_X1   g490(.A1(new_n599), .A2(new_n641), .A3(new_n670), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n525), .A2(new_n567), .A3(new_n564), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n567), .B1(new_n525), .B2(new_n564), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n248), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n674), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n695), .A2(G29gat), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT45), .Z(new_n698));
  INV_X1    g497(.A(new_n641), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n693), .B2(new_n694), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n641), .B1(new_n525), .B2(new_n564), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT44), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n599), .A2(new_n249), .A3(new_n670), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT108), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n701), .A2(new_n703), .A3(new_n707), .A4(new_n704), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n674), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G29gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n698), .A2(new_n710), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n695), .A2(G36gat), .A3(new_n404), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  INV_X1    g512(.A(new_n404), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n706), .A2(new_n714), .A3(new_n708), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G36gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(new_n685), .ZN(new_n720));
  OAI21_X1  g519(.A(G43gat), .B1(new_n705), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  INV_X1    g521(.A(new_n352), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(G43gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n722), .B1(new_n695), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n569), .A2(KEYINPUT110), .A3(new_n692), .A4(new_n724), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n721), .A2(new_n728), .A3(KEYINPUT47), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n726), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n726), .B2(new_n727), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n706), .A2(new_n685), .A3(new_n708), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G43gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT112), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n739), .B(KEYINPUT47), .C1(new_n733), .C2(new_n735), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n729), .B1(new_n738), .B2(new_n740), .ZN(G1330gat));
  NOR3_X1   g540(.A1(new_n695), .A2(G50gat), .A3(new_n516), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G50gat), .B1(new_n705), .B2(new_n516), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n706), .A2(new_n562), .A3(new_n708), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n742), .B1(new_n747), .B2(G50gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n748), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g548(.A1(new_n599), .A2(new_n641), .A3(new_n249), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n671), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n565), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n696), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT113), .B(G57gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1332gat));
  AOI211_X1 g554(.A(new_n404), .B(new_n752), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT114), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n756), .B(new_n758), .ZN(G1333gat));
  INV_X1    g558(.A(new_n752), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(G71gat), .A3(new_n685), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n752), .A2(new_n723), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(G71gat), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n760), .A2(new_n562), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n599), .A2(new_n248), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n701), .A2(new_n703), .A3(new_n670), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n696), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n702), .A2(new_n768), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT51), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n670), .A2(new_n609), .A3(new_n674), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n769), .B2(new_n404), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n670), .A2(new_n610), .A3(new_n714), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n769), .B2(new_n720), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n723), .A2(G99gat), .A3(new_n671), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n772), .B2(new_n780), .ZN(G1338gat));
  OAI21_X1  g580(.A(G106gat), .B1(new_n769), .B2(new_n516), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n671), .A2(G106gat), .A3(new_n516), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n772), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g584(.A(new_n599), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n655), .B1(new_n667), .B2(KEYINPUT54), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT54), .B1(new_n666), .B2(new_n649), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n664), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n665), .B1(new_n790), .B2(KEYINPUT55), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n650), .B1(new_n658), .B2(new_n660), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n656), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n663), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n650), .B1(new_n795), .B2(new_n661), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n794), .B(KEYINPUT55), .C1(new_n796), .C2(new_n788), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n225), .A2(new_n226), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n231), .A2(new_n232), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n242), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n246), .A2(new_n802), .ZN(new_n803));
  AND4_X1   g602(.A1(new_n640), .A2(new_n799), .A3(new_n637), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n794), .B1(new_n796), .B2(new_n788), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n805), .A2(new_n806), .B1(new_n664), .B2(new_n657), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n248), .A3(new_n797), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n803), .A2(new_n670), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n637), .A2(new_n640), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n786), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n599), .A2(new_n641), .A3(new_n249), .A4(new_n671), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n696), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n404), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n522), .ZN(new_n817));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n248), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n518), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n249), .A2(new_n294), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(G1340gat));
  AOI21_X1  g620(.A(G120gat), .B1(new_n817), .B2(new_n670), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n671), .A2(new_n292), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n819), .B2(new_n823), .ZN(G1341gat));
  NAND3_X1  g623(.A1(new_n817), .A2(new_n284), .A3(new_n599), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n816), .A2(new_n518), .A3(new_n786), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n284), .ZN(G1342gat));
  NOR2_X1   g626(.A1(new_n641), .A2(new_n714), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n815), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(G134gat), .A3(new_n522), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT56), .ZN(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n829), .B2(new_n518), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1343gat));
  NOR2_X1   g632(.A1(new_n685), .A2(new_n516), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT118), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n249), .A2(G141gat), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n815), .A2(new_n838), .A3(new_n834), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n836), .A2(new_n404), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT116), .B1(new_n791), .B2(new_n798), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n807), .A2(new_n842), .A3(new_n797), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n249), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n809), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n641), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n804), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n599), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n812), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n562), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT57), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n720), .A2(new_n674), .A3(new_n404), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n516), .B1(new_n811), .B2(new_n812), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n248), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  XOR2_X1   g656(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n858));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n856), .A2(new_n860), .A3(G141gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n856), .B2(G141gat), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n835), .A2(G141gat), .A3(new_n249), .A4(new_n714), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n859), .B1(new_n864), .B2(new_n865), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n425), .A2(KEYINPUT59), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n855), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT120), .B(new_n867), .C1(new_n868), .C2(new_n671), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n562), .A2(new_n854), .ZN(new_n870));
  INV_X1    g669(.A(new_n803), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  INV_X1    g671(.A(new_n799), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n641), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n637), .A2(new_n799), .A3(new_n640), .A4(KEYINPUT121), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n841), .A2(new_n843), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n248), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n699), .B1(new_n878), .B2(new_n809), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n786), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n870), .B1(new_n880), .B2(new_n812), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n853), .A2(new_n854), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n852), .A2(new_n671), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n425), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n869), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n868), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n670), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT120), .B1(new_n889), .B2(new_n867), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n836), .A2(new_n839), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n404), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n670), .A2(new_n425), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n887), .A2(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n868), .B2(new_n786), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n786), .A2(G155gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n892), .B2(new_n896), .ZN(G1346gat));
  NOR2_X1   g696(.A1(new_n413), .A2(new_n414), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n891), .A2(new_n898), .A3(new_n828), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n888), .A2(new_n699), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n900), .A2(KEYINPUT122), .B1(new_n414), .B2(new_n413), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(KEYINPUT122), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n674), .A2(new_n404), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n813), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(new_n518), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(new_n239), .A3(new_n249), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n905), .A2(new_n522), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n248), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n910), .B2(new_n239), .ZN(G1348gat));
  OAI21_X1  g710(.A(G176gat), .B1(new_n906), .B2(new_n671), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n671), .A2(G176gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n908), .B2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n906), .B2(new_n786), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n599), .A2(new_n264), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n906), .B2(new_n641), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n909), .A2(new_n265), .A3(new_n699), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1351gat));
  OR3_X1    g723(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT124), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT124), .B1(new_n881), .B2(new_n882), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n720), .A2(new_n904), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n371), .A3(new_n249), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n813), .A2(new_n834), .A3(new_n904), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n248), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n930), .A2(new_n933), .ZN(G1352gat));
  OAI21_X1  g733(.A(G204gat), .B1(new_n929), .B2(new_n671), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n670), .A2(new_n369), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n931), .A2(KEYINPUT125), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n931), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n935), .B(new_n940), .C1(new_n943), .C2(new_n944), .ZN(G1353gat));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n373), .A3(new_n599), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n786), .A2(new_n927), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  OR3_X1    g747(.A1(new_n881), .A2(new_n882), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n881), .A2(new_n882), .A3(new_n948), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n373), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n950), .A2(new_n953), .A3(KEYINPUT63), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n950), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n946), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n929), .B2(new_n641), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n932), .A2(new_n374), .A3(new_n699), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


