//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT67), .B(G96), .Z(G221));
  XOR2_X1   g012(.A(KEYINPUT68), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT69), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n461), .B1(new_n466), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AOI211_X1 g043(.A(KEYINPUT70), .B(new_n468), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n468), .C1(new_n462), .C2(new_n463), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G137), .A4(new_n468), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n471), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n462), .A2(new_n463), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n468), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT73), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n474), .A2(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n474), .A2(new_n486), .A3(new_n468), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n468), .A2(G112), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n483), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT74), .ZN(G162));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(KEYINPUT75), .A3(new_n499), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n468), .C1(new_n462), .C2(new_n463), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n474), .A2(new_n506), .A3(G138), .A4(new_n468), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n502), .A2(new_n503), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT6), .B1(new_n510), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(new_n509), .ZN(new_n518));
  NAND3_X1  g093(.A1(KEYINPUT77), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n512), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n520), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n514), .A2(G51), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n524), .A2(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n520), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n514), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT79), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n524), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n526), .B1(new_n548), .B2(KEYINPUT78), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n549), .B1(KEYINPUT78), .B2(new_n548), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n544), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT80), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n557), .B(new_n553), .C1(new_n546), .C2(new_n554), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(G651), .A3(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n520), .A2(G81), .B1(new_n514), .B2(G43), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT81), .Z(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(KEYINPUT82), .B2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(new_n513), .ZN(new_n571));
  OAI211_X1 g146(.A(G543), .B(new_n570), .C1(new_n571), .C2(new_n511), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n514), .A2(new_n576), .A3(new_n570), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n520), .A2(G91), .ZN(new_n578));
  INV_X1    g153(.A(G65), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n518), .B2(new_n519), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n583), .ZN(G299));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND2_X1  g160(.A1(new_n520), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n514), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AND2_X1   g164(.A1(new_n524), .A2(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT83), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n520), .A2(G86), .B1(new_n514), .B2(G48), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n526), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(new_n514), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI221_X1 g175(.A(new_n597), .B1(new_n598), .B2(new_n599), .C1(new_n600), .C2(new_n521), .ZN(G290));
  NAND2_X1  g176(.A1(new_n520), .A2(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n546), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT84), .B1(new_n610), .B2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  MUX2_X1   g187(.A(KEYINPUT84), .B(new_n611), .S(new_n612), .Z(G284));
  MUX2_X1   g188(.A(KEYINPUT84), .B(new_n611), .S(new_n612), .Z(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n610), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n610), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n562), .ZN(G323));
  XOR2_X1   g198(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n624));
  XNOR2_X1  g199(.A(G323), .B(new_n624), .ZN(G282));
  XNOR2_X1  g200(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n631), .A2(KEYINPUT87), .A3(G2105), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT87), .B1(new_n631), .B2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n481), .A2(G123), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n488), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n629), .A2(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(G2096), .ZN(new_n641));
  NAND4_X1  g216(.A1(new_n630), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT89), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2451), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT92), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT91), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2427), .B(G2430), .Z(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n648), .B(new_n655), .Z(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT90), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2454), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT93), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n664), .A2(new_n665), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT94), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n670), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n681), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  AOI211_X1 g260(.A(new_n683), .B(new_n685), .C1(new_n678), .C2(new_n682), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G305), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G6), .B2(G16), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G23), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G288), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n695), .A2(new_n696), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n697), .B(new_n702), .C1(new_n700), .C2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT97), .B(G16), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n703), .A2(new_n708), .A3(KEYINPUT34), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT34), .B1(new_n703), .B2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n481), .A2(G119), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n468), .A2(G107), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(G131), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n713), .B1(new_n714), .B2(new_n715), .C1(new_n488), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT95), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n712), .B1(new_n719), .B2(new_n711), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT96), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n720), .B(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G24), .B(G290), .S(new_n705), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT98), .B(G1986), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n709), .A2(new_n710), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT99), .A2(KEYINPUT36), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  NAND3_X1  g305(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT25), .Z(new_n732));
  INV_X1    g307(.A(G139), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n488), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT100), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n474), .A2(G127), .ZN(new_n736));
  AND2_X1   g311(.A1(G115), .A2(G2104), .ZN(new_n737));
  OAI21_X1  g312(.A(G2105), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G33), .B(new_n739), .S(G29), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT101), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2072), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT30), .B(G28), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n743), .A2(new_n711), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n638), .B2(new_n711), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT103), .Z(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT102), .B(KEYINPUT24), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(new_n711), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n478), .B2(new_n711), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n748), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n610), .B2(G16), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n754), .B1(G1348), .B2(new_n756), .C1(new_n749), .C2(new_n753), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n711), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n711), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT29), .B(G2090), .Z(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n757), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT26), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n765), .B(new_n767), .C1(G129), .C2(new_n481), .ZN(new_n768));
  INV_X1    g343(.A(G141), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n488), .B2(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G32), .B(new_n770), .S(G29), .Z(new_n771));
  XOR2_X1   g346(.A(KEYINPUT27), .B(G1996), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G21), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G168), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1966), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n562), .A2(new_n704), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G19), .B2(new_n704), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G1341), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n711), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n489), .A2(G140), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(G116), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G2105), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n481), .B2(G128), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(G2067), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G1348), .B2(new_n756), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n711), .A2(G27), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G164), .B2(new_n711), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G2078), .Z(new_n796));
  NAND4_X1  g371(.A1(new_n777), .A2(new_n781), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G171), .A2(new_n698), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G5), .B2(new_n698), .ZN(new_n799));
  INV_X1    g374(.A(G1961), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G1341), .B2(new_n780), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n704), .A2(G20), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT23), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n616), .B2(new_n698), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1956), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n797), .A2(new_n802), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n730), .A2(new_n742), .A3(new_n764), .A4(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  NAND2_X1  g385(.A1(new_n610), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT38), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n514), .A2(G55), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n521), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n526), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n561), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n559), .A3(new_n560), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n812), .B(new_n822), .Z(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n818), .A2(new_n825), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(G145));
  XNOR2_X1  g405(.A(G162), .B(new_n638), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n478), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n789), .B(new_n770), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n739), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n505), .A2(new_n507), .ZN(new_n835));
  INV_X1    g410(.A(new_n500), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n834), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n481), .A2(G130), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT104), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n489), .A2(G142), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n468), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n718), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n628), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n838), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT105), .ZN(new_n848));
  INV_X1    g423(.A(new_n838), .ZN(new_n849));
  INV_X1    g424(.A(new_n846), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(KEYINPUT105), .A3(new_n850), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n832), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n847), .A3(new_n832), .ZN(new_n855));
  INV_X1    g430(.A(G37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(G395));
  INV_X1    g435(.A(G868), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n819), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n863));
  XNOR2_X1  g438(.A(G290), .B(new_n693), .ZN(new_n864));
  XNOR2_X1  g439(.A(G166), .B(G288), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI211_X1 g441(.A(KEYINPUT107), .B(new_n863), .C1(new_n866), .C2(KEYINPUT108), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT107), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n866), .B2(KEYINPUT107), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n822), .B(new_n621), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n609), .A2(G299), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n616), .B1(new_n604), .B2(new_n608), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(new_n876), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(KEYINPUT41), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n875), .B2(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n878), .B(KEYINPUT106), .C1(new_n874), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(KEYINPUT106), .B2(new_n878), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n873), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n862), .B1(new_n887), .B2(new_n861), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT109), .ZN(G295));
  XNOR2_X1  g464(.A(new_n888), .B(KEYINPUT110), .ZN(G331));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n820), .A2(G301), .A3(new_n821), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G301), .B1(new_n820), .B2(new_n821), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n893), .A2(G286), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n822), .A2(G171), .ZN(new_n896));
  AOI21_X1  g471(.A(G168), .B1(new_n896), .B2(new_n892), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n895), .A2(new_n897), .A3(new_n884), .ZN(new_n898));
  INV_X1    g473(.A(new_n877), .ZN(new_n899));
  OAI21_X1  g474(.A(G286), .B1(new_n893), .B2(new_n894), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(G168), .A3(new_n892), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n869), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n856), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n877), .B1(new_n895), .B2(new_n897), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n900), .A2(new_n901), .A3(new_n883), .A4(new_n881), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n866), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT111), .B1(new_n908), .B2(G37), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n907), .A3(new_n866), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n905), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(new_n856), .A3(new_n911), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n891), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n905), .A2(new_n909), .A3(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT43), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n916), .B2(KEYINPUT43), .ZN(new_n919));
  AND4_X1   g494(.A1(new_n910), .A2(new_n903), .A3(new_n856), .A4(new_n911), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n915), .B1(new_n921), .B2(new_n891), .ZN(G397));
  NAND2_X1  g497(.A1(new_n789), .A2(G2067), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n784), .A2(new_n791), .A3(new_n788), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n719), .A2(new_n723), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n770), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n718), .A2(new_n722), .ZN(new_n929));
  AND4_X1   g504(.A1(new_n925), .A2(new_n926), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G1384), .B1(new_n835), .B2(new_n836), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT45), .B1(new_n932), .B2(KEYINPUT113), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(KEYINPUT113), .B2(new_n932), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n477), .B(G40), .C1(new_n467), .C2(new_n469), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  OR3_X1    g513(.A1(new_n937), .A2(G1986), .A3(G290), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(KEYINPUT48), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(KEYINPUT48), .B2(new_n940), .ZN(new_n942));
  INV_X1    g517(.A(new_n925), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n936), .B1(new_n943), .B2(new_n770), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n937), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n936), .B2(new_n927), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n925), .A2(new_n928), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n924), .B1(new_n926), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n936), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n942), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n932), .A2(new_n935), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1981), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n693), .A2(KEYINPUT116), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n593), .A2(new_n594), .A3(new_n958), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n959), .A2(new_n962), .B1(G1981), .B2(G305), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(KEYINPUT49), .ZN(new_n967));
  AOI211_X1 g542(.A(G1976), .B(G288), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n959), .A2(new_n962), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n956), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G164), .B2(G1384), .ZN(new_n973));
  INV_X1    g548(.A(new_n935), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n931), .A2(KEYINPUT45), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1971), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n502), .A2(new_n503), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n835), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n495), .A2(KEYINPUT75), .A3(new_n499), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT75), .B1(new_n495), .B2(new_n499), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n835), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n837), .A2(new_n982), .A3(new_n987), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT114), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n931), .A2(new_n993), .A3(new_n982), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n935), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n978), .B1(new_n996), .B2(G2090), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(G303), .A2(G8), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT55), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n956), .B(new_n1003), .C1(new_n1002), .C2(G288), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n956), .B1(new_n1002), .B2(G288), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n966), .B2(new_n967), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n971), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1012));
  NAND3_X1  g587(.A1(new_n986), .A2(new_n982), .A3(new_n987), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n500), .B1(new_n505), .B2(new_n507), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT50), .B1(new_n1014), .B2(G1384), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n974), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n978), .B1(G2090), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1000), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1001), .A2(new_n1009), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n974), .B(new_n1021), .C1(KEYINPUT45), .C2(new_n931), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n990), .A2(new_n749), .A3(new_n995), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(KEYINPUT117), .A3(new_n1023), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(G8), .A3(G168), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1012), .B1(new_n1020), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT63), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n998), .A2(new_n1000), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1001), .A3(new_n1009), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1011), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT62), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1029), .A2(G286), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1026), .A2(new_n1027), .A3(G168), .A4(new_n1028), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(KEYINPUT51), .A3(G8), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT127), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(G8), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1037), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT127), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT62), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n996), .A2(new_n800), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n976), .B2(G2078), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1022), .A2(new_n1053), .A3(G2078), .ZN(new_n1056));
  OAI21_X1  g631(.A(G171), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1020), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1047), .A2(new_n1051), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1036), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G2078), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n466), .B2(G2105), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n975), .A2(new_n1063), .A3(new_n477), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n934), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1052), .A2(G301), .A3(new_n1054), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT54), .B1(new_n1057), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1020), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G301), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1055), .B1(new_n934), .B2(new_n1064), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1070), .B(KEYINPUT54), .C1(G301), .C2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1068), .A2(new_n1049), .A3(new_n1050), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1348), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT115), .B1(new_n988), .B2(KEYINPUT50), .ZN(new_n1075));
  AOI211_X1 g650(.A(new_n979), .B(new_n982), .C1(new_n986), .C2(new_n987), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n993), .B1(new_n931), .B2(new_n982), .ZN(new_n1078));
  NOR4_X1   g653(.A1(new_n1014), .A2(KEYINPUT114), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n974), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1074), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n954), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(G2067), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1348), .B1(new_n990), .B2(new_n995), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1083), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n610), .B1(new_n1090), .B2(KEYINPUT124), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1086), .A3(new_n609), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1087), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1088), .A2(new_n1083), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT125), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1087), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1085), .A2(new_n1086), .A3(new_n609), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n609), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1095), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n973), .A2(new_n974), .A3(new_n927), .A4(new_n975), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n932), .B2(new_n935), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n559), .A2(KEYINPUT119), .A3(new_n560), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT120), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1113), .A3(new_n1109), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT120), .B(new_n1108), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT59), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1016), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  XNOR2_X1  g699(.A(G299), .B(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1120), .A2(new_n1125), .A3(new_n1122), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(KEYINPUT121), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT61), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1115), .A2(new_n1118), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1128), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1120), .A2(KEYINPUT122), .A3(new_n1125), .A4(new_n1122), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1135), .A2(KEYINPUT123), .A3(KEYINPUT61), .A4(new_n1136), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1133), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1096), .A2(new_n1103), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1127), .B1(new_n1094), .B2(new_n609), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1128), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1073), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(KEYINPUT126), .A3(new_n1144), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1060), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(G290), .B(G1986), .Z(new_n1150));
  AOI21_X1  g725(.A(new_n937), .B1(new_n930), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n953), .B1(new_n1149), .B2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g727(.A1(new_n854), .A2(new_n857), .ZN(new_n1154));
  OR2_X1    g728(.A1(G227), .A2(new_n459), .ZN(new_n1155));
  NOR3_X1   g729(.A1(G229), .A2(G401), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g731(.A1(new_n1157), .A2(new_n921), .ZN(G308));
  OR2_X1    g732(.A1(new_n919), .A2(new_n920), .ZN(new_n1159));
  OAI211_X1 g733(.A(new_n1154), .B(new_n1156), .C1(new_n1159), .C2(new_n918), .ZN(G225));
endmodule


