//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G232), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n202), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G77), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n212), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n206), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n225), .B(new_n228), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n208), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  INV_X1    g0052(.A(G20), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n252), .A2(new_n253), .A3(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n229), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  AND3_X1   g0059(.A1(new_n257), .A2(G50), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n203), .A2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n253), .A2(G33), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT68), .B1(G20), .B2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR3_X1   g0065(.A1(KEYINPUT68), .A2(G20), .A3(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G150), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n261), .B1(new_n262), .B2(new_n263), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n260), .B1(new_n269), .B2(new_n256), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n254), .A2(new_n202), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT72), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n272), .B(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(KEYINPUT67), .B2(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G223), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G222), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n290), .B(new_n283), .C1(G77), .C2(new_n286), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n283), .A2(new_n279), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G226), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(G200), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n273), .A2(new_n274), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n276), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n302), .A3(new_n297), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n301), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n276), .A2(new_n305), .A3(new_n299), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n208), .A2(G1698), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n308), .B1(G226), .B2(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G97), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n283), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n282), .A2(new_n284), .B1(G238), .B2(new_n292), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT14), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(G179), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(G169), .C1(new_n320), .C2(new_n321), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n266), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n264), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n331));
  INV_X1    g0131(.A(G77), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n262), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n256), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT11), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n252), .A2(G1), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G20), .A3(new_n221), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT12), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT69), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n256), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n337), .A2(G20), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(G68), .A3(new_n259), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n333), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n336), .A2(new_n339), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n328), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n322), .A2(G190), .ZN(new_n351));
  INV_X1    g0151(.A(new_n349), .ZN(new_n352));
  OAI21_X1  g0152(.A(G200), .B1(new_n320), .B2(new_n321), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n294), .A2(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n294), .A2(new_n323), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n272), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n307), .A2(new_n350), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT3), .A2(G33), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n253), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(KEYINPUT7), .A3(new_n253), .A4(new_n360), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n221), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(G58), .B(G68), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G20), .ZN(new_n367));
  INV_X1    g0167(.A(G159), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n267), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT16), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n309), .A2(new_n310), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT7), .B1(new_n371), .B2(new_n253), .ZN(new_n372));
  NOR4_X1   g0172(.A1(new_n309), .A2(new_n310), .A3(new_n362), .A4(G20), .ZN(new_n373));
  OAI21_X1  g0173(.A(G68), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n330), .A2(G159), .B1(new_n366), .B2(G20), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT75), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n378), .A3(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n374), .A2(new_n378), .A3(new_n376), .A4(new_n375), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n256), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n263), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n259), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n384), .A2(new_n344), .B1(new_n343), .B2(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n213), .A2(G1698), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n286), .B(new_n388), .C1(G223), .C2(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n283), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n292), .A2(G232), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n392), .A2(new_n285), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n323), .B2(new_n394), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n387), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT18), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n387), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n389), .A2(new_n390), .ZN(new_n402));
  INV_X1    g0202(.A(new_n283), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n285), .B(new_n393), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G200), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G190), .B2(new_n404), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n386), .A3(new_n382), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n407), .A2(new_n382), .A3(KEYINPUT17), .A4(new_n386), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n288), .A2(G232), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n286), .B(new_n413), .C1(new_n222), .C2(new_n288), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n283), .C1(G107), .C2(new_n286), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n292), .A2(new_n218), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n285), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G200), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n295), .B2(new_n417), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n346), .A2(G77), .A3(new_n259), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n254), .A2(new_n332), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n267), .A2(new_n263), .B1(new_n253), .B2(new_n332), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT15), .B(G87), .Z(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n262), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n256), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n417), .A2(new_n323), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT71), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT71), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n432), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G179), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n415), .A2(new_n285), .A3(new_n435), .A4(new_n416), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT70), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n428), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n401), .A2(new_n412), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n358), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n214), .A2(KEYINPUT6), .A3(G97), .ZN(new_n441));
  INV_X1    g0241(.A(G97), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(new_n214), .ZN(new_n443));
  NOR2_X1   g0243(.A1(G97), .A2(G107), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n441), .B1(new_n445), .B2(KEYINPUT6), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G20), .ZN(new_n447));
  OAI21_X1  g0247(.A(G107), .B1(new_n372), .B2(new_n373), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n330), .A2(G77), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(new_n256), .B1(new_n442), .B2(new_n254), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n258), .A2(G33), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n257), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G97), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(G244), .B(new_n288), .C1(new_n309), .C2(new_n310), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT4), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(G250), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT76), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n286), .A2(KEYINPUT76), .A3(G250), .A4(G1698), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n283), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n258), .B(G45), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n403), .A2(new_n472), .A3(G257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT77), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT77), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n403), .A2(new_n472), .A3(new_n475), .A4(G257), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n278), .A2(G1), .ZN(new_n478));
  OAI211_X1 g0278(.A(G274), .B(new_n478), .C1(new_n470), .C2(new_n471), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n323), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n468), .A2(new_n477), .A3(new_n435), .A4(new_n479), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n456), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(G200), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n468), .A2(new_n477), .A3(G190), .A4(new_n479), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n451), .A3(new_n455), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n461), .B(new_n253), .C1(G33), .C2(new_n442), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT79), .B(G116), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n256), .B(new_n488), .C1(new_n489), .C2(new_n253), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT20), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n491), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT69), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n257), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G116), .B(new_n452), .C1(new_n496), .C2(new_n340), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n343), .A2(new_n489), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n288), .A2(G257), .ZN(new_n500));
  OAI221_X1 g0300(.A(new_n500), .B1(new_n215), .B2(new_n288), .C1(new_n309), .C2(new_n310), .ZN(new_n501));
  INV_X1    g0301(.A(G303), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n371), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n503), .A3(new_n283), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n403), .A2(new_n472), .A3(G270), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n479), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n506), .A2(G169), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT82), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(KEYINPUT21), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n510), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n499), .A2(new_n512), .A3(new_n507), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n504), .A2(new_n505), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n499), .A2(G179), .A3(new_n479), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n341), .B2(new_n345), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(new_n452), .B1(new_n492), .B2(new_n493), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(G190), .A3(new_n479), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n506), .A2(G200), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n498), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n511), .A2(new_n513), .A3(new_n515), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n487), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n214), .A2(G20), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT23), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n253), .B(G87), .C1(new_n309), .C2(new_n310), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n286), .A2(new_n528), .A3(new_n253), .A4(G87), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n489), .A2(new_n253), .A3(G33), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n256), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n524), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n337), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT25), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n454), .A2(G107), .B1(new_n540), .B2(new_n539), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n536), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n403), .A2(new_n472), .A3(G264), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n545), .A2(new_n479), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n210), .A2(new_n288), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n286), .B(new_n547), .C1(G257), .C2(new_n288), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n403), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT83), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI211_X1 g0352(.A(KEYINPUT83), .B(new_n403), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n546), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G169), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n545), .A2(new_n479), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n550), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G179), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n544), .A2(new_n559), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n554), .A2(G190), .B1(G200), .B2(new_n557), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(new_n536), .A3(new_n542), .A4(new_n543), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT78), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n286), .A2(new_n566), .A3(G244), .A4(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n489), .A2(G33), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n286), .A2(G238), .A3(new_n288), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n565), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n283), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n258), .A2(G45), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n403), .A2(G250), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n281), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AND4_X1   g0375(.A1(KEYINPUT80), .A2(new_n571), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n574), .B1(new_n570), .B2(new_n283), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT80), .B1(new_n577), .B2(new_n573), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n435), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(KEYINPUT80), .A3(new_n573), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n323), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n253), .B1(new_n312), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n209), .A2(new_n442), .A3(new_n214), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT81), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n286), .A2(new_n253), .A3(G68), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n587), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n585), .B1(new_n262), .B2(new_n442), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n256), .B1(new_n254), .B2(new_n424), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n424), .B2(new_n453), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n579), .A2(new_n584), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(G190), .B1(new_n576), .B2(new_n578), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n582), .A2(G200), .A3(new_n583), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n595), .B1(new_n209), .B2(new_n453), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n440), .A2(new_n523), .A3(new_n563), .A4(new_n603), .ZN(G372));
  AOI21_X1  g0404(.A(G179), .B1(new_n582), .B2(new_n583), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n580), .A2(new_n323), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT84), .B1(new_n579), .B2(new_n606), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n596), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT26), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n582), .A2(new_n583), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(G190), .B1(G200), .B2(new_n580), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n600), .B(KEYINPUT85), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n483), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n527), .A2(new_n529), .ZN(new_n619));
  INV_X1    g0419(.A(new_n525), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n532), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT24), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n342), .B1(new_n622), .B2(new_n533), .ZN(new_n623));
  INV_X1    g0423(.A(new_n543), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(new_n541), .A3(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n554), .A2(G169), .B1(G179), .B2(new_n557), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT86), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n499), .A2(new_n512), .A3(new_n507), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n512), .B1(new_n499), .B2(new_n507), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n514), .A2(G179), .A3(new_n479), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n518), .B2(new_n498), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT86), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n544), .A2(new_n559), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n627), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n562), .A2(new_n486), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n618), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n617), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n597), .A2(new_n602), .A3(new_n618), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n608), .B1(new_n605), .B2(new_n607), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n579), .A2(KEYINPUT84), .A3(new_n606), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT87), .B1(new_n643), .B2(new_n596), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  INV_X1    g0445(.A(new_n596), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n645), .B(new_n646), .C1(new_n641), .C2(new_n642), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n440), .B1(new_n638), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n357), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n427), .A2(new_n432), .A3(new_n429), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n432), .B1(new_n427), .B2(new_n429), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n437), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n350), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n354), .A3(new_n412), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n401), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n650), .B1(new_n656), .B2(new_n307), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n649), .A2(new_n657), .ZN(G369));
  NOR2_X1   g0458(.A1(new_n252), .A2(G20), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n258), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G343), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT88), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n499), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n632), .A2(new_n521), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n632), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n670), .A2(KEYINPUT89), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(KEYINPUT89), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n544), .A2(new_n666), .ZN(new_n675));
  INV_X1    g0475(.A(new_n560), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n563), .A2(new_n675), .B1(new_n676), .B2(new_n666), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n627), .A2(new_n634), .ZN(new_n680));
  INV_X1    g0480(.A(new_n666), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n632), .A2(new_n666), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n563), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n226), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n587), .A2(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n232), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n611), .A2(new_n616), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n632), .A2(new_n560), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n636), .A2(new_n694), .A3(new_n483), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n693), .A2(new_n695), .B1(new_n644), .B2(new_n647), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n643), .A2(new_n596), .B1(new_n615), .B2(new_n614), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n483), .A2(new_n612), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n612), .B2(new_n639), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT29), .B(new_n681), .C1(new_n696), .C2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n636), .A2(new_n483), .A3(new_n694), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n611), .A2(new_n645), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n643), .A2(KEYINPUT87), .A3(new_n596), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n703), .A2(new_n697), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n639), .A2(new_n612), .ZN(new_n707));
  INV_X1    g0507(.A(new_n698), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n693), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT90), .A3(KEYINPUT29), .A4(new_n681), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n681), .B1(new_n638), .B2(new_n648), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n702), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n480), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n557), .A2(G179), .A3(new_n514), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n716), .B(new_n717), .C1(new_n576), .C2(new_n578), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(G179), .B1(new_n577), .B2(new_n573), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n480), .A3(new_n506), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(new_n557), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n613), .A2(KEYINPUT30), .A3(new_n716), .A4(new_n717), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n666), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n603), .A2(new_n523), .A3(new_n563), .A4(new_n681), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n715), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n692), .B1(new_n733), .B2(G1), .ZN(G364));
  NAND2_X1  g0534(.A1(new_n659), .A2(G45), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n688), .A2(G1), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT91), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n673), .B(new_n738), .C1(G330), .C2(new_n669), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT92), .Z(new_n740));
  NOR2_X1   g0540(.A1(new_n253), .A2(G190), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n435), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT96), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n253), .A2(new_n295), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n742), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n749), .A2(G77), .B1(G58), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT97), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n435), .A2(new_n405), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n741), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n405), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n221), .A2(new_n757), .B1(new_n759), .B2(new_n209), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n253), .B1(new_n761), .B2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n442), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n758), .A2(new_n741), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n214), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n760), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n754), .A2(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n741), .A2(new_n761), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G159), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n750), .A2(new_n756), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n371), .B(new_n771), .C1(G50), .C2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n755), .A2(new_n766), .A3(new_n767), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n764), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  INV_X1    g0578(.A(G329), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n751), .A2(new_n778), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n749), .B2(G311), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT33), .B(G317), .Z(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n757), .ZN(new_n783));
  INV_X1    g0583(.A(G326), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n371), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n762), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n783), .B(new_n785), .C1(G294), .C2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n781), .B(new_n787), .C1(new_n502), .C2(new_n759), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n775), .B1(new_n777), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n229), .B1(G20), .B2(new_n323), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n738), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n790), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n686), .A2(new_n286), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n232), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT95), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n250), .ZN(new_n799));
  XOR2_X1   g0599(.A(G355), .B(KEYINPUT93), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n286), .A2(new_n226), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(G116), .B2(new_n226), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  OAI21_X1  g0603(.A(new_n795), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n794), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n791), .B(new_n804), .C1(new_n669), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n740), .A2(new_n806), .ZN(G396));
  AND2_X1   g0607(.A1(new_n666), .A2(new_n427), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n653), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n428), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n808), .B1(new_n653), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT99), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT99), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n809), .C1(new_n438), .C2(new_n808), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n712), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n681), .B(new_n816), .C1(new_n638), .C2(new_n648), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(new_n732), .Z(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n738), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n790), .A2(new_n792), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n332), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G137), .A2(new_n773), .B1(new_n752), .B2(G143), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n825), .B1(new_n268), .B2(new_n757), .C1(new_n748), .C2(new_n368), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n286), .B1(new_n768), .B2(new_n828), .C1(new_n202), .C2(new_n759), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G58), .B2(new_n786), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n827), .B(new_n830), .C1(new_n221), .C2(new_n764), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n768), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n764), .A2(new_n209), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G294), .B2(new_n752), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n502), .B2(new_n772), .ZN(new_n836));
  INV_X1    g0636(.A(new_n757), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n763), .B(new_n836), .C1(G283), .C2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n371), .B1(new_n759), .B2(new_n214), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT98), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n749), .A2(new_n489), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n831), .B1(new_n833), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n738), .B1(new_n843), .B2(new_n790), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n824), .B(new_n844), .C1(new_n816), .C2(new_n793), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n822), .A2(new_n845), .ZN(G384));
  OAI211_X1 g0646(.A(G20), .B(new_n230), .C1(new_n446), .C2(KEYINPUT35), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n516), .B(new_n847), .C1(KEYINPUT35), .C2(new_n446), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT36), .Z(new_n849));
  OAI21_X1  g0649(.A(G77), .B1(new_n207), .B2(new_n221), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n850), .A2(new_n232), .B1(G50), .B2(new_n221), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(G1), .A3(new_n252), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT100), .Z(new_n854));
  NAND4_X1  g0654(.A1(new_n398), .A2(new_n400), .A3(new_n410), .A4(new_n411), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n342), .B1(new_n370), .B2(new_n377), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT101), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n386), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT101), .B1(new_n856), .B2(new_n385), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n855), .A2(new_n664), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n395), .B(new_n663), .C1(new_n323), .C2(new_n394), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n387), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n408), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n863), .A2(new_n859), .A3(new_n860), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n408), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n868), .B2(new_n865), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT102), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n855), .A2(new_n387), .A3(new_n664), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n864), .A2(new_n408), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(new_n865), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n862), .A2(new_n869), .A3(KEYINPUT102), .A4(KEYINPUT38), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n872), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n350), .A2(new_n666), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n862), .A2(new_n869), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n873), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n870), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n401), .A2(new_n664), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n349), .A2(new_n666), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n350), .A2(new_n354), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n354), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n349), .B(new_n666), .C1(new_n890), .C2(new_n328), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n434), .A2(new_n437), .A3(new_n681), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n819), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n884), .A2(new_n870), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n887), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n886), .A2(new_n897), .A3(KEYINPUT103), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT103), .B1(new_n886), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n702), .A2(new_n711), .A3(new_n440), .A4(new_n714), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n657), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n900), .B(new_n902), .Z(new_n903));
  NAND3_X1  g0703(.A1(new_n731), .A2(new_n816), .A3(new_n892), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n879), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT40), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n884), .A2(new_n908), .A3(new_n870), .ZN(new_n909));
  INV_X1    g0709(.A(new_n904), .ZN(new_n910));
  NAND2_X1  g0710(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n440), .A2(new_n731), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(G330), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n903), .B(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n659), .A2(new_n258), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n854), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT105), .Z(G367));
  OR2_X1    g0720(.A1(new_n615), .A2(new_n681), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n693), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n704), .B2(new_n705), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT106), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT106), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  XNOR2_X1  g0725(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n666), .A2(new_n456), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n483), .A3(new_n486), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n684), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n483), .B1(new_n929), .B2(new_n560), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT108), .Z(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n666), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT109), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n924), .A2(new_n925), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT43), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n927), .B(new_n934), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT110), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n929), .B1(new_n483), .B2(new_n681), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n679), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n679), .A2(new_n945), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n936), .B(new_n947), .C1(new_n941), .C2(new_n942), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n687), .B(KEYINPUT41), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n684), .B1(new_n678), .B2(new_n683), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n673), .B(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n733), .A2(KEYINPUT112), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT112), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n715), .A2(new_n732), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n952), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n684), .A2(new_n682), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n945), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT44), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(new_n945), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n674), .A2(KEYINPUT111), .A3(new_n678), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n954), .A2(new_n957), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n950), .B1(new_n966), .B2(new_n733), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n735), .A2(G1), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n946), .B(new_n948), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n937), .A2(new_n794), .ZN(new_n970));
  INV_X1    g0770(.A(new_n796), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n795), .B1(new_n226), .B2(new_n424), .C1(new_n242), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n762), .A2(new_n221), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n286), .B1(new_n757), .B2(new_n368), .C1(new_n268), .C2(new_n751), .ZN(new_n974));
  INV_X1    g0774(.A(new_n764), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n973), .B(new_n974), .C1(G77), .C2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(G143), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n772), .A2(new_n977), .B1(new_n759), .B2(new_n207), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n749), .B2(G50), .ZN(new_n979));
  INV_X1    g0779(.A(G137), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n976), .B(new_n979), .C1(new_n980), .C2(new_n768), .ZN(new_n981));
  INV_X1    g0781(.A(new_n759), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT46), .B1(new_n982), .B2(new_n489), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(KEYINPUT46), .A3(G116), .ZN(new_n984));
  INV_X1    g0784(.A(G294), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(new_n985), .B2(new_n757), .C1(new_n502), .C2(new_n751), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n983), .B(new_n986), .C1(G107), .C2(new_n786), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n371), .B1(new_n768), .B2(new_n988), .C1(new_n442), .C2(new_n764), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT113), .Z(new_n990));
  OAI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(new_n776), .C2(new_n748), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n772), .A2(new_n832), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n738), .B1(new_n994), .B2(new_n790), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n970), .A2(new_n972), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n969), .A2(new_n996), .ZN(G387));
  NAND2_X1  g0797(.A1(new_n954), .A2(new_n957), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n687), .C1(new_n733), .C2(new_n953), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n975), .A2(new_n489), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G322), .A2(new_n773), .B1(new_n837), .B2(G311), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n988), .B2(new_n751), .C1(new_n748), .C2(new_n502), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT48), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n776), .B2(new_n762), .C1(new_n985), .C2(new_n759), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n286), .B(new_n1000), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n1004), .C1(new_n784), .C2(new_n768), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n772), .A2(new_n368), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n982), .A2(G77), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n202), .B2(new_n751), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n749), .B2(G68), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n286), .B1(new_n764), .B2(new_n442), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n424), .A2(new_n762), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n383), .C2(new_n837), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1011), .B(new_n1014), .C1(new_n268), .C2(new_n768), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1007), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n738), .B1(new_n1016), .B2(new_n790), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n678), .B2(new_n805), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n238), .A2(G45), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n263), .A2(G50), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n221), .A2(new_n332), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n689), .ZN(new_n1023));
  AOI211_X1 g0823(.A(G45), .B(new_n1022), .C1(new_n1023), .C2(KEYINPUT114), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(KEYINPUT114), .C2(new_n1023), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1019), .A2(new_n796), .A3(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(G107), .B2(new_n226), .C1(new_n689), .C2(new_n801), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1018), .B1(new_n795), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n953), .B2(new_n968), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n999), .A2(new_n1029), .ZN(G393));
  XOR2_X1   g0830(.A(new_n963), .B(new_n679), .Z(new_n1031));
  INV_X1    g0831(.A(new_n968), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n837), .A2(G50), .B1(new_n769), .B2(G143), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n221), .B2(new_n759), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n762), .A2(new_n332), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1035), .A2(new_n371), .A3(new_n834), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT51), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n772), .A2(new_n268), .B1(new_n751), .B2(new_n368), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n749), .A2(new_n383), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n757), .A2(new_n502), .B1(new_n768), .B2(new_n778), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n765), .B(new_n1042), .C1(G283), .C2(new_n982), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n749), .A2(G294), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n772), .A2(new_n988), .B1(new_n751), .B2(new_n832), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n286), .B1(new_n786), .B2(new_n489), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n790), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n246), .A2(new_n796), .B1(G97), .B2(new_n686), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n795), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n737), .A3(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n945), .A2(new_n794), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n688), .B1(new_n998), .B2(new_n1031), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT116), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n966), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1058), .B1(new_n1057), .B2(new_n966), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1033), .B(new_n1056), .C1(new_n1060), .C2(new_n1061), .ZN(G390));
  OAI221_X1 g0862(.A(new_n371), .B1(new_n759), .B2(new_n209), .C1(new_n776), .C2(new_n772), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1036), .B(new_n1063), .C1(G68), .C2(new_n975), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n751), .A2(new_n516), .B1(new_n757), .B2(new_n214), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n749), .B2(G97), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(new_n985), .C2(new_n768), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G50), .A2(new_n975), .B1(new_n769), .B2(G125), .ZN(new_n1068));
  INV_X1    g0868(.A(G128), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n772), .C1(new_n980), .C2(new_n757), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n371), .B(new_n1070), .C1(G159), .C2(new_n786), .ZN(new_n1071));
  XOR2_X1   g0871(.A(KEYINPUT54), .B(G143), .Z(new_n1072));
  NAND2_X1  g0872(.A1(new_n749), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(new_n828), .C2(new_n751), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n982), .A2(G150), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT53), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1067), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n738), .B1(new_n1077), .B2(new_n790), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n881), .A2(new_n885), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n793), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n263), .B2(new_n823), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n731), .A2(new_n816), .A3(new_n892), .A4(G330), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n819), .A2(new_n894), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n892), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n882), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1085), .A2(new_n1086), .B1(new_n881), .B2(new_n885), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n681), .B(new_n816), .C1(new_n696), .C2(new_n699), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n893), .B1(new_n1088), .B2(new_n894), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n879), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n882), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1083), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1088), .A2(new_n894), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1086), .B(new_n879), .C1(new_n1093), .C2(new_n893), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n895), .A2(new_n882), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1082), .C1(new_n1079), .C2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1096), .A3(new_n968), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT117), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT117), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1092), .A2(new_n1096), .A3(new_n1099), .A4(new_n968), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1081), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n731), .A2(new_n816), .A3(G330), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n893), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1082), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1084), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1093), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n1105), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n440), .A2(G330), .A3(new_n731), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1108), .A2(new_n657), .A3(new_n901), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1102), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n901), .A2(new_n657), .A3(new_n1109), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1104), .A2(new_n1082), .B1(new_n819), .B2(new_n894), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1105), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n1093), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1111), .A2(new_n687), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1101), .A2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(new_n1112), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT119), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n304), .A2(new_n306), .A3(new_n357), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT55), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT55), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n304), .A2(new_n306), .A3(new_n1127), .A4(new_n357), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n272), .A2(new_n664), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1132), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n1123), .A3(new_n1130), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n908), .B1(new_n879), .B2(new_n905), .ZN(new_n1138));
  OAI211_X1 g0938(.A(G330), .B(new_n1136), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(G330), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n900), .A2(new_n1122), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n886), .A2(new_n897), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT103), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n886), .A2(new_n897), .A3(KEYINPUT103), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1122), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1142), .A2(new_n1139), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1121), .A2(new_n1143), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1136), .B1(new_n913), .B2(G330), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1139), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1154), .A2(new_n1155), .B1(new_n898), .B2(new_n899), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1146), .A2(new_n1142), .A3(new_n1147), .A4(new_n1139), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n1121), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT120), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT57), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1153), .A2(new_n1159), .A3(new_n1163), .A4(new_n687), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1143), .A2(new_n968), .A3(new_n1150), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n823), .A2(new_n202), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n748), .A2(new_n980), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G125), .A2(new_n773), .B1(new_n752), .B2(G128), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n828), .B2(new_n757), .C1(new_n268), .C2(new_n762), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n982), .C2(new_n1072), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT59), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G41), .B1(new_n769), .B2(G124), .ZN(new_n1172));
  AOI21_X1  g0972(.A(G33), .B1(new_n975), .B2(G159), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n202), .B1(new_n309), .B2(G41), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1009), .B1(new_n442), .B2(new_n757), .C1(new_n214), .C2(new_n751), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1176), .A2(G41), .A3(new_n286), .A4(new_n973), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n764), .A2(new_n207), .B1(new_n768), .B2(new_n776), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n749), .B2(new_n423), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n516), .C2(new_n772), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT58), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1174), .A2(new_n1175), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n738), .B1(new_n1182), .B2(new_n790), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1166), .B(new_n1183), .C1(new_n1136), .C2(new_n793), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1165), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1164), .A2(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1110), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n949), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT121), .Z(new_n1191));
  AOI22_X1  g0991(.A1(new_n749), .A2(G107), .B1(new_n489), .B2(new_n837), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n985), .B2(new_n772), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT123), .Z(new_n1194));
  AOI22_X1  g0994(.A1(new_n982), .A2(G97), .B1(new_n769), .B2(G303), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n332), .B2(new_n764), .C1(new_n776), .C2(new_n751), .ZN(new_n1196));
  OR4_X1    g0996(.A1(new_n286), .A2(new_n1194), .A3(new_n1013), .A4(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n772), .A2(new_n828), .B1(new_n751), .B2(new_n980), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n749), .B2(G150), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n837), .A2(new_n1072), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n982), .A2(G159), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n286), .B1(new_n768), .B2(new_n1069), .C1(new_n207), .C2(new_n764), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G50), .B2(new_n786), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1197), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n738), .B1(new_n1205), .B2(new_n790), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n893), .A2(KEYINPUT122), .A3(new_n792), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n823), .A2(new_n221), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT122), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n892), .B2(new_n793), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1108), .B2(new_n968), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1191), .A2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT124), .ZN(G381));
  OR2_X1    g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(G381), .A2(G384), .A3(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G375), .A2(G378), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1057), .A2(new_n966), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT116), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1220), .A2(new_n1059), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1221), .A2(new_n996), .A3(new_n969), .A4(new_n1033), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1217), .A2(new_n1218), .A3(new_n1223), .ZN(G407));
  AND2_X1   g1024(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n688), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1185), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  INV_X1    g1030(.A(G384), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT60), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1110), .B2(new_n1188), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n688), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1213), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1231), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1234), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n687), .B(new_n1238), .C1(new_n1189), .C2(new_n1232), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(G384), .A3(new_n1213), .ZN(new_n1240));
  INV_X1    g1040(.A(G213), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(G343), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(G2897), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1237), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1228), .B1(new_n1164), .B2(new_n1186), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1156), .A2(new_n1157), .A3(new_n968), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(KEYINPUT125), .A3(new_n1184), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1121), .A2(new_n1143), .A3(new_n949), .A4(new_n1150), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1118), .A4(new_n1101), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1248), .A2(new_n1184), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT125), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n1251), .A2(new_n1253), .B1(new_n1241), .B2(G343), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1246), .B1(new_n1247), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT63), .ZN(new_n1256));
  AND4_X1   g1056(.A1(new_n1118), .A2(new_n1249), .A3(new_n1250), .A4(new_n1101), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1252), .A2(KEYINPUT125), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1242), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1216), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(G390), .B2(G387), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1221), .A2(new_n1033), .B1(new_n996), .B2(new_n969), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1265), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G390), .A2(G387), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1222), .A2(new_n1270), .A3(new_n1266), .A4(new_n1264), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1247), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1274), .A2(KEYINPUT63), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1262), .A2(new_n1273), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1274), .A2(new_n1278), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT127), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1255), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1255), .B2(new_n1282), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1280), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1276), .B1(new_n1285), .B2(new_n1273), .ZN(G405));
  NOR2_X1   g1086(.A1(new_n1218), .A2(new_n1247), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1272), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1269), .B(new_n1271), .C1(new_n1218), .C2(new_n1247), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1288), .A2(new_n1260), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1260), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


