//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n464), .A2(new_n467), .A3(G137), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n468), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(G160));
  AND3_X1   g052(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n472), .B2(G112), .ZN(new_n482));
  OAI22_X1  g057(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n472), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n483), .B1(G136), .B2(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(new_n472), .B2(G114), .ZN(new_n487));
  NOR2_X1   g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT67), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n488), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n473), .A2(new_n468), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n472), .A2(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n472), .A2(KEYINPUT4), .A3(G138), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n502), .A2(new_n468), .A3(new_n464), .A4(new_n467), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n495), .A2(new_n497), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  XOR2_X1   g080(.A(KEYINPUT5), .B(G543), .Z(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT68), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n508), .A2(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n506), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G651), .B1(G50), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  AND2_X1   g100(.A1(new_n515), .A2(G63), .ZN(new_n526));
  AND3_X1   g101(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(G651), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT69), .B(G51), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n523), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n517), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n517), .A2(G90), .B1(G52), .B2(new_n523), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT70), .ZN(new_n539));
  INV_X1    g114(.A(G77), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI221_X1 g116(.A(KEYINPUT70), .B1(new_n540), .B2(new_n522), .C1(new_n506), .C2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(G651), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n537), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n517), .A2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n506), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G651), .B1(G43), .B2(new_n523), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  AOI22_X1  g133(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n507), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n512), .A2(new_n516), .A3(G91), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n508), .A2(new_n510), .A3(G53), .A4(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(G299));
  NAND2_X1  g139(.A1(new_n537), .A2(new_n543), .ZN(G301));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n535), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT73), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G286));
  NAND2_X1  g145(.A1(new_n518), .A2(new_n524), .ZN(G303));
  OR2_X1    g146(.A1(new_n515), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n523), .B2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n512), .A2(new_n516), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n506), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(new_n580), .A3(G651), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT74), .B1(new_n582), .B2(new_n507), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n523), .A2(G48), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n512), .A2(new_n516), .A3(G86), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n517), .A2(G85), .B1(G47), .B2(new_n523), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n506), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n507), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(new_n591), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n588), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n513), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G54), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n597), .A2(new_n507), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n574), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n602), .A2(new_n603), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n596), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n596), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n569), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(KEYINPUT77), .B1(new_n611), .B2(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(KEYINPUT77), .B2(new_n613), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(KEYINPUT77), .B2(new_n613), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n550), .A2(new_n611), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n608), .A2(new_n617), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n621), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g198(.A(KEYINPUT3), .B(G2104), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n466), .A2(G2105), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n630), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n479), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(G135), .B2(new_n485), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT80), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT81), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(KEYINPUT82), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n659), .A2(new_n662), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n659), .A2(new_n662), .ZN(new_n669));
  INV_X1    g244(.A(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(new_n661), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n664), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT83), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  AOI211_X1 g259(.A(new_n682), .B(new_n684), .C1(new_n677), .C2(new_n681), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT84), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(G229));
  INV_X1    g270(.A(KEYINPUT24), .ZN(new_n696));
  INV_X1    g271(.A(G34), .ZN(new_n697));
  AOI21_X1  g272(.A(G29), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(G160), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G2084), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(G33), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n624), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(new_n472), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT91), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT25), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n485), .B2(G139), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(new_n700), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n702), .B1(new_n711), .B2(G2072), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G2072), .B2(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT26), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n716), .A2(new_n717), .B1(G105), .B2(new_n625), .ZN(new_n718));
  INV_X1    g293(.A(G141), .ZN(new_n719));
  INV_X1    g294(.A(G129), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n718), .B1(new_n484), .B2(new_n719), .C1(new_n720), .C2(new_n479), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT93), .ZN(new_n728));
  INV_X1    g303(.A(G32), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n700), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT27), .B(G1996), .Z(new_n731));
  OAI21_X1  g306(.A(new_n713), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT94), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G4), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n608), .B2(new_n734), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT89), .B(G1348), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(G5), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G171), .B2(new_n734), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT96), .B(G1961), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n700), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n700), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT29), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n742), .B1(G2084), .B2(new_n701), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n738), .B(new_n748), .C1(new_n747), .C2(new_n746), .ZN(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n734), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n734), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G1341), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n551), .A2(new_n734), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n734), .B2(G19), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n754), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n751), .A2(new_n752), .ZN(new_n759));
  NOR2_X1   g334(.A1(G164), .A2(new_n700), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G27), .B2(new_n700), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT97), .B(G2078), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT95), .B(G28), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT31), .B(G11), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n637), .B2(G29), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n761), .A2(new_n762), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n759), .A2(new_n763), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n700), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n485), .A2(G140), .ZN(new_n775));
  INV_X1    g350(.A(G104), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n776), .A2(new_n472), .A3(KEYINPUT90), .ZN(new_n777));
  AOI21_X1  g352(.A(KEYINPUT90), .B1(new_n776), .B2(new_n472), .ZN(new_n778));
  OAI221_X1 g353(.A(G2104), .B1(G116), .B2(new_n472), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G128), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n479), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n700), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2067), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n734), .A2(G20), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT23), .Z(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n758), .A2(new_n772), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n730), .A2(new_n731), .ZN(new_n792));
  AND3_X1   g367(.A1(new_n749), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n733), .A2(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  INV_X1    g371(.A(G1981), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G23), .B(G288), .S(G16), .Z(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT33), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G1976), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(G1976), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n734), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n734), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT88), .B(G1971), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n798), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(G16), .Z(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1986), .Z(new_n812));
  INV_X1    g387(.A(KEYINPUT87), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n700), .A2(G25), .ZN(new_n816));
  INV_X1    g391(.A(G95), .ZN(new_n817));
  AND3_X1   g392(.A1(new_n817), .A2(new_n472), .A3(KEYINPUT86), .ZN(new_n818));
  AOI21_X1  g393(.A(KEYINPUT86), .B1(new_n817), .B2(new_n472), .ZN(new_n819));
  OAI221_X1 g394(.A(G2104), .B1(G107), .B2(new_n472), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G119), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n479), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G131), .B2(new_n485), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n816), .B1(new_n823), .B2(new_n700), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  XOR2_X1   g400(.A(new_n824), .B(new_n825), .Z(new_n826));
  NOR3_X1   g401(.A1(new_n814), .A2(new_n815), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n809), .A2(new_n810), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n794), .B1(new_n829), .B2(new_n830), .ZN(G311));
  XNOR2_X1  g406(.A(new_n828), .B(KEYINPUT36), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n832), .A2(new_n733), .A3(new_n793), .ZN(G150));
  AOI22_X1  g408(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n507), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT99), .B(G55), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n523), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n574), .A2(new_n840), .B1(new_n835), .B2(KEYINPUT98), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n545), .A2(KEYINPUT100), .A3(new_n549), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT100), .B1(new_n545), .B2(new_n549), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n551), .A2(new_n842), .A3(KEYINPUT100), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n600), .B(new_n601), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n604), .A2(new_n607), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n617), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n849), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(G860), .B1(new_n839), .B2(new_n841), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n725), .B(new_n783), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n823), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n504), .A2(KEYINPUT101), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n478), .A2(new_n502), .B1(new_n489), .B2(new_n494), .ZN(new_n864));
  AND4_X1   g439(.A1(new_n468), .A2(new_n464), .A3(new_n467), .A4(new_n496), .ZN(new_n865));
  INV_X1    g440(.A(new_n500), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT4), .B1(new_n624), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n710), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n875));
  OAI22_X1  g450(.A1(new_n479), .A2(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(G142), .B2(new_n485), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n627), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n872), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n862), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n637), .B(G160), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(G162), .Z(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n882), .B2(new_n880), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g460(.A(new_n848), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n620), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  INV_X1    g463(.A(G299), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n852), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n608), .A2(KEYINPUT102), .A3(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n608), .B2(G299), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n852), .A2(KEYINPUT103), .A3(new_n889), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n892), .A2(new_n900), .A3(new_n894), .A4(new_n895), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n898), .B1(new_n902), .B2(new_n887), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  XOR2_X1   g479(.A(G290), .B(G305), .Z(new_n905));
  XNOR2_X1  g480(.A(G166), .B(G288), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n898), .B(new_n909), .C1(new_n902), .C2(new_n887), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n904), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n908), .B1(new_n904), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(G868), .B2(new_n842), .ZN(G295));
  OAI21_X1  g489(.A(new_n913), .B1(G868), .B2(new_n842), .ZN(G331));
  AOI21_X1  g490(.A(G301), .B1(new_n567), .B2(new_n568), .ZN(new_n916));
  NAND2_X1  g491(.A1(G301), .A2(new_n535), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n846), .A2(new_n847), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n568), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT73), .B1(new_n533), .B2(new_n534), .ZN(new_n921));
  OAI21_X1  g496(.A(G171), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n844), .A2(new_n845), .ZN(new_n923));
  INV_X1    g498(.A(new_n845), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n843), .A3(new_n842), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .A4(new_n917), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n899), .A2(new_n901), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n916), .A2(new_n918), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n848), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(KEYINPUT105), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n896), .A4(new_n919), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n907), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n907), .B1(new_n928), .B2(new_n933), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n931), .A2(new_n932), .A3(new_n919), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n899), .A3(new_n901), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n897), .B2(new_n927), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n919), .A4(new_n926), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n936), .B1(new_n908), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n940), .B(KEYINPUT44), .C1(new_n941), .C2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n934), .A2(new_n935), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n908), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n937), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT107), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n957), .B(KEYINPUT44), .C1(new_n952), .C2(new_n953), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n949), .B1(new_n956), .B2(new_n958), .ZN(G397));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  NAND4_X1  g535(.A1(G160), .A2(new_n504), .A3(G40), .A4(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1976), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n961), .B(G8), .C1(new_n962), .C2(G288), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT52), .ZN(new_n964));
  NAND2_X1  g539(.A1(G288), .A2(new_n962), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n964), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n581), .A2(new_n583), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n586), .A2(new_n585), .ZN(new_n971));
  OAI21_X1  g546(.A(G1981), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n584), .A2(new_n797), .A3(new_n585), .A4(new_n586), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n961), .A2(G8), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n974), .B2(new_n975), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n968), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n980));
  AND2_X1   g555(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n981));
  OAI211_X1 g556(.A(G303), .B(G8), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  NOR2_X1   g558(.A1(G166), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n984), .B2(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n469), .A2(new_n470), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n472), .ZN(new_n987));
  INV_X1    g562(.A(new_n476), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G40), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n466), .B1(new_n491), .B2(G2105), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n493), .B1(new_n991), .B2(new_n490), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n487), .A2(KEYINPUT67), .A3(new_n488), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n503), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n501), .A2(new_n497), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n960), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n989), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT108), .B(G1384), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n863), .A2(new_n870), .A3(KEYINPUT45), .A4(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G1971), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(G40), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n471), .A2(new_n1002), .A3(new_n476), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n504), .A2(new_n1004), .A3(new_n960), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G2090), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n985), .B(G8), .C1(new_n1000), .C2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1007), .B2(new_n1000), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n984), .A2(new_n981), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n982), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n979), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G2084), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1001), .A2(new_n1013), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n864), .B2(new_n868), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT45), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1966), .B1(new_n997), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(G8), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G286), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1011), .A2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g599(.A(G8), .B1(new_n1000), .B2(new_n1007), .C1(new_n985), .C2(new_n1023), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1025), .A2(new_n979), .A3(KEYINPUT63), .A4(new_n1020), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1022), .A2(KEYINPUT63), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n973), .B(KEYINPUT113), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n976), .A2(new_n978), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(G1976), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n1030), .B(KEYINPUT114), .Z(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n977), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1008), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1032), .A2(new_n1033), .B1(new_n1034), .B2(new_n979), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT126), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT123), .B1(new_n1019), .B2(KEYINPUT51), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n983), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1003), .B1(new_n1016), .B2(KEYINPUT45), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n996), .A2(new_n990), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n752), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n983), .B1(new_n1043), .B2(new_n1014), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1043), .A2(new_n1014), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(G8), .C1(new_n1049), .C2(new_n535), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1039), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1047), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1052), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1039), .B1(new_n1019), .B2(KEYINPUT123), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1045), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2078), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n997), .A2(new_n999), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  INV_X1    g637(.A(G1961), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1061), .A2(new_n1062), .B1(new_n1063), .B2(new_n1006), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(G2078), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n997), .A2(new_n1065), .A3(new_n1017), .ZN(new_n1066));
  AOI21_X1  g641(.A(G301), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n979), .A2(new_n1011), .A3(new_n1067), .A4(new_n1008), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1053), .A2(new_n1059), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT125), .B1(new_n1071), .B2(KEYINPUT62), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1037), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1052), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1058), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1068), .B1(new_n1075), .B2(new_n1058), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(KEYINPUT126), .A4(new_n1053), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1036), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n863), .A2(new_n870), .A3(new_n998), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1080), .A2(new_n990), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n999), .A2(new_n1003), .A3(new_n1065), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1064), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1084), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT124), .B1(new_n1084), .B2(G171), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1067), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(G171), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1064), .A2(G301), .A3(new_n1066), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(KEYINPUT54), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1075), .A2(new_n1012), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1090), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1006), .A2(new_n789), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n997), .A2(new_n999), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n560), .A2(new_n561), .A3(new_n563), .A4(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n961), .ZN(new_n1104));
  INV_X1    g679(.A(G2067), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  INV_X1    g682(.A(G1348), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1106), .A2(new_n1107), .B1(new_n1006), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(KEYINPUT116), .A3(new_n1105), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n608), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1103), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n1110), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n608), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n852), .A4(new_n1110), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1116), .A2(new_n1113), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1102), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1117), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1129));
  INV_X1    g704(.A(G1996), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n997), .A2(new_n999), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT118), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  AND3_X1   g708(.A1(new_n961), .A2(KEYINPUT119), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT119), .B1(new_n961), .B2(new_n1133), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n997), .A2(new_n999), .A3(new_n1137), .A4(new_n1130), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1140));
  AND3_X1   g715(.A1(new_n1139), .A2(new_n551), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1140), .B1(new_n1139), .B2(new_n551), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1128), .B(new_n1129), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1124), .B1(new_n1143), .B2(KEYINPUT121), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1127), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1102), .A2(new_n1145), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1146), .B(new_n1147), .C1(new_n1142), .C2(new_n1141), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1118), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1095), .B1(new_n1149), .B2(KEYINPUT122), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n1151), .B(new_n1118), .C1(new_n1144), .C2(new_n1148), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1079), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1081), .A2(new_n1003), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n823), .A2(new_n825), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n823), .A2(new_n825), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n782), .B(new_n1105), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n726), .B2(new_n1130), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1154), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1154), .A2(new_n1130), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT110), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1161), .B1(new_n1163), .B2(new_n725), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT109), .B1(G290), .B2(G1986), .ZN(new_n1165));
  NAND2_X1  g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1158), .B(new_n1164), .C1(new_n1154), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1153), .A2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1155), .A2(G1986), .A3(G290), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(KEYINPUT48), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1170), .A2(KEYINPUT48), .ZN(new_n1172));
  NOR4_X1   g747(.A1(new_n1164), .A2(new_n1158), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1164), .A2(new_n1157), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n783), .A2(new_n1105), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1155), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1155), .B1(new_n726), .B2(new_n1159), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1163), .A2(KEYINPUT46), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1163), .A2(KEYINPUT46), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT47), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1173), .B(new_n1176), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1169), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g760(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n693), .A2(new_n694), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n1188), .A2(new_n884), .A3(new_n954), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


