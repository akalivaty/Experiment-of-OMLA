//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0006(.A(new_n201), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n213), .B1(new_n220), .B2(KEYINPUT0), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n218), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G68), .ZN(new_n230));
  INV_X1    g0030(.A(G238), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n215), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n221), .B(new_n234), .C1(KEYINPUT0), .C2(new_n220), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n230), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n247), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n210), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(KEYINPUT67), .A3(new_n210), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(G58), .B(G68), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n260), .A2(G20), .B1(G159), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(G20), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT7), .ZN(new_n268));
  OAI21_X1  g0068(.A(G68), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n264), .A2(new_n266), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT75), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n270), .A2(new_n274), .A3(new_n211), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT16), .B(new_n262), .C1(new_n269), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n260), .A2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n261), .A2(G159), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n274), .B1(new_n280), .B2(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(new_n283), .B2(G68), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n259), .B(new_n276), .C1(new_n284), .C2(KEYINPUT16), .ZN(new_n285));
  XOR2_X1   g0085(.A(KEYINPUT8), .B(G58), .Z(new_n286));
  INV_X1    g0086(.A(G1), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G13), .A3(G20), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n259), .B1(new_n287), .B2(G20), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n286), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G87), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT76), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n264), .A2(new_n266), .A3(G223), .A4(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n264), .A2(new_n266), .A3(G226), .A4(G1698), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  OAI211_X1 g0100(.A(G1), .B(G13), .C1(new_n263), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n287), .B1(G41), .B2(G45), .ZN(new_n304));
  INV_X1    g0104(.A(G274), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(KEYINPUT66), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT66), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n287), .C1(G41), .C2(G45), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(new_n229), .ZN(new_n312));
  OAI21_X1  g0112(.A(G169), .B1(new_n303), .B2(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n308), .A2(new_n301), .A3(new_n310), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n306), .B1(new_n314), .B2(G232), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n299), .A2(new_n302), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G179), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n292), .A2(KEYINPUT18), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT77), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n285), .A2(new_n291), .B1(new_n313), .B2(new_n317), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT77), .A3(KEYINPUT18), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n292), .A2(new_n318), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT18), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(G200), .B1(new_n303), .B2(new_n312), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n315), .A2(G190), .A3(new_n316), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n285), .A2(new_n328), .A3(new_n291), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT17), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n303), .A2(new_n332), .A3(new_n312), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n315), .B2(new_n316), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT17), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n291), .A4(new_n285), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n280), .A2(G226), .A3(new_n296), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n280), .A2(G1698), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n342), .B1(new_n263), .B2(new_n225), .C1(new_n343), .C2(new_n229), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n302), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n306), .B1(new_n314), .B2(G238), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n345), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g0150(.A(G200), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n259), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(G68), .C1(G1), .C2(new_n211), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT73), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n263), .A2(G20), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G77), .B1(G20), .B2(new_n230), .ZN(new_n356));
  INV_X1    g0156(.A(new_n261), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n202), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT11), .B1(new_n358), .B2(new_n259), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT74), .B1(new_n288), .B2(G68), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT12), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n354), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n345), .A2(new_n347), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT13), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(G190), .A3(new_n348), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n351), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G169), .B1(new_n349), .B2(new_n350), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT14), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT14), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(G169), .C1(new_n349), .C2(new_n350), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n349), .A2(new_n350), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G179), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n365), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n369), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n270), .A2(G107), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n280), .A2(new_n296), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n379), .B1(new_n380), .B2(new_n229), .C1(new_n231), .C2(new_n343), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n302), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n307), .B1(new_n311), .B2(new_n224), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n383), .A2(KEYINPUT69), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(KEYINPUT69), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n290), .A2(G77), .ZN(new_n389));
  INV_X1    g0189(.A(new_n286), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n390), .A2(new_n357), .B1(new_n211), .B2(new_n223), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n211), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n259), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n288), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n223), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT70), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n389), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n388), .B(new_n399), .C1(G179), .C2(new_n386), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n386), .B2(G200), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n332), .B2(new_n386), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n341), .A2(new_n378), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n280), .A2(G222), .A3(new_n296), .ZN(new_n404));
  INV_X1    g0204(.A(G223), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n404), .B1(new_n223), .B2(new_n280), .C1(new_n343), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n302), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n306), .B1(new_n314), .B2(G226), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G200), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT10), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(G190), .A3(new_n408), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n203), .A2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT68), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n286), .A2(new_n355), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n203), .A2(KEYINPUT68), .A3(G20), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n261), .A2(G150), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n259), .B1(new_n202), .B2(new_n396), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n290), .A2(G50), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n421), .A2(KEYINPUT9), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT9), .B1(new_n421), .B2(new_n422), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT71), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n422), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT9), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT71), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n421), .A2(KEYINPUT9), .A3(new_n422), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n413), .A2(new_n425), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT72), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n413), .A2(new_n425), .A3(new_n431), .A4(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n428), .A2(new_n430), .A3(new_n410), .A4(new_n412), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n433), .A2(new_n435), .B1(KEYINPUT10), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n409), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n426), .C1(G169), .C2(new_n438), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n403), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT21), .ZN(new_n444));
  INV_X1    g0244(.A(G303), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n343), .A2(new_n219), .B1(new_n445), .B2(new_n280), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n380), .A2(new_n218), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n302), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n287), .B(G45), .C1(new_n300), .C2(KEYINPUT5), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n300), .A2(KEYINPUT5), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G274), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n301), .B(G270), .C1(new_n449), .C2(new_n450), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n452), .A2(KEYINPUT79), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT79), .B1(new_n452), .B2(new_n453), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n448), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G169), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n254), .A2(new_n210), .B1(G20), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n211), .C1(G33), .C2(new_n225), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n459), .A2(KEYINPUT20), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n396), .A2(new_n458), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n288), .B1(G1), .B2(new_n263), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n352), .A2(G116), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n259), .A2(new_n469), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT80), .A3(G116), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n468), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n444), .B1(new_n457), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT81), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT81), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n444), .C1(new_n457), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n264), .A2(new_n266), .A3(new_n211), .A4(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n280), .A2(new_n484), .A3(new_n211), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(G20), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT82), .B1(new_n211), .B2(G107), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT23), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT23), .ZN(new_n491));
  OAI211_X1 g0291(.A(KEYINPUT82), .B(new_n491), .C1(new_n211), .C2(G107), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT83), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT24), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n486), .A2(new_n497), .A3(new_n493), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n494), .B2(KEYINPUT24), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n259), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n288), .A2(G107), .ZN(new_n502));
  OR2_X1    g0302(.A1(new_n502), .A2(KEYINPUT25), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT84), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n502), .B2(KEYINPUT25), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n474), .A2(G107), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(new_n505), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n449), .A2(new_n450), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(G264), .A4(new_n301), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n301), .B(G264), .C1(new_n449), .C2(new_n450), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n280), .A2(G250), .A3(new_n296), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n280), .A2(G257), .A3(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G294), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n514), .A2(new_n516), .B1(new_n520), .B2(new_n302), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G179), .A3(new_n452), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n387), .B1(new_n521), .B2(new_n452), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT86), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n524), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT86), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(new_n522), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n511), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n448), .B(G179), .C1(new_n454), .C2(new_n455), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n457), .B2(new_n444), .ZN(new_n531));
  INV_X1    g0331(.A(new_n476), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n481), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(G200), .B1(new_n521), .B2(new_n452), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n521), .A2(new_n452), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n535), .A2(KEYINPUT87), .B1(new_n536), .B2(G190), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(KEYINPUT87), .A3(new_n334), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n501), .B(new_n510), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT6), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n540), .A2(new_n225), .A3(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(G97), .B(G107), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n543), .A2(new_n211), .B1(new_n223), .B2(new_n357), .ZN(new_n544));
  INV_X1    g0344(.A(G107), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n281), .B2(new_n282), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n259), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n288), .A2(G97), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n474), .B2(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n280), .A2(G244), .A3(new_n296), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n553), .A2(new_n460), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n302), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n451), .A2(new_n302), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(G257), .B1(G274), .B2(new_n451), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n550), .B1(G200), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n452), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n302), .B2(new_n556), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n560), .A2(new_n387), .B1(new_n547), .B2(new_n549), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n439), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n561), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n569));
  NAND2_X1  g0369(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n225), .B2(new_n393), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n280), .A2(new_n211), .A3(G68), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(G33), .A3(G97), .A4(new_n570), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(new_n211), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n259), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n474), .A2(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n392), .A2(new_n396), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G45), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n301), .B(G250), .C1(G1), .C2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(G1), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G274), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n280), .A2(G244), .A3(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n587), .B(new_n487), .C1(new_n380), .C2(new_n231), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n586), .B1(new_n588), .B2(new_n302), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G190), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n581), .B(new_n590), .C1(new_n334), .C2(new_n589), .ZN(new_n591));
  INV_X1    g0391(.A(new_n474), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n578), .B(new_n580), .C1(new_n592), .C2(new_n392), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n589), .A2(new_n439), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(G169), .C2(new_n589), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n456), .A2(G200), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n598), .B(new_n476), .C1(new_n332), .C2(new_n456), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n539), .A2(new_n568), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n534), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n443), .A2(new_n601), .ZN(G372));
  AND2_X1   g0402(.A1(new_n568), .A2(new_n597), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n481), .A2(new_n533), .ZN(new_n604));
  INV_X1    g0404(.A(new_n511), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n523), .A2(new_n524), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n603), .B(new_n539), .C1(new_n604), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n566), .A2(new_n567), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n596), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g0410(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT26), .B1(new_n596), .B2(new_n609), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n612), .A2(new_n595), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n443), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g0416(.A(new_n616), .B(KEYINPUT89), .Z(new_n617));
  AOI22_X1  g0417(.A1(new_n370), .A2(KEYINPUT14), .B1(new_n374), .B2(G179), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n365), .B1(new_n618), .B2(new_n373), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n369), .A2(new_n400), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n339), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n326), .A2(new_n319), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n433), .A2(new_n435), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n436), .A2(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n442), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT90), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n617), .A2(new_n628), .ZN(G369));
  AND2_X1   g0429(.A1(new_n211), .A2(G13), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n287), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G213), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G343), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n476), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n604), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n599), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(KEYINPUT91), .A3(G330), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  INV_X1    g0443(.A(G330), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n529), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n636), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n529), .B(new_n539), .C1(new_n605), .C2(new_n637), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n604), .A2(new_n637), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n607), .A2(new_n637), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(G399));
  NOR2_X1   g0457(.A1(new_n217), .A2(G41), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n575), .A2(new_n458), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n658), .A2(new_n287), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n209), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g0461(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n560), .A2(new_n536), .ZN(new_n664));
  INV_X1    g0464(.A(new_n589), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n456), .A2(new_n665), .A3(new_n439), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT93), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n456), .A2(new_n665), .A3(new_n668), .A4(new_n439), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n664), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n530), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n521), .A2(new_n589), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT30), .A4(new_n564), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n557), .A2(new_n521), .A3(new_n589), .A4(new_n559), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n530), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(KEYINPUT31), .B(new_n636), .C1(new_n670), .C2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n601), .B2(new_n637), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n636), .B1(new_n670), .B2(new_n677), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n644), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n534), .A2(new_n539), .A3(new_n603), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n610), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n687), .B(new_n595), .C1(new_n610), .C2(new_n611), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n637), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n636), .B1(new_n608), .B2(new_n614), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n684), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n663), .B1(new_n694), .B2(G1), .ZN(G364));
  INV_X1    g0495(.A(new_n646), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n287), .B1(new_n630), .B2(G45), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n658), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n696), .B(new_n700), .C1(G330), .C2(new_n641), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n210), .B1(G20), .B2(new_n387), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G179), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G190), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n225), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n211), .A2(G190), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n704), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G159), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT32), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n211), .A2(new_n439), .A3(new_n334), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n332), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n708), .B(new_n713), .C1(G50), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n439), .A2(G200), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT95), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n211), .A2(new_n332), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G87), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n439), .A2(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n709), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n280), .B1(new_n725), .B2(new_n223), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n719), .A2(new_n709), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n545), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n720), .A2(new_n724), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n726), .B(new_n728), .C1(G58), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n715), .A2(G190), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G68), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n717), .A2(new_n723), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n725), .ZN(new_n735));
  AOI22_X1  g0535(.A1(G311), .A2(new_n735), .B1(new_n711), .B2(G329), .ZN(new_n736));
  INV_X1    g0536(.A(G322), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n270), .C1(new_n737), .C2(new_n729), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(G294), .B2(new_n706), .ZN(new_n739));
  INV_X1    g0539(.A(new_n727), .ZN(new_n740));
  AOI22_X1  g0540(.A1(G283), .A2(new_n740), .B1(new_n722), .B2(G303), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT33), .B(G317), .ZN(new_n742));
  AOI22_X1  g0542(.A1(G326), .A2(new_n716), .B1(new_n732), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n703), .B1(new_n734), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n702), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n217), .A2(new_n270), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G355), .A2(new_n750), .B1(new_n458), .B2(new_n217), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n252), .A2(new_n582), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n217), .A2(new_n280), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G45), .B2(new_n208), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n700), .B(new_n745), .C1(new_n749), .C2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n748), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n756), .B1(new_n641), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n701), .A2(new_n758), .ZN(G396));
  NAND2_X1  g0559(.A1(new_n399), .A2(new_n636), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n402), .A2(new_n400), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT99), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT99), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n402), .A2(new_n400), .A3(new_n763), .A4(new_n760), .ZN(new_n764));
  AOI221_X4 g0564(.A(new_n636), .B1(new_n762), .B2(new_n764), .C1(new_n608), .C2(new_n614), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n400), .A2(new_n637), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n762), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n766), .B1(new_n692), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n684), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n699), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n702), .A2(new_n746), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n699), .B1(G77), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n740), .A2(G87), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G107), .B2(new_n722), .ZN(new_n778));
  INV_X1    g0578(.A(G294), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n270), .B1(new_n729), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n725), .A2(new_n458), .B1(new_n710), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n708), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT96), .B(G283), .Z(new_n784));
  AOI22_X1  g0584(.A1(G303), .A2(new_n716), .B1(new_n732), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n778), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n740), .A2(G68), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n202), .B2(new_n721), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT98), .Z(new_n789));
  INV_X1    g0589(.A(G132), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n280), .B1(new_n710), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G58), .B2(new_n706), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G143), .A2(new_n730), .B1(new_n735), .B2(G159), .ZN(new_n793));
  INV_X1    g0593(.A(new_n716), .ZN(new_n794));
  INV_X1    g0594(.A(G137), .ZN(new_n795));
  INV_X1    g0595(.A(G150), .ZN(new_n796));
  INV_X1    g0596(.A(new_n732), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n793), .B1(new_n794), .B2(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n799));
  OAI211_X1 g0599(.A(new_n789), .B(new_n792), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n786), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n776), .B1(new_n802), .B2(new_n702), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n769), .B2(new_n747), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n773), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G384));
  INV_X1    g0606(.A(new_n543), .ZN(new_n807));
  OAI211_X1 g0607(.A(G116), .B(new_n212), .C1(new_n807), .C2(KEYINPUT35), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(KEYINPUT35), .B2(new_n807), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT36), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n209), .B(G77), .C1(new_n228), .C2(new_n230), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n287), .B(G13), .C1(new_n811), .C2(new_n248), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT100), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n400), .A2(new_n636), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n762), .A2(new_n764), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n692), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n377), .A2(new_n636), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n378), .A2(new_n818), .B1(new_n619), .B2(new_n636), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n814), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n819), .ZN(new_n821));
  OAI211_X1 g0621(.A(KEYINPUT100), .B(new_n821), .C1(new_n765), .C2(new_n815), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n634), .B1(new_n285), .B2(new_n291), .ZN(new_n823));
  INV_X1    g0623(.A(new_n292), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n336), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT37), .B1(new_n322), .B2(KEYINPUT104), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(KEYINPUT104), .C2(new_n322), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n262), .B1(new_n269), .B2(new_n275), .ZN(new_n828));
  NOR2_X1   g0628(.A1(KEYINPUT101), .A2(KEYINPUT16), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n259), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n829), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n267), .A2(new_n274), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n832), .B(G68), .C1(new_n268), .C2(new_n267), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(new_n262), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n291), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n318), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n836), .A2(KEYINPUT103), .A3(new_n330), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT103), .B1(new_n836), .B2(new_n330), .ZN(new_n838));
  INV_X1    g0638(.A(new_n634), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n837), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n827), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT102), .B1(new_n340), .B2(new_n841), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT102), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n846), .B(new_n840), .C1(new_n327), .C2(new_n339), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n844), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT105), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  OAI211_X1 g0652(.A(KEYINPUT38), .B(new_n844), .C1(new_n845), .C2(new_n847), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(KEYINPUT105), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n820), .A2(new_n822), .A3(new_n851), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n326), .A2(new_n319), .A3(new_n634), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n619), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(new_n636), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n854), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT106), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n292), .A2(new_n839), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n330), .C1(KEYINPUT104), .C2(new_n322), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT104), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n843), .B1(new_n324), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n843), .B1(new_n825), .B2(new_n324), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n324), .A2(new_n863), .A3(new_n330), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n827), .A2(KEYINPUT106), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT107), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n326), .A2(new_n319), .B1(new_n331), .B2(new_n338), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n863), .ZN(new_n875));
  INV_X1    g0675(.A(new_n319), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n322), .A2(KEYINPUT18), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n339), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(KEYINPUT107), .A3(new_n823), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n869), .A2(new_n872), .A3(new_n875), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n850), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n853), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n860), .B1(new_n861), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n857), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n691), .A2(new_n443), .A3(new_n693), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n628), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT108), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n683), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n681), .A2(KEYINPUT108), .A3(new_n682), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n768), .B(new_n819), .C1(new_n680), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n854), .A2(new_n851), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n882), .A2(KEYINPUT109), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT109), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n881), .A2(new_n853), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n680), .A2(new_n892), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n769), .A3(new_n821), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n895), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n896), .A2(new_n904), .A3(G330), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n443), .A2(new_n901), .A3(G330), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n895), .A2(new_n894), .B1(new_n900), .B2(new_n903), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n443), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n888), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n287), .B2(new_n630), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n888), .B1(new_n907), .B2(new_n909), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n813), .B1(new_n911), .B2(new_n912), .ZN(G367));
  INV_X1    g0713(.A(new_n550), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n568), .B1(new_n914), .B2(new_n637), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n609), .B2(new_n637), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT110), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n653), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n609), .B1(new_n918), .B2(new_n529), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n637), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT111), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n581), .A2(new_n637), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n597), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n595), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n925), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n920), .A2(new_n921), .B1(new_n637), .B2(new_n923), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n931), .B1(new_n934), .B2(KEYINPUT111), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n926), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n651), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n916), .B(KEYINPUT110), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n935), .A3(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n941), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n943), .A2(new_n936), .B1(new_n651), .B2(new_n918), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n658), .B(KEYINPUT41), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n650), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n652), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n646), .A2(new_n653), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n646), .B1(new_n653), .B2(new_n948), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n656), .B2(new_n939), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n655), .A2(new_n918), .A3(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n656), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n655), .B2(new_n918), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n651), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n938), .A2(new_n960), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n951), .A2(new_n962), .A3(new_n694), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n946), .B1(new_n964), .B2(new_n694), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n942), .B(new_n944), .C1(new_n965), .C2(new_n698), .ZN(new_n966));
  INV_X1    g0766(.A(new_n753), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n242), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n749), .B1(new_n216), .B2(new_n392), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n699), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G143), .A2(new_n716), .B1(new_n732), .B2(G159), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n706), .A2(G68), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n729), .A2(new_n796), .B1(new_n710), .B2(new_n795), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n270), .B(new_n973), .C1(G50), .C2(new_n735), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G58), .A2(new_n722), .B1(new_n740), .B2(G77), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n722), .A2(G116), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT46), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n779), .B2(new_n797), .C1(new_n781), .C2(new_n794), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n740), .A2(G97), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n706), .A2(G107), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n280), .B1(new_n735), .B2(new_n784), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n730), .A2(G303), .B1(new_n711), .B2(G317), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n976), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT47), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n703), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n970), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n757), .B2(new_n931), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT112), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n966), .A2(new_n991), .ZN(G387));
  NAND2_X1  g0792(.A1(new_n951), .A2(new_n694), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT114), .B1(new_n993), .B2(new_n658), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n951), .A2(new_n694), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(KEYINPUT114), .A3(new_n658), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n951), .A2(new_n698), .ZN(new_n999));
  AOI211_X1 g0799(.A(G45), .B(new_n659), .C1(G68), .C2(G77), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT113), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(KEYINPUT113), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT50), .B1(new_n390), .B2(G50), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n390), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1005), .B(new_n753), .C1(new_n582), .C2(new_n239), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n750), .A2(new_n659), .B1(new_n545), .B2(new_n217), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n748), .B(new_n702), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G159), .A2(new_n716), .B1(new_n732), .B2(new_n286), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n707), .A2(new_n392), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n729), .A2(new_n202), .B1(new_n725), .B2(new_n230), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n280), .B1(new_n710), .B2(new_n796), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n722), .A2(G77), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1009), .A2(new_n980), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n280), .B1(new_n711), .B2(G326), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n721), .A2(new_n779), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G317), .A2(new_n730), .B1(new_n735), .B2(G303), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n794), .B2(new_n737), .C1(new_n781), .C2(new_n797), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT48), .Z(new_n1020));
  AOI211_X1 g0820(.A(new_n1017), .B(new_n1020), .C1(new_n706), .C2(new_n784), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1016), .B1(new_n458), .B2(new_n727), .C1(new_n1021), .C2(KEYINPUT49), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT49), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1015), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n700), .B(new_n1008), .C1(new_n1024), .C2(new_n702), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n947), .A2(new_n748), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n999), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n998), .A2(new_n1028), .ZN(G393));
  NOR2_X1   g0829(.A1(new_n938), .A2(new_n960), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n961), .A2(new_n651), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n993), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n964), .A2(new_n658), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT117), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1036), .A3(new_n658), .A4(new_n964), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n939), .A2(new_n757), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(KEYINPUT115), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(KEYINPUT115), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n716), .A2(G150), .B1(G159), .B2(new_n730), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT51), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n270), .B1(new_n711), .B2(G143), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n223), .B2(new_n707), .C1(new_n390), .C2(new_n725), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1046), .B(new_n777), .C1(G68), .C2(new_n722), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1044), .B(new_n1047), .C1(new_n202), .C2(new_n797), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n716), .A2(G317), .B1(G311), .B2(new_n730), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT52), .Z(new_n1050));
  AOI21_X1  g0850(.A(new_n280), .B1(new_n711), .B2(G322), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n458), .B2(new_n707), .C1(new_n779), .C2(new_n725), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n728), .B(new_n1052), .C1(new_n722), .C2(new_n784), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1050), .B(new_n1053), .C1(new_n445), .C2(new_n797), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n703), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n749), .B1(new_n225), .B2(new_n216), .C1(new_n247), .C2(new_n967), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT116), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n700), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1041), .A2(new_n1042), .A3(new_n1055), .A4(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1031), .A2(new_n1030), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n698), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1038), .A2(new_n1062), .ZN(G390));
  OAI21_X1  g0863(.A(new_n860), .B1(new_n817), .B2(new_n819), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n861), .A2(new_n883), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n684), .A2(new_n769), .A3(new_n821), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n816), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n689), .A2(new_n1067), .B1(new_n400), .B2(new_n636), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n859), .B1(new_n1068), .B2(new_n821), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n900), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1065), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT118), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT118), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1065), .A2(new_n1073), .A3(new_n1066), .A4(new_n1070), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1065), .A2(new_n1070), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n893), .A2(G330), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1072), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n628), .A2(new_n886), .A3(new_n906), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n680), .A2(new_n683), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(G330), .A3(new_n769), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n819), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n817), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1068), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n644), .B(new_n768), .C1(new_n680), .C2(new_n892), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1066), .B(new_n1087), .C1(new_n1088), .C2(new_n821), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1080), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1079), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1072), .A2(new_n1078), .A3(new_n1074), .A4(new_n1090), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(new_n658), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1072), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n861), .A2(new_n746), .A3(new_n883), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n699), .B1(new_n286), .B2(new_n775), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n716), .A2(G128), .B1(G132), .B2(new_n730), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT119), .Z(new_n1099));
  NOR2_X1   g0899(.A1(new_n721), .A2(new_n796), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n270), .B1(new_n711), .B2(G125), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n706), .A2(G159), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  NAND2_X1  g0904(.A1(new_n735), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n727), .A2(new_n202), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G137), .C2(new_n732), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1099), .A2(new_n1101), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n270), .B1(new_n710), .B2(new_n779), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n729), .A2(new_n458), .B1(new_n725), .B2(new_n225), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G77), .C2(new_n706), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n723), .A3(new_n787), .ZN(new_n1113));
  INV_X1    g0913(.A(G283), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n545), .A2(new_n797), .B1(new_n794), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1109), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1097), .B1(new_n1116), .B2(new_n702), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1095), .A2(new_n698), .B1(new_n1096), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1094), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT120), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1094), .A2(new_n1118), .A3(KEYINPUT120), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(new_n884), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n856), .A3(new_n855), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n426), .A2(new_n839), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT55), .B1(new_n626), .B2(new_n441), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT55), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n437), .A2(new_n1129), .A3(new_n442), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1127), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n626), .A2(KEYINPUT55), .A3(new_n441), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1129), .B1(new_n437), .B2(new_n442), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n1126), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1131), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1132), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n908), .B2(G330), .ZN(new_n1139));
  AND4_X1   g0939(.A1(G330), .A2(new_n896), .A3(new_n904), .A4(new_n1138), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1125), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n905), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n908), .A2(G330), .A3(new_n1138), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n885), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(KEYINPUT122), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1080), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1093), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT122), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1143), .A2(new_n885), .A3(new_n1144), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n658), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1152), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n1148), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1146), .A2(new_n698), .A3(new_n1150), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1142), .A2(new_n746), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n730), .B1(new_n735), .B2(G137), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n796), .B2(new_n707), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n722), .B2(new_n1104), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n716), .A2(G125), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n790), .C2(new_n797), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n740), .A2(G159), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G33), .B(G41), .C1(new_n711), .C2(G124), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G97), .A2(new_n732), .B1(new_n716), .B2(G116), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n300), .B(new_n270), .C1(new_n729), .C2(new_n545), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n725), .A2(new_n392), .B1(new_n710), .B2(new_n1114), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G58), .A2(new_n740), .B1(new_n722), .B2(G77), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1170), .A2(new_n972), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G50), .B1(new_n263), .B2(new_n300), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n280), .B2(G41), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1169), .A2(new_n1177), .A3(new_n1178), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n702), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n774), .A2(new_n202), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1159), .A2(new_n699), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1158), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1157), .A2(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n698), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n700), .B1(new_n230), .B2(new_n774), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n730), .A2(G137), .B1(new_n711), .B2(G128), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n202), .B2(new_n707), .C1(new_n796), .C2(new_n725), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G132), .A2(new_n716), .B1(new_n732), .B2(new_n1104), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(G159), .C2(new_n722), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n280), .B1(new_n727), .B2(new_n228), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT124), .Z(new_n1197));
  AOI22_X1  g0997(.A1(G77), .A2(new_n740), .B1(new_n722), .B2(G97), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n270), .B1(new_n710), .B2(new_n445), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n729), .A2(new_n1114), .B1(new_n725), .B2(new_n545), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1199), .A2(new_n1010), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G116), .A2(new_n732), .B1(new_n716), .B2(G294), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1195), .A2(new_n1197), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1190), .B1(new_n703), .B2(new_n1204), .C1(new_n821), .C2(new_n747), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1189), .A2(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n945), .B(KEYINPUT123), .Z(new_n1207));
  NOR2_X1   g1007(.A1(new_n1090), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1188), .A2(new_n1147), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1206), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(G381));
  NOR2_X1   g1012(.A1(G375), .A2(new_n1119), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n966), .A2(new_n1038), .A3(new_n991), .A4(new_n1062), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n998), .A2(new_n701), .A3(new_n758), .A4(new_n1028), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1216), .A2(G384), .A3(G381), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1215), .A3(new_n1217), .ZN(G407));
  NAND2_X1  g1018(.A1(new_n1213), .A2(new_n635), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  AOI21_X1  g1020(.A(KEYINPUT120), .B1(new_n1094), .B2(new_n1118), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1094), .A2(new_n1118), .A3(KEYINPUT120), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1157), .B(new_n1186), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1207), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .A4(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1184), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n698), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1119), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1223), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G343), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n658), .B(new_n1091), .C1(new_n1209), .C2(KEYINPUT60), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT125), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1209), .A2(new_n1239), .A3(KEYINPUT60), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1236), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  OR3_X1    g1041(.A1(new_n1241), .A2(new_n805), .A3(new_n1206), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n805), .B1(new_n1241), .B2(new_n1206), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1233), .A2(G2897), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1244), .B(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT61), .B1(new_n1235), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1233), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1244), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT63), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(G390), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n997), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1255), .A2(new_n995), .A3(new_n994), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1028), .ZN(new_n1257));
  OAI21_X1  g1057(.A(G396), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1216), .A2(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1254), .A2(new_n1214), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1254), .B2(new_n1214), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1247), .A2(new_n1252), .A3(new_n1253), .A4(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1244), .A2(G2897), .A3(new_n1233), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1264), .B1(new_n1267), .B2(new_n1248), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1185), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1229), .B1(new_n1271), .B2(G378), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(new_n1272), .A2(KEYINPUT62), .A3(new_n1244), .A4(new_n1233), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1268), .A2(new_n1270), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1263), .B1(new_n1274), .B2(new_n1262), .ZN(G405));
  NAND3_X1  g1075(.A1(G375), .A2(new_n1094), .A3(new_n1118), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1223), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1262), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1223), .B(new_n1276), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1249), .A2(KEYINPUT126), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1278), .A2(new_n1279), .A3(KEYINPUT126), .A4(new_n1249), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(G402));
endmodule


