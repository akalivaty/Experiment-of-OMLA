

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752;

  AND2_X1 U375 ( .A1(n441), .A2(G224), .ZN(n407) );
  NOR2_X2 U376 ( .A1(n538), .A2(n600), .ZN(n539) );
  NOR2_X1 U377 ( .A1(n752), .A2(n751), .ZN(n576) );
  NOR2_X1 U378 ( .A1(n518), .A2(n693), .ZN(n474) );
  INV_X2 U379 ( .A(G953), .ZN(n441) );
  AND2_X1 U380 ( .A1(n401), .A2(n396), .ZN(n369) );
  XNOR2_X1 U381 ( .A(n374), .B(n575), .ZN(n751) );
  NOR2_X1 U382 ( .A1(n528), .A2(n354), .ZN(n371) );
  INV_X2 U383 ( .A(n518), .ZN(n535) );
  BUF_X2 U384 ( .A(n688), .Z(n353) );
  XNOR2_X1 U385 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n408) );
  XOR2_X1 U386 ( .A(KEYINPUT4), .B(G146), .Z(n440) );
  OR2_X1 U387 ( .A1(n418), .A2(n444), .ZN(n377) );
  XNOR2_X1 U388 ( .A(n515), .B(n438), .ZN(n528) );
  NOR2_X1 U389 ( .A1(n713), .A2(n528), .ZN(n529) );
  XNOR2_X1 U390 ( .A(n554), .B(n553), .ZN(n623) );
  NAND2_X1 U391 ( .A1(n395), .A2(n362), .ZN(n394) );
  XNOR2_X2 U392 ( .A(n534), .B(n533), .ZN(n647) );
  NAND2_X1 U393 ( .A1(n623), .A2(n742), .ZN(n402) );
  INV_X1 U394 ( .A(n395), .ZN(n352) );
  NAND2_X1 U395 ( .A1(n648), .A2(n621), .ZN(n372) );
  INV_X1 U396 ( .A(G128), .ZN(n415) );
  NAND2_X1 U397 ( .A1(n639), .A2(n638), .ZN(n548) );
  XNOR2_X1 U398 ( .A(n439), .B(n406), .ZN(n405) );
  XNOR2_X1 U399 ( .A(n404), .B(n440), .ZN(n403) );
  XNOR2_X1 U400 ( .A(n407), .B(n414), .ZN(n406) );
  XNOR2_X1 U401 ( .A(n379), .B(n355), .ZN(n578) );
  XNOR2_X1 U402 ( .A(G113), .B(KEYINPUT70), .ZN(n419) );
  XNOR2_X1 U403 ( .A(G101), .B(G110), .ZN(n416) );
  XNOR2_X1 U404 ( .A(G119), .B(G128), .ZN(n449) );
  XNOR2_X1 U405 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n450) );
  XNOR2_X1 U406 ( .A(G116), .B(G107), .ZN(n498) );
  XNOR2_X1 U407 ( .A(n385), .B(n502), .ZN(n741) );
  XNOR2_X1 U408 ( .A(n440), .B(n367), .ZN(n385) );
  XNOR2_X1 U409 ( .A(n368), .B(G137), .ZN(n367) );
  INV_X1 U410 ( .A(G131), .ZN(n368) );
  XNOR2_X1 U411 ( .A(n375), .B(n571), .ZN(n722) );
  NOR2_X1 U412 ( .A1(n709), .A2(n708), .ZN(n375) );
  NAND2_X1 U413 ( .A1(n562), .A2(n389), .ZN(n388) );
  AND2_X1 U414 ( .A1(n392), .A2(n391), .ZN(n390) );
  NOR2_X1 U415 ( .A1(n598), .A2(n393), .ZN(n389) );
  OR2_X1 U416 ( .A1(n597), .A2(KEYINPUT85), .ZN(n384) );
  INV_X1 U417 ( .A(KEYINPUT66), .ZN(n400) );
  XNOR2_X1 U418 ( .A(n408), .B(n409), .ZN(n404) );
  XNOR2_X1 U419 ( .A(n587), .B(KEYINPUT38), .ZN(n705) );
  XNOR2_X1 U420 ( .A(G119), .B(G116), .ZN(n420) );
  XOR2_X1 U421 ( .A(G122), .B(G104), .Z(n480) );
  NAND2_X1 U422 ( .A1(n399), .A2(n397), .ZN(n396) );
  NAND2_X1 U423 ( .A1(n621), .A2(n400), .ZN(n399) );
  NAND2_X1 U424 ( .A1(n622), .A2(n398), .ZN(n397) );
  NAND2_X1 U425 ( .A1(KEYINPUT2), .A2(n400), .ZN(n398) );
  INV_X1 U426 ( .A(KEYINPUT28), .ZN(n393) );
  NAND2_X1 U427 ( .A1(n598), .A2(n393), .ZN(n391) );
  XNOR2_X1 U428 ( .A(n373), .B(n735), .ZN(n648) );
  NOR2_X1 U429 ( .A1(n561), .A2(n572), .ZN(n585) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n641) );
  INV_X1 U431 ( .A(KEYINPUT98), .ZN(n370) );
  NOR2_X1 U432 ( .A1(n519), .A2(n535), .ZN(n544) );
  XOR2_X1 U433 ( .A(G101), .B(KEYINPUT5), .Z(n465) );
  XNOR2_X1 U434 ( .A(n491), .B(n456), .ZN(n660) );
  XNOR2_X1 U435 ( .A(n504), .B(n503), .ZN(n629) );
  XNOR2_X1 U436 ( .A(n445), .B(n741), .ZN(n663) );
  OR2_X2 U437 ( .A1(n580), .A2(n722), .ZN(n374) );
  NAND2_X1 U438 ( .A1(n532), .A2(n588), .ZN(n534) );
  AND2_X1 U439 ( .A1(n475), .A2(n699), .ZN(n476) );
  AND2_X1 U440 ( .A1(n387), .A2(n386), .ZN(n582) );
  NOR2_X1 U441 ( .A1(n579), .A2(n472), .ZN(n386) );
  OR2_X1 U442 ( .A1(n561), .A2(n562), .ZN(n354) );
  XNOR2_X1 U443 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n355) );
  XOR2_X1 U444 ( .A(G110), .B(G137), .Z(n356) );
  AND2_X1 U445 ( .A1(n352), .A2(n620), .ZN(n357) );
  XOR2_X1 U446 ( .A(KEYINPUT91), .B(KEYINPUT0), .Z(n358) );
  XNOR2_X1 U447 ( .A(KEYINPUT15), .B(G902), .ZN(n621) );
  XOR2_X1 U448 ( .A(n656), .B(n655), .Z(n359) );
  XOR2_X1 U449 ( .A(n634), .B(n633), .Z(n360) );
  XOR2_X1 U450 ( .A(n651), .B(n650), .Z(n361) );
  AND2_X1 U451 ( .A1(n622), .A2(n400), .ZN(n362) );
  AND2_X1 U452 ( .A1(n620), .A2(KEYINPUT66), .ZN(n363) );
  XNOR2_X1 U453 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n364) );
  NOR2_X1 U454 ( .A1(n744), .A2(G952), .ZN(n666) );
  XOR2_X1 U455 ( .A(KEYINPUT124), .B(KEYINPUT56), .Z(n365) );
  XNOR2_X1 U456 ( .A(n405), .B(n403), .ZN(n418) );
  NAND2_X1 U457 ( .A1(n369), .A2(n394), .ZN(n628) );
  NAND2_X1 U458 ( .A1(n366), .A2(n552), .ZN(n554) );
  NOR2_X1 U459 ( .A1(n551), .A2(n550), .ZN(n366) );
  XNOR2_X2 U460 ( .A(n417), .B(n416), .ZN(n733) );
  BUF_X1 U461 ( .A(n441), .Z(n744) );
  NOR2_X2 U462 ( .A1(n578), .A2(n437), .ZN(n378) );
  XNOR2_X2 U463 ( .A(n372), .B(n429), .ZN(n555) );
  NAND2_X1 U464 ( .A1(n377), .A2(n376), .ZN(n373) );
  NAND2_X1 U465 ( .A1(n418), .A2(n444), .ZN(n376) );
  XNOR2_X2 U466 ( .A(n378), .B(n358), .ZN(n515) );
  NAND2_X1 U467 ( .A1(n555), .A2(n704), .ZN(n379) );
  XNOR2_X2 U468 ( .A(n517), .B(n516), .ZN(n540) );
  XNOR2_X2 U469 ( .A(n733), .B(KEYINPUT72), .ZN(n444) );
  NAND2_X1 U470 ( .A1(n402), .A2(n363), .ZN(n401) );
  BUF_X2 U471 ( .A(n659), .Z(n661) );
  XNOR2_X1 U472 ( .A(n380), .B(n365), .ZN(G51) );
  NAND2_X1 U473 ( .A1(n654), .A2(n653), .ZN(n380) );
  XNOR2_X1 U474 ( .A(n381), .B(n364), .ZN(G60) );
  NAND2_X1 U475 ( .A1(n658), .A2(n653), .ZN(n381) );
  XNOR2_X1 U476 ( .A(n382), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U477 ( .A1(n636), .A2(n653), .ZN(n382) );
  NAND2_X1 U478 ( .A1(n383), .A2(n685), .ZN(n606) );
  NAND2_X1 U479 ( .A1(n384), .A2(n577), .ZN(n383) );
  XNOR2_X1 U480 ( .A(n439), .B(G134), .ZN(n502) );
  XNOR2_X2 U481 ( .A(n410), .B(n415), .ZN(n439) );
  NAND2_X1 U482 ( .A1(n387), .A2(n574), .ZN(n580) );
  NAND2_X1 U483 ( .A1(n390), .A2(n388), .ZN(n387) );
  NAND2_X1 U484 ( .A1(n692), .A2(n393), .ZN(n392) );
  INV_X1 U485 ( .A(n402), .ZN(n395) );
  XNOR2_X2 U486 ( .A(G125), .B(KEYINPUT18), .ZN(n409) );
  XNOR2_X2 U487 ( .A(G143), .B(KEYINPUT65), .ZN(n410) );
  AND2_X1 U488 ( .A1(n411), .A2(n653), .ZN(G66) );
  XNOR2_X1 U489 ( .A(n412), .B(n660), .ZN(n411) );
  NAND2_X1 U490 ( .A1(n661), .A2(G217), .ZN(n412) );
  INV_X1 U491 ( .A(n624), .ZN(n627) );
  NAND2_X1 U492 ( .A1(n624), .A2(n744), .ZN(n732) );
  XNOR2_X1 U493 ( .A(n630), .B(n629), .ZN(n631) );
  XOR2_X1 U494 ( .A(n453), .B(n452), .Z(n413) );
  INV_X1 U495 ( .A(KEYINPUT87), .ZN(n566) );
  XNOR2_X1 U496 ( .A(n566), .B(KEYINPUT39), .ZN(n567) );
  XNOR2_X2 U497 ( .A(KEYINPUT17), .B(KEYINPUT81), .ZN(n414) );
  XOR2_X1 U498 ( .A(G104), .B(G107), .Z(n417) );
  XNOR2_X1 U499 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U500 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n421) );
  XNOR2_X1 U501 ( .A(n422), .B(n421), .ZN(n467) );
  XNOR2_X1 U502 ( .A(KEYINPUT16), .B(G122), .ZN(n423) );
  XNOR2_X1 U503 ( .A(n423), .B(KEYINPUT73), .ZN(n424) );
  XNOR2_X1 U504 ( .A(n467), .B(n424), .ZN(n735) );
  NOR2_X1 U505 ( .A1(G237), .A2(G902), .ZN(n425) );
  XNOR2_X1 U506 ( .A(n425), .B(KEYINPUT76), .ZN(n431) );
  INV_X1 U507 ( .A(G210), .ZN(n426) );
  OR2_X1 U508 ( .A1(n431), .A2(n426), .ZN(n428) );
  XNOR2_X1 U509 ( .A(KEYINPUT84), .B(KEYINPUT93), .ZN(n427) );
  XNOR2_X1 U510 ( .A(n428), .B(n427), .ZN(n429) );
  INV_X1 U511 ( .A(G214), .ZN(n430) );
  OR2_X1 U512 ( .A1(n431), .A2(n430), .ZN(n704) );
  XOR2_X1 U513 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n433) );
  NAND2_X1 U514 ( .A1(G234), .A2(G237), .ZN(n432) );
  XOR2_X1 U515 ( .A(n433), .B(n432), .Z(n435) );
  AND2_X1 U516 ( .A1(n435), .A2(G953), .ZN(n434) );
  NAND2_X1 U517 ( .A1(G902), .A2(n434), .ZN(n557) );
  NOR2_X1 U518 ( .A1(n557), .A2(G898), .ZN(n436) );
  NAND2_X1 U519 ( .A1(G952), .A2(n435), .ZN(n719) );
  NOR2_X1 U520 ( .A1(n719), .A2(G953), .ZN(n560) );
  NOR2_X1 U521 ( .A1(n436), .A2(n560), .ZN(n437) );
  INV_X1 U522 ( .A(KEYINPUT94), .ZN(n438) );
  NAND2_X1 U523 ( .A1(G227), .A2(n744), .ZN(n442) );
  INV_X1 U524 ( .A(G140), .ZN(n644) );
  XNOR2_X1 U525 ( .A(n442), .B(n644), .ZN(n443) );
  XNOR2_X1 U526 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U527 ( .A(G902), .ZN(n505) );
  NAND2_X1 U528 ( .A1(n663), .A2(n505), .ZN(n447) );
  INV_X1 U529 ( .A(G469), .ZN(n446) );
  XNOR2_X2 U530 ( .A(n447), .B(n446), .ZN(n472) );
  XOR2_X1 U531 ( .A(G125), .B(KEYINPUT10), .Z(n448) );
  XNOR2_X1 U532 ( .A(G140), .B(n448), .ZN(n740) );
  XNOR2_X1 U533 ( .A(n740), .B(G146), .ZN(n491) );
  XNOR2_X1 U534 ( .A(n356), .B(n449), .ZN(n453) );
  XOR2_X1 U535 ( .A(KEYINPUT78), .B(KEYINPUT95), .Z(n451) );
  XNOR2_X1 U536 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U537 ( .A1(G234), .A2(n441), .ZN(n454) );
  XOR2_X1 U538 ( .A(KEYINPUT8), .B(n454), .Z(n495) );
  NAND2_X1 U539 ( .A1(G221), .A2(n495), .ZN(n455) );
  XNOR2_X1 U540 ( .A(n413), .B(n455), .ZN(n456) );
  NAND2_X1 U541 ( .A1(n660), .A2(n505), .ZN(n460) );
  NAND2_X1 U542 ( .A1(G234), .A2(n621), .ZN(n457) );
  XNOR2_X1 U543 ( .A(KEYINPUT20), .B(n457), .ZN(n461) );
  AND2_X1 U544 ( .A1(G217), .A2(n461), .ZN(n458) );
  XNOR2_X1 U545 ( .A(KEYINPUT25), .B(n458), .ZN(n459) );
  XNOR2_X2 U546 ( .A(n460), .B(n459), .ZN(n688) );
  AND2_X1 U547 ( .A1(n461), .A2(G221), .ZN(n463) );
  XNOR2_X1 U548 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n462) );
  XNOR2_X1 U549 ( .A(n463), .B(n462), .ZN(n689) );
  NAND2_X1 U550 ( .A1(n353), .A2(n689), .ZN(n693) );
  OR2_X1 U551 ( .A1(n472), .A2(n693), .ZN(n561) );
  NOR2_X1 U552 ( .A1(G953), .A2(G237), .ZN(n485) );
  NAND2_X1 U553 ( .A1(n485), .A2(G210), .ZN(n464) );
  XOR2_X1 U554 ( .A(n465), .B(n464), .Z(n466) );
  XNOR2_X1 U555 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U556 ( .A(n741), .B(n468), .ZN(n634) );
  NAND2_X1 U557 ( .A1(n634), .A2(n505), .ZN(n471) );
  INV_X1 U558 ( .A(KEYINPUT97), .ZN(n469) );
  XNOR2_X1 U559 ( .A(n469), .B(G472), .ZN(n470) );
  XNOR2_X2 U560 ( .A(n471), .B(n470), .ZN(n562) );
  INV_X1 U561 ( .A(n562), .ZN(n692) );
  AND2_X1 U562 ( .A1(n515), .A2(n562), .ZN(n475) );
  XNOR2_X1 U563 ( .A(n472), .B(KEYINPUT1), .ZN(n518) );
  INV_X1 U564 ( .A(KEYINPUT75), .ZN(n473) );
  XNOR2_X1 U565 ( .A(n474), .B(n473), .ZN(n699) );
  XNOR2_X2 U566 ( .A(n476), .B(KEYINPUT31), .ZN(n681) );
  NAND2_X1 U567 ( .A1(n641), .A2(n681), .ZN(n478) );
  INV_X1 U568 ( .A(KEYINPUT99), .ZN(n477) );
  XNOR2_X1 U569 ( .A(n478), .B(n477), .ZN(n511) );
  XNOR2_X1 U570 ( .A(G113), .B(G131), .ZN(n479) );
  XNOR2_X1 U571 ( .A(n480), .B(n479), .ZN(n484) );
  XOR2_X1 U572 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n482) );
  XNOR2_X1 U573 ( .A(G143), .B(KEYINPUT102), .ZN(n481) );
  XNOR2_X1 U574 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U575 ( .A(n484), .B(n483), .ZN(n489) );
  XOR2_X1 U576 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n487) );
  NAND2_X1 U577 ( .A1(G214), .A2(n485), .ZN(n486) );
  XNOR2_X1 U578 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U579 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U580 ( .A(n491), .B(n490), .ZN(n656) );
  NOR2_X1 U581 ( .A1(G902), .A2(n656), .ZN(n493) );
  XNOR2_X1 U582 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n492) );
  XNOR2_X1 U583 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U584 ( .A(n494), .B(G475), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G217), .A2(n495), .ZN(n497) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n496) );
  XNOR2_X1 U587 ( .A(n497), .B(n496), .ZN(n501) );
  XOR2_X1 U588 ( .A(KEYINPUT9), .B(G122), .Z(n499) );
  XNOR2_X1 U589 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n504) );
  INV_X1 U591 ( .A(n502), .ZN(n503) );
  NAND2_X1 U592 ( .A1(n629), .A2(n505), .ZN(n507) );
  INV_X1 U593 ( .A(G478), .ZN(n506) );
  XNOR2_X1 U594 ( .A(n507), .B(n506), .ZN(n530) );
  INV_X1 U595 ( .A(n530), .ZN(n508) );
  AND2_X1 U596 ( .A1(n531), .A2(n508), .ZN(n673) );
  INV_X1 U597 ( .A(n673), .ZN(n668) );
  OR2_X1 U598 ( .A1(n531), .A2(n508), .ZN(n680) );
  NAND2_X1 U599 ( .A1(n668), .A2(n680), .ZN(n510) );
  INV_X1 U600 ( .A(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n510), .B(n509), .ZN(n577) );
  NAND2_X1 U602 ( .A1(n511), .A2(n577), .ZN(n512) );
  XNOR2_X1 U603 ( .A(n512), .B(KEYINPUT106), .ZN(n524) );
  NAND2_X1 U604 ( .A1(n531), .A2(n530), .ZN(n708) );
  INV_X1 U605 ( .A(n689), .ZN(n513) );
  NOR2_X1 U606 ( .A1(n708), .A2(n513), .ZN(n514) );
  NAND2_X1 U607 ( .A1(n515), .A2(n514), .ZN(n517) );
  XOR2_X1 U608 ( .A(KEYINPUT68), .B(KEYINPUT22), .Z(n516) );
  INV_X1 U609 ( .A(n540), .ZN(n519) );
  INV_X1 U610 ( .A(n544), .ZN(n521) );
  INV_X1 U611 ( .A(KEYINPUT6), .ZN(n520) );
  XNOR2_X1 U612 ( .A(n562), .B(n520), .ZN(n600) );
  NOR2_X1 U613 ( .A1(n521), .A2(n600), .ZN(n522) );
  XNOR2_X1 U614 ( .A(n522), .B(KEYINPUT88), .ZN(n523) );
  NAND2_X1 U615 ( .A1(n523), .A2(n353), .ZN(n646) );
  NAND2_X1 U616 ( .A1(n524), .A2(n646), .ZN(n525) );
  XNOR2_X1 U617 ( .A(n525), .B(KEYINPUT107), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n699), .A2(n600), .ZN(n527) );
  XNOR2_X1 U619 ( .A(KEYINPUT109), .B(KEYINPUT33), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n527), .B(n526), .ZN(n713) );
  XNOR2_X1 U621 ( .A(n529), .B(KEYINPUT34), .ZN(n532) );
  NOR2_X1 U622 ( .A1(n531), .A2(n530), .ZN(n588) );
  INV_X1 U623 ( .A(KEYINPUT35), .ZN(n533) );
  XNOR2_X1 U624 ( .A(n647), .B(KEYINPUT44), .ZN(n547) );
  INV_X1 U625 ( .A(KEYINPUT108), .ZN(n537) );
  INV_X1 U626 ( .A(n535), .ZN(n694) );
  NOR2_X1 U627 ( .A1(n694), .A2(n353), .ZN(n536) );
  XNOR2_X1 U628 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U629 ( .A(n539), .B(KEYINPUT82), .ZN(n541) );
  NAND2_X1 U630 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X2 U631 ( .A(n542), .B(KEYINPUT32), .ZN(n639) );
  NOR2_X1 U632 ( .A1(n562), .A2(n353), .ZN(n543) );
  NAND2_X1 U633 ( .A1(n544), .A2(n543), .ZN(n638) );
  XNOR2_X1 U634 ( .A(n548), .B(KEYINPUT89), .ZN(n545) );
  NOR2_X1 U635 ( .A1(n545), .A2(KEYINPUT44), .ZN(n546) );
  NOR2_X1 U636 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U637 ( .A1(n548), .A2(KEYINPUT44), .ZN(n549) );
  XNOR2_X1 U638 ( .A(n549), .B(KEYINPUT67), .ZN(n550) );
  XNOR2_X1 U639 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n553) );
  BUF_X1 U640 ( .A(n555), .Z(n556) );
  INV_X1 U641 ( .A(n556), .ZN(n587) );
  XNOR2_X1 U642 ( .A(n557), .B(KEYINPUT110), .ZN(n558) );
  NOR2_X1 U643 ( .A1(G900), .A2(n558), .ZN(n559) );
  NOR2_X1 U644 ( .A1(n560), .A2(n559), .ZN(n572) );
  AND2_X1 U645 ( .A1(n705), .A2(n585), .ZN(n565) );
  NAND2_X1 U646 ( .A1(n562), .A2(n704), .ZN(n563) );
  XNOR2_X1 U647 ( .A(n563), .B(KEYINPUT30), .ZN(n564) );
  XNOR2_X1 U648 ( .A(KEYINPUT113), .B(n564), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n565), .A2(n586), .ZN(n568) );
  XNOR2_X1 U650 ( .A(n568), .B(n567), .ZN(n611) );
  INV_X1 U651 ( .A(n680), .ZN(n677) );
  AND2_X1 U652 ( .A1(n611), .A2(n677), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n569), .B(KEYINPUT40), .ZN(n752) );
  XNOR2_X1 U654 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n570) );
  XNOR2_X1 U655 ( .A(n570), .B(KEYINPUT42), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n705), .A2(n704), .ZN(n709) );
  XNOR2_X1 U657 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n571) );
  NOR2_X1 U658 ( .A1(n572), .A2(n353), .ZN(n573) );
  NAND2_X1 U659 ( .A1(n689), .A2(n573), .ZN(n598) );
  INV_X1 U660 ( .A(n472), .ZN(n574) );
  XNOR2_X1 U661 ( .A(n576), .B(KEYINPUT46), .ZN(n609) );
  INV_X1 U662 ( .A(n577), .ZN(n710) );
  INV_X1 U663 ( .A(KEYINPUT85), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n710), .A2(n591), .ZN(n583) );
  BUF_X1 U665 ( .A(n578), .Z(n579) );
  INV_X1 U666 ( .A(KEYINPUT83), .ZN(n581) );
  XNOR2_X1 U667 ( .A(n582), .B(n581), .ZN(n678) );
  NAND2_X1 U668 ( .A1(n583), .A2(n678), .ZN(n584) );
  NAND2_X1 U669 ( .A1(n584), .A2(KEYINPUT47), .ZN(n595) );
  AND2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n590) );
  INV_X1 U671 ( .A(n587), .ZN(n615) );
  AND2_X1 U672 ( .A1(n588), .A2(n615), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n637) );
  INV_X1 U674 ( .A(n637), .ZN(n593) );
  NOR2_X1 U675 ( .A1(KEYINPUT47), .A2(n591), .ZN(n592) );
  NOR2_X1 U676 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U677 ( .A1(n595), .A2(n594), .ZN(n607) );
  INV_X1 U678 ( .A(n678), .ZN(n596) );
  NOR2_X1 U679 ( .A1(n596), .A2(KEYINPUT47), .ZN(n597) );
  NOR2_X1 U680 ( .A1(n680), .A2(n598), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U682 ( .A(n601), .B(KEYINPUT111), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n602), .A2(n704), .ZN(n612) );
  INV_X1 U684 ( .A(n615), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n612), .A2(n603), .ZN(n604) );
  XNOR2_X1 U686 ( .A(n604), .B(KEYINPUT36), .ZN(n605) );
  NAND2_X1 U687 ( .A1(n605), .A2(n535), .ZN(n685) );
  NOR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n608) );
  AND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U690 ( .A(n610), .B(KEYINPUT48), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n673), .A2(n611), .ZN(n686) );
  INV_X1 U692 ( .A(n686), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT112), .B(n612), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n535), .A2(n613), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n614), .B(KEYINPUT43), .ZN(n616) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n645) );
  NOR2_X1 U697 ( .A1(n617), .A2(n645), .ZN(n618) );
  AND2_X2 U698 ( .A1(n619), .A2(n618), .ZN(n742) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n620) );
  INV_X1 U700 ( .A(n621), .ZN(n622) );
  BUF_X1 U701 ( .A(n623), .Z(n624) );
  NAND2_X1 U702 ( .A1(n742), .A2(KEYINPUT2), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT86), .ZN(n626) );
  NOR2_X2 U704 ( .A1(n627), .A2(n626), .ZN(n687) );
  NOR2_X4 U705 ( .A1(n628), .A2(n687), .ZN(n659) );
  NAND2_X1 U706 ( .A1(n661), .A2(G478), .ZN(n630) );
  AND2_X1 U707 ( .A1(n631), .A2(n653), .ZN(G63) );
  NAND2_X1 U708 ( .A1(n659), .A2(G472), .ZN(n635) );
  XNOR2_X1 U709 ( .A(KEYINPUT92), .B(KEYINPUT117), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n632), .B(KEYINPUT62), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n635), .B(n360), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n637), .B(G143), .ZN(G45) );
  XNOR2_X1 U713 ( .A(n638), .B(G110), .ZN(G12) );
  XNOR2_X1 U714 ( .A(n639), .B(G119), .ZN(G21) );
  NOR2_X1 U715 ( .A1(n681), .A2(n668), .ZN(n640) );
  XOR2_X1 U716 ( .A(G116), .B(n640), .Z(G18) );
  BUF_X1 U717 ( .A(n641), .Z(n642) );
  NOR2_X1 U718 ( .A1(n642), .A2(n680), .ZN(n643) );
  XOR2_X1 U719 ( .A(G104), .B(n643), .Z(G6) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(G42) );
  XNOR2_X1 U721 ( .A(n646), .B(G101), .ZN(G3) );
  XNOR2_X1 U722 ( .A(n647), .B(G122), .ZN(G24) );
  NAND2_X1 U723 ( .A1(n659), .A2(G210), .ZN(n652) );
  BUF_X1 U724 ( .A(n648), .Z(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n649), .B(KEYINPUT55), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n652), .B(n361), .ZN(n654) );
  INV_X1 U728 ( .A(n666), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n659), .A2(G475), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT125), .B(KEYINPUT59), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n657), .B(n359), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n661), .A2(G469), .ZN(n665) );
  XNOR2_X1 U733 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(G54) );
  XNOR2_X1 U737 ( .A(G107), .B(KEYINPUT27), .ZN(n672) );
  XOR2_X1 U738 ( .A(KEYINPUT118), .B(KEYINPUT26), .Z(n670) );
  NOR2_X1 U739 ( .A1(n642), .A2(n668), .ZN(n669) );
  XOR2_X1 U740 ( .A(n670), .B(n669), .Z(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(G9) );
  XOR2_X1 U742 ( .A(KEYINPUT29), .B(KEYINPUT119), .Z(n675) );
  NAND2_X1 U743 ( .A1(n678), .A2(n673), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(n676) );
  XOR2_X1 U745 ( .A(G128), .B(n676), .Z(G30) );
  NAND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n679), .B(G146), .ZN(G48) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U749 ( .A(KEYINPUT120), .B(n682), .Z(n683) );
  XNOR2_X1 U750 ( .A(G113), .B(n683), .ZN(G15) );
  XOR2_X1 U751 ( .A(G125), .B(KEYINPUT37), .Z(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(n684), .ZN(G27) );
  XNOR2_X1 U753 ( .A(G134), .B(n686), .ZN(G36) );
  NOR2_X1 U754 ( .A1(n357), .A2(n687), .ZN(n721) );
  NOR2_X1 U755 ( .A1(n689), .A2(n353), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT49), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n697) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U759 ( .A(KEYINPUT50), .B(n695), .Z(n696) );
  NOR2_X1 U760 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n698), .B(KEYINPUT121), .ZN(n701) );
  NAND2_X1 U762 ( .A1(n699), .A2(n562), .ZN(n700) );
  NAND2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U764 ( .A(KEYINPUT51), .B(n702), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n722), .A2(n703), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n706), .B(KEYINPUT122), .ZN(n707) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n714) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U773 ( .A(n717), .B(KEYINPUT52), .ZN(n718) );
  NOR2_X1 U774 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n722), .A2(n713), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(KEYINPUT123), .ZN(n724) );
  NAND2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n726), .A2(G953), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n727), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U781 ( .A1(G224), .A2(G953), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n728), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U783 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U784 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n732), .A2(n731), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n733), .B(KEYINPUT127), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n735), .B(n734), .ZN(n737) );
  NOR2_X1 U788 ( .A1(G898), .A2(n744), .ZN(n736) );
  NOR2_X1 U789 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n739), .B(n738), .ZN(G69) );
  XNOR2_X1 U791 ( .A(n741), .B(n740), .ZN(n746) );
  INV_X1 U792 ( .A(n746), .ZN(n743) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n750) );
  XNOR2_X1 U795 ( .A(G227), .B(n746), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U799 ( .A(G137), .B(n751), .Z(G39) );
  XOR2_X1 U800 ( .A(n752), .B(G131), .Z(G33) );
endmodule

