//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(G116), .B(G119), .Z(new_n193));
  OAI21_X1  g007(.A(KEYINPUT68), .B1(new_n193), .B2(new_n188), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(G107), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n197), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n196), .A2(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n199), .A2(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT5), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G116), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n191), .A2(KEYINPUT5), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n213), .A2(new_n214), .A3(G113), .A4(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n195), .A2(new_n208), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G110), .B(G122), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n197), .A2(new_n200), .A3(new_n202), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G101), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n192), .A2(new_n194), .B1(new_n193), .B2(new_n188), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n217), .B(new_n218), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT6), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n193), .A2(new_n188), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n195), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n223), .A3(new_n221), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n218), .B1(new_n230), .B2(new_n217), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n187), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n217), .B1(new_n224), .B2(new_n225), .ZN(new_n233));
  INV_X1    g047(.A(new_n218), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n235), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n226), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G125), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  AOI21_X1  g059(.A(G146), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n241), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n242), .A2(G146), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT64), .B(G143), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G146), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n249), .A2(KEYINPUT65), .B1(new_n239), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n254), .B(new_n241), .C1(new_n246), .C2(new_n248), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n238), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  OAI21_X1  g071(.A(G128), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n246), .B2(new_n248), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n243), .A2(new_n245), .A3(G146), .ZN(new_n260));
  INV_X1    g074(.A(new_n250), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G125), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G224), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G953), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n267), .B(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n231), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n237), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n256), .A2(new_n266), .B1(new_n276), .B2(new_n269), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n218), .B(KEYINPUT8), .ZN(new_n278));
  INV_X1    g092(.A(new_n217), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n208), .B1(new_n195), .B2(new_n216), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NOR4_X1   g096(.A1(new_n256), .A2(new_n276), .A3(new_n266), .A4(new_n269), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n275), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n270), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(KEYINPUT83), .A3(new_n281), .A4(new_n277), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n286), .A3(new_n226), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n274), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n274), .A2(new_n287), .A3(new_n288), .A4(new_n290), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G134), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n262), .A2(G143), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n243), .A2(new_n245), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n262), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT89), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n251), .A2(G128), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT89), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n296), .A4(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n305));
  INV_X1    g119(.A(G122), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G116), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G122), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n305), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n309), .A3(new_n305), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G107), .ZN(new_n313));
  INV_X1    g127(.A(new_n312), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n199), .B1(new_n314), .B2(new_n310), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n301), .A2(KEYINPUT13), .A3(new_n297), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT13), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n243), .A2(new_n245), .A3(new_n318), .A4(G128), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n319), .A2(G134), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n304), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT90), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n313), .A2(new_n315), .B1(new_n317), .B2(new_n320), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n304), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n315), .A2(KEYINPUT91), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n301), .A2(new_n297), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n299), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n308), .A2(KEYINPUT14), .A3(G122), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n307), .A2(new_n309), .ZN(new_n333));
  OAI211_X1 g147(.A(G107), .B(new_n332), .C1(new_n333), .C2(KEYINPUT14), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n315), .A2(KEYINPUT91), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n328), .A2(new_n331), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT9), .B(G234), .ZN(new_n337));
  INV_X1    g151(.A(G217), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n337), .A2(new_n338), .A3(G953), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n327), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n327), .B2(new_n336), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n288), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G478), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(KEYINPUT15), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(KEYINPUT92), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT92), .ZN(new_n347));
  INV_X1    g161(.A(new_n326), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n325), .B1(new_n324), .B2(new_n304), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n336), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n339), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n352), .B2(new_n340), .ZN(new_n353));
  INV_X1    g167(.A(new_n345), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n346), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n288), .B(new_n354), .C1(new_n341), .C2(new_n342), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(KEYINPUT93), .A3(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G475), .A2(G902), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n362), .B(KEYINPUT87), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(KEYINPUT66), .A2(G131), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT66), .A2(G131), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G237), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT71), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT71), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G237), .ZN(new_n372));
  AOI21_X1  g186(.A(G953), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(G143), .A3(G214), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n298), .B1(new_n373), .B2(G214), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n376), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n367), .A3(new_n374), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT17), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n238), .B2(KEYINPUT75), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(G125), .A3(G140), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n238), .B2(G140), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n386), .A2(new_n247), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n247), .B1(new_n386), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n378), .A2(new_n374), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n368), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G113), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n196), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  INV_X1    g211(.A(G214), .ZN(new_n398));
  AOI211_X1 g212(.A(new_n398), .B(G953), .C1(new_n370), .C2(new_n372), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n374), .B(new_n397), .C1(new_n399), .C2(new_n298), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n378), .A2(KEYINPUT85), .A3(new_n397), .A4(new_n374), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n397), .ZN(new_n405));
  XOR2_X1   g219(.A(G125), .B(G140), .Z(new_n406));
  OR2_X1    g220(.A1(new_n406), .A2(G146), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n383), .A2(G146), .A3(new_n385), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n392), .A2(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n394), .A2(new_n396), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n377), .A2(new_n379), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n383), .A2(KEYINPUT19), .A3(new_n385), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(new_n414), .C1(new_n406), .C2(KEYINPUT19), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n414), .B2(new_n413), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n390), .B1(new_n416), .B2(new_n247), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n396), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n364), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n410), .A2(new_n418), .ZN(new_n424));
  INV_X1    g238(.A(new_n396), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n394), .A2(new_n410), .A3(new_n396), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n364), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n396), .B1(new_n394), .B2(new_n410), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n288), .B1(new_n411), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n423), .A2(new_n430), .B1(G475), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n356), .A2(new_n361), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT78), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(KEYINPUT79), .Z(new_n437));
  INV_X1    g251(.A(G953), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n438), .A2(G952), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(G902), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(G898), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR4_X1   g260(.A1(new_n295), .A2(new_n434), .A3(new_n437), .A4(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G140), .ZN(new_n448));
  INV_X1    g262(.A(G227), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(G953), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n448), .B(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT10), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n264), .B2(new_n259), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G128), .B1(new_n246), .B2(new_n257), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n260), .A2(new_n261), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n207), .B1(new_n457), .B2(new_n264), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n458), .B2(KEYINPUT10), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n253), .A2(new_n255), .A3(new_n223), .A4(new_n221), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT11), .B1(new_n296), .B2(G137), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT11), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(G134), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n296), .A2(G137), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n367), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G131), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n462), .A2(new_n465), .B1(new_n296), .B2(G137), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n459), .A2(new_n461), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n252), .B1(G128), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n208), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT10), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n453), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n473), .B1(new_n479), .B2(new_n460), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n451), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n451), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n473), .A3(new_n460), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n259), .A2(new_n207), .A3(new_n264), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT77), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n458), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n259), .A2(new_n207), .A3(new_n488), .A4(new_n264), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n471), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n476), .B1(new_n456), .B2(new_n455), .ZN(new_n492));
  OAI211_X1 g306(.A(KEYINPUT77), .B(new_n484), .C1(new_n492), .C2(new_n207), .ZN(new_n493));
  INV_X1    g307(.A(new_n490), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT12), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n482), .B(new_n483), .C1(new_n491), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n481), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G469), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n288), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n288), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n471), .B1(new_n459), .B2(new_n461), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n482), .A3(new_n483), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n459), .A2(new_n461), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n487), .B1(new_n486), .B2(new_n490), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT12), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n473), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(G469), .B(new_n503), .C1(new_n507), .C2(new_n482), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G221), .B1(new_n337), .B2(G902), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n447), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT32), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n464), .B2(G134), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n464), .A2(G134), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n296), .A2(KEYINPUT67), .A3(G137), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n468), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n468), .A2(new_n520), .A3(KEYINPUT69), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n265), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n248), .B1(new_n298), .B2(new_n247), .ZN(new_n526));
  INV_X1    g340(.A(new_n241), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT65), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n252), .A2(new_n239), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n471), .A2(new_n528), .A3(new_n255), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(KEYINPUT30), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT70), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n525), .A2(KEYINPUT70), .A3(new_n530), .A4(KEYINPUT30), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n265), .A2(new_n468), .A3(new_n520), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n225), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT31), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n373), .A2(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT27), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n525), .A2(new_n530), .A3(new_n225), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n541), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(KEYINPUT28), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n525), .A2(new_n551), .A3(new_n530), .A4(new_n225), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n537), .A2(new_n229), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n545), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT72), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n547), .B1(new_n535), .B2(new_n539), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n559), .B1(new_n560), .B2(new_n541), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n537), .A2(new_n538), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n229), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n533), .B2(new_n534), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT72), .B(KEYINPUT31), .C1(new_n564), .C2(new_n547), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n558), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n514), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n546), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n535), .B2(new_n539), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT73), .B1(new_n571), .B2(new_n545), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n573), .B(new_n556), .C1(new_n564), .C2(new_n570), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n550), .A2(new_n552), .B1(new_n229), .B2(new_n537), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT29), .B1(new_n575), .B2(new_n545), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n525), .A2(new_n530), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n229), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n553), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n545), .A2(KEYINPUT29), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n565), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n549), .A2(new_n557), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n567), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n569), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT74), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n569), .A2(new_n584), .A3(new_n588), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n338), .B1(G234), .B2(new_n288), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT25), .ZN(new_n596));
  INV_X1    g410(.A(new_n390), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT23), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n210), .B2(G128), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n599), .B(new_n600), .C1(G119), .C2(new_n262), .ZN(new_n601));
  XNOR2_X1  g415(.A(G119), .B(G128), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT24), .B(G110), .Z(new_n603));
  OAI22_X1  g417(.A1(new_n601), .A2(G110), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n597), .A2(new_n604), .A3(new_n407), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n601), .A2(G110), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n389), .B2(new_n390), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT22), .B(G137), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n438), .A2(G221), .A3(G234), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n605), .A2(new_n607), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n596), .B1(new_n615), .B2(G902), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n613), .A2(KEYINPUT25), .A3(new_n288), .A4(new_n614), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n595), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n615), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n594), .A2(G902), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n593), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT76), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n593), .A2(KEYINPUT76), .A3(new_n621), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n513), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n201), .ZN(G3));
  AOI21_X1  g441(.A(G902), .B1(new_n585), .B2(new_n586), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(KEYINPUT94), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n628), .B(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n621), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n511), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT95), .Z(new_n635));
  INV_X1    g449(.A(new_n436), .ZN(new_n636));
  INV_X1    g450(.A(new_n446), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n294), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n352), .A2(new_n340), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n350), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT33), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n352), .A2(new_n641), .A3(KEYINPUT33), .A4(new_n340), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n344), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n344), .A2(new_n288), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n343), .B2(G478), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n638), .A2(new_n433), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n635), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  NAND3_X1  g468(.A1(new_n428), .A2(new_n421), .A3(new_n364), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n423), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n423), .A2(KEYINPUT97), .A3(new_n655), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n658), .A2(new_n659), .B1(G475), .B2(new_n432), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n356), .A2(new_n361), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n638), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n635), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n612), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n608), .B(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(new_n620), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n618), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n511), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n447), .A2(new_n631), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AOI21_X1  g488(.A(new_n436), .B1(new_n292), .B2(new_n293), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n444), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n441), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n676), .A2(new_n662), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n593), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  AOI21_X1  g497(.A(new_n433), .B1(new_n356), .B2(new_n361), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n636), .A3(new_n670), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n679), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n512), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n685), .B1(KEYINPUT40), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n545), .B1(new_n579), .B2(new_n546), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n288), .B1(new_n560), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G472), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n568), .B1(new_n585), .B2(new_n586), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(KEYINPUT32), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n566), .A2(new_n514), .A3(new_n568), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n294), .B(KEYINPUT38), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n690), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n298), .ZN(G45));
  NOR4_X1   g515(.A1(new_n433), .A2(new_n645), .A3(new_n648), .A4(new_n680), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n671), .A2(new_n702), .A3(new_n675), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n587), .A2(new_n567), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n704), .A2(new_n514), .B1(G472), .B2(new_n583), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n591), .B1(new_n705), .B2(new_n588), .ZN(new_n706));
  INV_X1    g520(.A(new_n592), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  INV_X1    g523(.A(new_n510), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n497), .A2(new_n288), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT99), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n499), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n711), .A2(KEYINPUT99), .A3(G469), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT100), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(new_n593), .A3(new_n651), .A4(new_n621), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n593), .A3(new_n621), .A4(new_n663), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND2_X1  g540(.A1(new_n716), .A2(new_n675), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n434), .A2(new_n446), .A3(new_n670), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n593), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT101), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n556), .B1(new_n580), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n553), .A2(new_n732), .A3(new_n579), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n560), .B(new_n541), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n567), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(new_n621), .C1(new_n628), .C2(new_n629), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n684), .A2(new_n675), .A3(new_n637), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n718), .A2(new_n739), .A3(new_n740), .A4(new_n720), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  OAI21_X1  g556(.A(G472), .B1(new_n566), .B2(G902), .ZN(new_n743));
  INV_X1    g557(.A(new_n670), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n702), .A2(new_n743), .A3(new_n744), .A4(new_n737), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n727), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n238), .ZN(G27));
  NAND2_X1  g561(.A1(new_n696), .A2(KEYINPUT103), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n588), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n705), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n621), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n294), .A2(new_n436), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT102), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n511), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n509), .A2(KEYINPUT102), .A3(new_n510), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n702), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT42), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n650), .A2(KEYINPUT42), .A3(new_n433), .A4(new_n680), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n593), .A2(new_n758), .A3(new_n621), .A4(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NOR2_X1   g578(.A1(new_n662), .A2(new_n680), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n593), .A2(new_n758), .A3(new_n621), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT104), .B(G134), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G36));
  NAND2_X1  g582(.A1(new_n649), .A2(new_n433), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n744), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n772), .A2(new_n773), .A3(new_n631), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n772), .B2(new_n631), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n753), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT105), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n472), .A2(new_n480), .A3(new_n451), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n483), .B1(new_n491), .B2(new_n495), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n451), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n784), .B2(new_n501), .ZN(new_n785));
  AOI211_X1 g599(.A(G469), .B(G902), .C1(new_n481), .C2(new_n496), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n501), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n710), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n687), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n774), .A2(KEYINPUT105), .A3(new_n775), .A4(new_n753), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n778), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  OR2_X1    g607(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n753), .A2(new_n702), .A3(new_n632), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n593), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n442), .A2(new_n771), .A3(new_n716), .A4(new_n753), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n744), .A3(new_n743), .A4(new_n737), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n753), .A2(new_n716), .A3(new_n621), .A4(new_n442), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n698), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n433), .A3(new_n650), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n801), .B1(new_n808), .B2(KEYINPUT110), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(KEYINPUT110), .B2(new_n808), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n771), .A2(new_n442), .A3(new_n739), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n699), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n716), .A2(new_n436), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT109), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n714), .A2(new_n715), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n796), .B1(new_n710), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n753), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n811), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n817), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n810), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n801), .B1(new_n822), .B2(new_n807), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n423), .A2(new_n430), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n432), .A2(G475), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n805), .A2(new_n827), .A3(new_n649), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n828), .B(new_n439), .C1(new_n727), .C2(new_n811), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n802), .A2(new_n621), .A3(new_n751), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT48), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT48), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n823), .A2(new_n824), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT111), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n823), .A2(new_n836), .A3(new_n824), .A4(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n746), .B1(new_n593), .B2(new_n681), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n618), .A2(new_n669), .A3(new_n680), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n508), .A2(new_n501), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n510), .B(new_n842), .C1(new_n843), .C2(new_n786), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT107), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n509), .A2(KEYINPUT107), .A3(new_n510), .A4(new_n842), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n675), .A3(new_n684), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n697), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n593), .B2(new_n703), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n841), .A2(new_n850), .A3(KEYINPUT108), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT108), .B1(new_n841), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n840), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n746), .ZN(new_n854));
  INV_X1    g668(.A(new_n849), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n682), .A2(new_n708), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n827), .B1(new_n645), .B2(new_n648), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n434), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n446), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n295), .A2(new_n437), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n631), .A3(new_n862), .A4(new_n633), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n741), .A2(new_n672), .A3(new_n863), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n722), .A2(new_n864), .A3(new_n725), .A4(new_n730), .ZN(new_n865));
  INV_X1    g679(.A(new_n626), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n745), .A2(new_n757), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n661), .A2(new_n680), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n660), .A2(new_n753), .A3(new_n868), .A4(new_n671), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n593), .B2(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n760), .A2(new_n870), .A3(new_n762), .A4(new_n766), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n865), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n839), .B1(new_n858), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n864), .A2(new_n722), .A3(new_n725), .A4(new_n730), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n760), .A2(new_n870), .A3(new_n762), .A4(new_n766), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n626), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT108), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n856), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n841), .A2(new_n850), .A3(KEYINPUT108), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(KEYINPUT52), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n876), .A2(KEYINPUT53), .A3(new_n853), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT54), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n853), .A2(new_n880), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n839), .B1(new_n884), .B2(new_n872), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n876), .A2(KEYINPUT53), .A3(new_n853), .A4(new_n857), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n838), .A2(new_n889), .B1(G952), .B2(G953), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n769), .A2(new_n632), .A3(new_n710), .A4(new_n437), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT49), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n818), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT106), .Z(new_n894));
  AOI21_X1  g708(.A(new_n699), .B1(new_n892), .B2(new_n818), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n697), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n890), .A2(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n438), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n288), .B1(new_n885), .B2(new_n887), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n237), .A2(new_n273), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n271), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n899), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n900), .A2(KEYINPUT113), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n900), .A2(KEYINPUT113), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n291), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n906), .B1(new_n910), .B2(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n500), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n886), .B1(new_n885), .B2(new_n887), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT115), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n888), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g732(.A(KEYINPUT115), .B(new_n886), .C1(new_n885), .C2(new_n887), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n497), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n907), .A2(new_n908), .A3(new_n784), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n898), .B1(new_n921), .B2(new_n922), .ZN(G54));
  NAND2_X1  g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n428), .B1(new_n909), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n428), .ZN(new_n927));
  NOR4_X1   g741(.A1(new_n907), .A2(new_n908), .A3(new_n927), .A4(new_n924), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n928), .A3(new_n898), .ZN(G60));
  INV_X1    g743(.A(new_n643), .ZN(new_n930));
  INV_X1    g744(.A(new_n644), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n646), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n918), .B2(new_n919), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n899), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n936), .B2(new_n899), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n932), .B1(new_n889), .B2(new_n934), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G63));
  OAI21_X1  g755(.A(new_n899), .B1(KEYINPUT119), .B2(KEYINPUT61), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n943));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n885), .B2(new_n887), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n946), .B2(new_n668), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n619), .B2(new_n946), .ZN(new_n948));
  NAND2_X1  g762(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n445), .B2(new_n268), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n865), .A2(new_n866), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT120), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n902), .B1(G898), .B2(new_n438), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  NAND2_X1  g770(.A1(new_n792), .A2(new_n799), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n789), .A2(new_n675), .A3(new_n687), .A4(new_n684), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n959), .A2(KEYINPUT121), .A3(new_n752), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n841), .A2(new_n708), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT121), .B1(new_n959), .B2(new_n752), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n766), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n958), .A2(KEYINPUT122), .A3(new_n763), .A4(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n763), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n957), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n967), .A3(new_n438), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n535), .A2(new_n562), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(new_n416), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n624), .A2(new_n625), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n820), .A2(new_n688), .A3(new_n860), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n792), .A2(new_n799), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n961), .A2(new_n700), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT62), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(G953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n449), .B2(new_n677), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT123), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n981), .B(new_n983), .ZN(G72));
  NAND3_X1  g798(.A1(new_n964), .A2(new_n967), .A3(new_n953), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n571), .B(KEYINPUT125), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n545), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n898), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n979), .A2(new_n953), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n987), .ZN(new_n994));
  INV_X1    g808(.A(new_n987), .ZN(new_n995));
  AOI211_X1 g809(.A(KEYINPUT124), .B(new_n995), .C1(new_n979), .C2(new_n953), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n545), .B(new_n989), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n572), .A2(new_n574), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n987), .B1(new_n998), .B2(new_n560), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT126), .Z(new_n1000));
  AOI211_X1 g814(.A(KEYINPUT127), .B(new_n1000), .C1(new_n873), .C2(new_n881), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1000), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n882), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n991), .B(new_n997), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(G57));
endmodule


