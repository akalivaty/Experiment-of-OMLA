

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(KEYINPUT15), .B(n591), .Z(n924) );
  NAND2_X2 U552 ( .A1(n603), .A2(n726), .ZN(n664) );
  XNOR2_X2 U553 ( .A(n672), .B(KEYINPUT32), .ZN(n694) );
  NOR2_X1 U554 ( .A1(n652), .A2(n677), .ZN(n654) );
  XNOR2_X1 U555 ( .A(KEYINPUT108), .B(n759), .ZN(n518) );
  AND2_X1 U556 ( .A1(n600), .A2(n726), .ZN(n602) );
  NOR2_X1 U557 ( .A1(n617), .A2(n933), .ZN(n619) );
  INV_X1 U558 ( .A(KEYINPUT30), .ZN(n653) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n643) );
  AND2_X1 U560 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U561 ( .A(KEYINPUT1), .B(n525), .Z(n788) );
  NAND2_X1 U562 ( .A1(n760), .A2(n518), .ZN(n761) );
  NOR2_X1 U563 ( .A1(n546), .A2(n545), .ZN(G164) );
  NOR2_X1 U564 ( .A1(G651), .A2(G543), .ZN(n791) );
  NAND2_X1 U565 ( .A1(n791), .A2(G89), .ZN(n519) );
  XNOR2_X1 U566 ( .A(n519), .B(KEYINPUT4), .ZN(n522) );
  INV_X1 U567 ( .A(G651), .ZN(n524) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n566) );
  OR2_X1 U569 ( .A1(n524), .A2(n566), .ZN(n520) );
  XNOR2_X2 U570 ( .A(KEYINPUT67), .B(n520), .ZN(n787) );
  NAND2_X1 U571 ( .A1(G76), .A2(n787), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT5), .ZN(n531) );
  NOR2_X1 U574 ( .A1(G543), .A2(n524), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n788), .A2(G63), .ZN(n526) );
  XNOR2_X1 U576 ( .A(n526), .B(KEYINPUT72), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G651), .A2(n566), .ZN(n792) );
  NAND2_X1 U578 ( .A1(G51), .A2(n792), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U582 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U584 ( .A(G2104), .ZN(n541) );
  NOR2_X2 U585 ( .A1(G2105), .A2(n541), .ZN(n887) );
  NAND2_X1 U586 ( .A1(n887), .A2(G102), .ZN(n533) );
  XNOR2_X1 U587 ( .A(n533), .B(KEYINPUT88), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XOR2_X2 U589 ( .A(KEYINPUT17), .B(n534), .Z(n886) );
  NAND2_X1 U590 ( .A1(G138), .A2(n886), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n538) );
  INV_X1 U592 ( .A(KEYINPUT89), .ZN(n537) );
  XNOR2_X1 U593 ( .A(n538), .B(n537), .ZN(n546) );
  INV_X1 U594 ( .A(G2105), .ZN(n540) );
  NOR2_X1 U595 ( .A1(G2104), .A2(n540), .ZN(n882) );
  NAND2_X1 U596 ( .A1(G126), .A2(n882), .ZN(n539) );
  XNOR2_X1 U597 ( .A(n539), .B(KEYINPUT86), .ZN(n544) );
  NOR2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n883) );
  NAND2_X1 U599 ( .A1(G114), .A2(n883), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT87), .B(n542), .Z(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n791), .A2(G90), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n787), .A2(G77), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n549), .Z(n552) );
  NAND2_X1 U606 ( .A1(G64), .A2(n788), .ZN(n550) );
  XOR2_X1 U607 ( .A(KEYINPUT68), .B(n550), .Z(n551) );
  NOR2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n792), .A2(G52), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(G301) );
  INV_X1 U611 ( .A(G301), .ZN(G171) );
  NAND2_X1 U612 ( .A1(G62), .A2(n788), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G75), .A2(n787), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G88), .A2(n791), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G50), .A2(n792), .ZN(n557) );
  XNOR2_X1 U617 ( .A(KEYINPUT79), .B(n557), .ZN(n558) );
  NOR2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n562), .B(KEYINPUT80), .ZN(G303) );
  NAND2_X1 U621 ( .A1(G49), .A2(n792), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G74), .A2(G651), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U624 ( .A1(n788), .A2(n565), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n566), .A2(G87), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(G288) );
  NAND2_X1 U627 ( .A1(G86), .A2(n791), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G61), .A2(n788), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G73), .A2(n787), .ZN(n571) );
  XNOR2_X1 U631 ( .A(n571), .B(KEYINPUT2), .ZN(n572) );
  XNOR2_X1 U632 ( .A(n572), .B(KEYINPUT77), .ZN(n573) );
  NOR2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U634 ( .A(n575), .B(KEYINPUT78), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G48), .A2(n792), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(G305) );
  NAND2_X1 U637 ( .A1(G72), .A2(n787), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G60), .A2(n788), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G85), .A2(n791), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G47), .A2(n792), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(G290) );
  NAND2_X1 U644 ( .A1(G79), .A2(n787), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G54), .A2(n792), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G92), .A2(n791), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G66), .A2(n788), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U650 ( .A(KEYINPUT71), .B(n588), .Z(n589) );
  NOR2_X1 U651 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G125), .A2(n882), .ZN(n592) );
  XOR2_X1 U653 ( .A(KEYINPUT65), .B(n592), .Z(n762) );
  AND2_X1 U654 ( .A1(G40), .A2(n762), .ZN(n599) );
  NAND2_X1 U655 ( .A1(G101), .A2(n887), .ZN(n593) );
  XOR2_X1 U656 ( .A(n593), .B(KEYINPUT23), .Z(n596) );
  NAND2_X1 U657 ( .A1(G137), .A2(n886), .ZN(n594) );
  XNOR2_X1 U658 ( .A(KEYINPUT66), .B(n594), .ZN(n595) );
  AND2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U660 ( .A1(n883), .A2(G113), .ZN(n597) );
  AND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n763) );
  NAND2_X1 U662 ( .A1(n599), .A2(n763), .ZN(n725) );
  INV_X1 U663 ( .A(G1996), .ZN(n746) );
  NOR2_X1 U664 ( .A1(n725), .A2(n746), .ZN(n600) );
  NOR2_X2 U665 ( .A1(G164), .A2(G1384), .ZN(n726) );
  XOR2_X1 U666 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n601) );
  XNOR2_X1 U667 ( .A(n602), .B(n601), .ZN(n605) );
  INV_X1 U668 ( .A(n725), .ZN(n603) );
  NAND2_X1 U669 ( .A1(n664), .A2(G1341), .ZN(n604) );
  NAND2_X1 U670 ( .A1(n605), .A2(n604), .ZN(n617) );
  NAND2_X1 U671 ( .A1(G56), .A2(n788), .ZN(n606) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n606), .Z(n614) );
  NAND2_X1 U673 ( .A1(n787), .A2(G68), .ZN(n607) );
  XNOR2_X1 U674 ( .A(n607), .B(KEYINPUT70), .ZN(n611) );
  XOR2_X1 U675 ( .A(KEYINPUT69), .B(KEYINPUT12), .Z(n609) );
  NAND2_X1 U676 ( .A1(G81), .A2(n791), .ZN(n608) );
  XNOR2_X1 U677 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U678 ( .A(KEYINPUT13), .B(n612), .ZN(n613) );
  NOR2_X1 U679 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U680 ( .A1(n792), .A2(G43), .ZN(n615) );
  NAND2_X1 U681 ( .A1(n616), .A2(n615), .ZN(n933) );
  NOR2_X1 U682 ( .A1(n924), .A2(n619), .ZN(n618) );
  XNOR2_X1 U683 ( .A(KEYINPUT100), .B(n618), .ZN(n627) );
  NAND2_X1 U684 ( .A1(n619), .A2(n924), .ZN(n624) );
  NAND2_X1 U685 ( .A1(n664), .A2(G1348), .ZN(n620) );
  XNOR2_X1 U686 ( .A(n620), .B(KEYINPUT98), .ZN(n622) );
  INV_X1 U687 ( .A(n664), .ZN(n646) );
  NAND2_X1 U688 ( .A1(n646), .A2(G2067), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U691 ( .A(n625), .B(KEYINPUT99), .ZN(n626) );
  OR2_X1 U692 ( .A1(n627), .A2(n626), .ZN(n638) );
  NAND2_X1 U693 ( .A1(G65), .A2(n788), .ZN(n629) );
  NAND2_X1 U694 ( .A1(G53), .A2(n792), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U696 ( .A1(G78), .A2(n787), .ZN(n631) );
  NAND2_X1 U697 ( .A1(G91), .A2(n791), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U699 ( .A1(n633), .A2(n632), .ZN(n803) );
  NAND2_X1 U700 ( .A1(n646), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U701 ( .A(n634), .B(KEYINPUT27), .ZN(n636) );
  INV_X1 U702 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U703 ( .A1(n998), .A2(n646), .ZN(n635) );
  NOR2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U705 ( .A1(n803), .A2(n639), .ZN(n637) );
  NAND2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U707 ( .A1(n803), .A2(n639), .ZN(n640) );
  XOR2_X1 U708 ( .A(n640), .B(KEYINPUT28), .Z(n641) );
  NAND2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n644) );
  XNOR2_X1 U710 ( .A(n644), .B(n643), .ZN(n650) );
  OR2_X1 U711 ( .A1(n646), .A2(G1961), .ZN(n648) );
  XOR2_X1 U712 ( .A(G2078), .B(KEYINPUT25), .Z(n645) );
  XNOR2_X1 U713 ( .A(KEYINPUT97), .B(n645), .ZN(n949) );
  NAND2_X1 U714 ( .A1(n646), .A2(n949), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n657) );
  NAND2_X1 U716 ( .A1(n657), .A2(G171), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n663) );
  XNOR2_X1 U718 ( .A(KEYINPUT102), .B(KEYINPUT31), .ZN(n661) );
  NOR2_X1 U719 ( .A1(n664), .A2(G2084), .ZN(n651) );
  XOR2_X1 U720 ( .A(KEYINPUT96), .B(n651), .Z(n673) );
  NAND2_X1 U721 ( .A1(G8), .A2(n673), .ZN(n652) );
  NAND2_X1 U722 ( .A1(G8), .A2(n664), .ZN(n702) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n702), .ZN(n677) );
  XNOR2_X1 U724 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(G168), .A2(n655), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n656), .B(KEYINPUT101), .ZN(n659) );
  OR2_X1 U727 ( .A1(n657), .A2(G171), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n675) );
  NAND2_X1 U731 ( .A1(G286), .A2(n675), .ZN(n670) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n702), .ZN(n666) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U735 ( .A(KEYINPUT103), .B(n667), .Z(n668) );
  NAND2_X1 U736 ( .A1(n668), .A2(G303), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n671), .A2(G8), .ZN(n672) );
  INV_X1 U739 ( .A(n673), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n674), .A2(G8), .ZN(n679) );
  INV_X1 U741 ( .A(n675), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n695) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n928) );
  AND2_X1 U745 ( .A1(n695), .A2(n928), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n694), .A2(n680), .ZN(n684) );
  INV_X1 U747 ( .A(n928), .ZN(n682) );
  NOR2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U749 ( .A1(G303), .A2(G1971), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n687), .A2(n681), .ZN(n931) );
  OR2_X1 U751 ( .A1(n682), .A2(n931), .ZN(n683) );
  AND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n685), .A2(n702), .ZN(n686) );
  OR2_X1 U754 ( .A1(n686), .A2(KEYINPUT33), .ZN(n692) );
  XOR2_X1 U755 ( .A(G1981), .B(G305), .Z(n920) );
  INV_X1 U756 ( .A(n920), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n687), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U758 ( .A1(n702), .A2(n688), .ZN(n689) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n693), .B(KEYINPUT104), .ZN(n706) );
  NAND2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n698) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n696) );
  NAND2_X1 U764 ( .A1(G8), .A2(n696), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  AND2_X1 U766 ( .A1(n699), .A2(n702), .ZN(n704) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U768 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n742) );
  XOR2_X1 U772 ( .A(KEYINPUT90), .B(G1986), .Z(n707) );
  XNOR2_X1 U773 ( .A(G290), .B(n707), .ZN(n925) );
  NAND2_X1 U774 ( .A1(G95), .A2(n887), .ZN(n709) );
  NAND2_X1 U775 ( .A1(G119), .A2(n882), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U777 ( .A1(n883), .A2(G107), .ZN(n710) );
  XOR2_X1 U778 ( .A(KEYINPUT94), .B(n710), .Z(n711) );
  NOR2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U780 ( .A1(n886), .A2(G131), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n893) );
  NAND2_X1 U782 ( .A1(G1991), .A2(n893), .ZN(n715) );
  XNOR2_X1 U783 ( .A(n715), .B(KEYINPUT95), .ZN(n724) );
  NAND2_X1 U784 ( .A1(G105), .A2(n887), .ZN(n716) );
  XNOR2_X1 U785 ( .A(n716), .B(KEYINPUT38), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n886), .A2(G141), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U788 ( .A1(G129), .A2(n882), .ZN(n720) );
  NAND2_X1 U789 ( .A1(G117), .A2(n883), .ZN(n719) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U791 ( .A1(n722), .A2(n721), .ZN(n864) );
  NOR2_X1 U792 ( .A1(n746), .A2(n864), .ZN(n723) );
  NOR2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n977) );
  NAND2_X1 U794 ( .A1(n925), .A2(n977), .ZN(n727) );
  NOR2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n758) );
  NAND2_X1 U796 ( .A1(n727), .A2(n758), .ZN(n740) );
  NAND2_X1 U797 ( .A1(n883), .A2(G116), .ZN(n728) );
  XNOR2_X1 U798 ( .A(n728), .B(KEYINPUT92), .ZN(n730) );
  NAND2_X1 U799 ( .A1(G128), .A2(n882), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U801 ( .A(KEYINPUT35), .B(n731), .ZN(n737) );
  NAND2_X1 U802 ( .A1(n886), .A2(G140), .ZN(n732) );
  XOR2_X1 U803 ( .A(KEYINPUT91), .B(n732), .Z(n734) );
  NAND2_X1 U804 ( .A1(n887), .A2(G104), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U806 ( .A(KEYINPUT34), .B(n735), .Z(n736) );
  NAND2_X1 U807 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U808 ( .A(KEYINPUT36), .B(n738), .Z(n865) );
  XNOR2_X1 U809 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  OR2_X1 U810 ( .A1(n865), .A2(n744), .ZN(n739) );
  XNOR2_X1 U811 ( .A(n739), .B(KEYINPUT93), .ZN(n987) );
  NAND2_X1 U812 ( .A1(n987), .A2(n758), .ZN(n753) );
  NAND2_X1 U813 ( .A1(n740), .A2(n753), .ZN(n741) );
  NOR2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U815 ( .A(n743), .ZN(n760) );
  NAND2_X1 U816 ( .A1(n865), .A2(n744), .ZN(n745) );
  XNOR2_X1 U817 ( .A(n745), .B(KEYINPUT106), .ZN(n985) );
  AND2_X1 U818 ( .A1(n746), .A2(n864), .ZN(n967) );
  INV_X1 U819 ( .A(n977), .ZN(n750) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U821 ( .A1(G1991), .A2(n893), .ZN(n970) );
  NOR2_X1 U822 ( .A1(n747), .A2(n970), .ZN(n748) );
  XOR2_X1 U823 ( .A(KEYINPUT105), .B(n748), .Z(n749) );
  NOR2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U825 ( .A1(n967), .A2(n751), .ZN(n752) );
  XNOR2_X1 U826 ( .A(n752), .B(KEYINPUT39), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n985), .A2(n755), .ZN(n756) );
  XOR2_X1 U829 ( .A(KEYINPUT107), .B(n756), .Z(n757) );
  NAND2_X1 U830 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U831 ( .A(n761), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U832 ( .A1(n763), .A2(n762), .ZN(G160) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G57), .ZN(G237) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  INV_X1 U837 ( .A(n803), .ZN(G299) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n830) );
  NAND2_X1 U841 ( .A1(n830), .A2(G567), .ZN(n765) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n765), .Z(G234) );
  INV_X1 U843 ( .A(G860), .ZN(n798) );
  OR2_X1 U844 ( .A1(n933), .A2(n798), .ZN(G153) );
  NAND2_X1 U845 ( .A1(G868), .A2(G301), .ZN(n767) );
  OR2_X1 U846 ( .A1(n924), .A2(G868), .ZN(n766) );
  NAND2_X1 U847 ( .A1(n767), .A2(n766), .ZN(G284) );
  INV_X1 U848 ( .A(G868), .ZN(n810) );
  NOR2_X1 U849 ( .A1(G286), .A2(n810), .ZN(n769) );
  NOR2_X1 U850 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U851 ( .A1(n769), .A2(n768), .ZN(G297) );
  NAND2_X1 U852 ( .A1(n798), .A2(G559), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n770), .A2(n924), .ZN(n771) );
  XNOR2_X1 U854 ( .A(n771), .B(KEYINPUT16), .ZN(n772) );
  XOR2_X1 U855 ( .A(KEYINPUT73), .B(n772), .Z(G148) );
  NOR2_X1 U856 ( .A1(G868), .A2(n933), .ZN(n775) );
  NAND2_X1 U857 ( .A1(n924), .A2(G868), .ZN(n773) );
  NOR2_X1 U858 ( .A1(G559), .A2(n773), .ZN(n774) );
  NOR2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U860 ( .A(KEYINPUT74), .B(n776), .ZN(G282) );
  NAND2_X1 U861 ( .A1(G123), .A2(n882), .ZN(n777) );
  XNOR2_X1 U862 ( .A(n777), .B(KEYINPUT18), .ZN(n780) );
  NAND2_X1 U863 ( .A1(G111), .A2(n883), .ZN(n778) );
  XOR2_X1 U864 ( .A(KEYINPUT75), .B(n778), .Z(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n784) );
  NAND2_X1 U866 ( .A1(G135), .A2(n886), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G99), .A2(n887), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n969) );
  XNOR2_X1 U870 ( .A(G2096), .B(n969), .ZN(n786) );
  INV_X1 U871 ( .A(G2100), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G80), .A2(n787), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G67), .A2(n788), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n796) );
  NAND2_X1 U876 ( .A1(G93), .A2(n791), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G55), .A2(n792), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U879 ( .A1(n796), .A2(n795), .ZN(n811) );
  XNOR2_X1 U880 ( .A(n811), .B(KEYINPUT76), .ZN(n800) );
  NAND2_X1 U881 ( .A1(G559), .A2(n924), .ZN(n797) );
  XOR2_X1 U882 ( .A(n933), .B(n797), .Z(n807) );
  NAND2_X1 U883 ( .A1(n807), .A2(n798), .ZN(n799) );
  XNOR2_X1 U884 ( .A(n800), .B(n799), .ZN(G145) );
  XNOR2_X1 U885 ( .A(n811), .B(KEYINPUT19), .ZN(n801) );
  XNOR2_X1 U886 ( .A(G288), .B(n801), .ZN(n802) );
  XNOR2_X1 U887 ( .A(G290), .B(n802), .ZN(n805) );
  XNOR2_X1 U888 ( .A(n803), .B(G303), .ZN(n804) );
  XNOR2_X1 U889 ( .A(n805), .B(n804), .ZN(n806) );
  XOR2_X1 U890 ( .A(n806), .B(G305), .Z(n901) );
  XOR2_X1 U891 ( .A(n807), .B(n901), .Z(n808) );
  XNOR2_X1 U892 ( .A(KEYINPUT81), .B(n808), .ZN(n809) );
  NOR2_X1 U893 ( .A1(n810), .A2(n809), .ZN(n813) );
  NOR2_X1 U894 ( .A1(G868), .A2(n811), .ZN(n812) );
  NOR2_X1 U895 ( .A1(n813), .A2(n812), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2078), .A2(G2084), .ZN(n814) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n814), .Z(n815) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n815), .ZN(n816) );
  XNOR2_X1 U899 ( .A(n816), .B(KEYINPUT83), .ZN(n818) );
  XOR2_X1 U900 ( .A(KEYINPUT21), .B(KEYINPUT82), .Z(n817) );
  XNOR2_X1 U901 ( .A(n818), .B(n817), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U904 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U905 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U906 ( .A1(G218), .A2(n821), .ZN(n822) );
  XNOR2_X1 U907 ( .A(KEYINPUT84), .B(n822), .ZN(n823) );
  NAND2_X1 U908 ( .A1(n823), .A2(G96), .ZN(n834) );
  NAND2_X1 U909 ( .A1(n834), .A2(G2106), .ZN(n827) );
  NAND2_X1 U910 ( .A1(G69), .A2(G120), .ZN(n824) );
  NOR2_X1 U911 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U912 ( .A1(G108), .A2(n825), .ZN(n835) );
  NAND2_X1 U913 ( .A1(n835), .A2(G567), .ZN(n826) );
  NAND2_X1 U914 ( .A1(n827), .A2(n826), .ZN(n836) );
  NAND2_X1 U915 ( .A1(G483), .A2(G661), .ZN(n828) );
  NOR2_X1 U916 ( .A1(n836), .A2(n828), .ZN(n829) );
  XOR2_X1 U917 ( .A(KEYINPUT85), .B(n829), .Z(n833) );
  NAND2_X1 U918 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U921 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  INV_X1 U930 ( .A(n836), .ZN(G319) );
  XOR2_X1 U931 ( .A(G2096), .B(KEYINPUT43), .Z(n838) );
  XNOR2_X1 U932 ( .A(G2090), .B(KEYINPUT110), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U934 ( .A(n839), .B(G2678), .Z(n841) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2100), .Z(n843) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1986), .B(G1956), .Z(n847) );
  XNOR2_X1 U942 ( .A(G1966), .B(G1961), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U944 ( .A(G1991), .B(G1976), .Z(n849) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1971), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U947 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U948 ( .A(KEYINPUT111), .B(G2474), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U950 ( .A(G1981), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U952 ( .A1(G100), .A2(n887), .ZN(n857) );
  NAND2_X1 U953 ( .A1(G112), .A2(n883), .ZN(n856) );
  NAND2_X1 U954 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT112), .B(n858), .ZN(n863) );
  NAND2_X1 U956 ( .A1(G124), .A2(n882), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U958 ( .A1(n886), .A2(G136), .ZN(n860) );
  NAND2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U960 ( .A1(n863), .A2(n862), .ZN(G162) );
  XOR2_X1 U961 ( .A(G162), .B(n864), .Z(n867) );
  XOR2_X1 U962 ( .A(G164), .B(n865), .Z(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n869) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U967 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U968 ( .A(G160), .B(n969), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n873), .B(n872), .ZN(n897) );
  NAND2_X1 U970 ( .A1(G139), .A2(n886), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G103), .A2(n887), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U973 ( .A1(G127), .A2(n882), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G115), .A2(n883), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U976 ( .A(KEYINPUT47), .B(n878), .ZN(n879) );
  XNOR2_X1 U977 ( .A(KEYINPUT113), .B(n879), .ZN(n880) );
  NOR2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n978) );
  NAND2_X1 U979 ( .A1(G130), .A2(n882), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G118), .A2(n883), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U982 ( .A1(G142), .A2(n886), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G106), .A2(n887), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U985 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n978), .B(n895), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U990 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n933), .B(G286), .ZN(n900) );
  XNOR2_X1 U992 ( .A(G171), .B(n924), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U995 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U996 ( .A(G2454), .B(G2435), .Z(n905) );
  XNOR2_X1 U997 ( .A(G2438), .B(G2427), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n912) );
  XOR2_X1 U999 ( .A(KEYINPUT109), .B(G2446), .Z(n907) );
  XNOR2_X1 U1000 ( .A(G2443), .B(G2430), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1002 ( .A(n908), .B(G2451), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G1348), .B(G1341), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n919), .ZN(G401) );
  XNOR2_X1 U1016 ( .A(KEYINPUT56), .B(G16), .ZN(n944) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G168), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(n922), .B(KEYINPUT121), .ZN(n923) );
  XOR2_X1 U1020 ( .A(KEYINPUT57), .B(n923), .Z(n942) );
  XNOR2_X1 U1021 ( .A(G1348), .B(n924), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n939) );
  NAND2_X1 U1023 ( .A1(G303), .A2(G1971), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(G1956), .B(G299), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(G171), .B(G1961), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(G1341), .B(n933), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT122), .B(n940), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n996) );
  XOR2_X1 U1036 ( .A(G29), .B(KEYINPUT120), .Z(n964) );
  XOR2_X1 U1037 ( .A(G2084), .B(G34), .Z(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT54), .B(n945), .ZN(n960) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n958) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n953) );
  XOR2_X1 U1045 ( .A(n949), .B(G27), .Z(n951) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(n961), .B(KEYINPUT119), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n989) );
  XOR2_X1 U1055 ( .A(n962), .B(n989), .Z(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n965), .ZN(n994) );
  XOR2_X1 U1058 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1060 ( .A(KEYINPUT51), .B(n968), .Z(n972) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1063 ( .A(G2084), .B(G160), .Z(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT116), .B(n973), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n983) );
  XOR2_X1 U1067 ( .A(G2072), .B(n978), .Z(n980) );
  XOR2_X1 U1068 ( .A(G164), .B(G2078), .Z(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1070 ( .A(KEYINPUT50), .B(n981), .Z(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1073 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1074 ( .A(KEYINPUT52), .B(n988), .ZN(n990) );
  NAND2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1076 ( .A1(n991), .A2(G29), .ZN(n992) );
  XOR2_X1 U1077 ( .A(KEYINPUT118), .B(n992), .Z(n993) );
  NOR2_X1 U1078 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1079 ( .A1(n996), .A2(n995), .ZN(n1025) );
  XOR2_X1 U1080 ( .A(G1966), .B(G21), .Z(n1009) );
  XOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .Z(n997) );
  XNOR2_X1 U1082 ( .A(G4), .B(n997), .ZN(n1006) );
  XNOR2_X1 U1083 ( .A(G20), .B(n998), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(n999), .B(KEYINPUT123), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(G6), .B(G1981), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1089 ( .A(KEYINPUT124), .B(n1004), .Z(n1005) );
  NOR2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(n1007), .B(KEYINPUT60), .ZN(n1008) );
  NAND2_X1 U1092 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(n1010), .B(KEYINPUT125), .ZN(n1018) );
  XOR2_X1 U1094 ( .A(G1971), .B(KEYINPUT126), .Z(n1011) );
  XNOR2_X1 U1095 ( .A(G22), .B(n1011), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(G1976), .B(G23), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G1986), .B(G24), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1016), .Z(n1017) );
  NAND2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(G5), .B(G1961), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1021), .Z(n1022) );
  NOR2_X1 U1105 ( .A1(G16), .A2(n1022), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT127), .B(n1023), .Z(n1024) );
  NOR2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1026), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
  INV_X1 U1110 ( .A(G303), .ZN(G166) );
endmodule

