

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U547 ( .A1(n725), .A2(n510), .ZN(n726) );
  NAND2_X1 U548 ( .A1(G8), .A2(n706), .ZN(n764) );
  INV_X1 U549 ( .A(KEYINPUT31), .ZN(n697) );
  NOR2_X1 U550 ( .A1(G1966), .A2(n764), .ZN(n739) );
  INV_X1 U551 ( .A(n892), .ZN(n746) );
  XNOR2_X1 U552 ( .A(n761), .B(KEYINPUT103), .ZN(n765) );
  NOR2_X2 U553 ( .A1(n532), .A2(n531), .ZN(G160) );
  AND2_X1 U554 ( .A1(G171), .A2(n724), .ZN(n510) );
  XOR2_X1 U555 ( .A(KEYINPUT74), .B(n568), .Z(n511) );
  OR2_X1 U556 ( .A1(n764), .A2(n763), .ZN(n512) );
  AND2_X1 U557 ( .A1(n748), .A2(n747), .ZN(n749) );
  AND2_X1 U558 ( .A1(n765), .A2(n512), .ZN(n799) );
  INV_X1 U559 ( .A(G651), .ZN(n537) );
  NOR2_X1 U560 ( .A1(G651), .A2(n654), .ZN(n650) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n640) );
  NOR2_X2 U562 ( .A1(G2105), .A2(n519), .ZN(n976) );
  NOR2_X1 U563 ( .A1(n524), .A2(n523), .ZN(G164) );
  INV_X1 U564 ( .A(KEYINPUT93), .ZN(n518) );
  INV_X1 U565 ( .A(G2104), .ZN(n519) );
  INV_X1 U566 ( .A(G2105), .ZN(n513) );
  NOR2_X1 U567 ( .A1(n519), .A2(n513), .ZN(n972) );
  NAND2_X1 U568 ( .A1(n972), .A2(G114), .ZN(n516) );
  NOR2_X1 U569 ( .A1(n513), .A2(G2104), .ZN(n514) );
  XNOR2_X2 U570 ( .A(n514), .B(KEYINPUT64), .ZN(n973) );
  NAND2_X1 U571 ( .A1(G126), .A2(n973), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U573 ( .A(n518), .B(n517), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G102), .A2(n976), .ZN(n522) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X1 U576 ( .A(KEYINPUT17), .B(n520), .Z(n977) );
  NAND2_X1 U577 ( .A1(G138), .A2(n977), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U579 ( .A1(G101), .A2(n976), .ZN(n525) );
  XNOR2_X1 U580 ( .A(n525), .B(KEYINPUT65), .ZN(n526) );
  XNOR2_X1 U581 ( .A(n526), .B(KEYINPUT23), .ZN(n528) );
  NAND2_X1 U582 ( .A1(G113), .A2(n972), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n977), .A2(G137), .ZN(n530) );
  NAND2_X1 U585 ( .A1(G125), .A2(n973), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n654) );
  NAND2_X1 U588 ( .A1(n650), .A2(G52), .ZN(n536) );
  NOR2_X1 U589 ( .A1(G543), .A2(n537), .ZN(n533) );
  XOR2_X1 U590 ( .A(KEYINPUT68), .B(n533), .Z(n534) );
  XNOR2_X2 U591 ( .A(KEYINPUT1), .B(n534), .ZN(n657) );
  NAND2_X1 U592 ( .A1(G64), .A2(n657), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n544) );
  OR2_X1 U594 ( .A1(n537), .A2(n654), .ZN(n538) );
  XNOR2_X1 U595 ( .A(KEYINPUT67), .B(n538), .ZN(n643) );
  NAND2_X1 U596 ( .A1(n643), .A2(G77), .ZN(n539) );
  XNOR2_X1 U597 ( .A(n539), .B(KEYINPUT70), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G90), .A2(n640), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n542), .Z(n543) );
  NOR2_X1 U601 ( .A1(n544), .A2(n543), .ZN(G171) );
  XOR2_X1 U602 ( .A(G2443), .B(G2446), .Z(n546) );
  XNOR2_X1 U603 ( .A(G2427), .B(G2451), .ZN(n545) );
  XNOR2_X1 U604 ( .A(n546), .B(n545), .ZN(n552) );
  XOR2_X1 U605 ( .A(G2430), .B(G2454), .Z(n548) );
  XNOR2_X1 U606 ( .A(G1341), .B(G1348), .ZN(n547) );
  XNOR2_X1 U607 ( .A(n548), .B(n547), .ZN(n550) );
  XOR2_X1 U608 ( .A(G2435), .B(G2438), .Z(n549) );
  XNOR2_X1 U609 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U610 ( .A(n552), .B(n551), .Z(n553) );
  AND2_X1 U611 ( .A1(G14), .A2(n553), .ZN(G401) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G69), .ZN(G235) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U616 ( .A(G223), .ZN(n818) );
  NAND2_X1 U617 ( .A1(n818), .A2(G567), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  XOR2_X1 U619 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n557) );
  NAND2_X1 U620 ( .A1(G56), .A2(n657), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n640), .A2(G81), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G68), .A2(n643), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n561), .Z(n562) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n650), .A2(G43), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n994) );
  INV_X1 U630 ( .A(G860), .ZN(n616) );
  OR2_X1 U631 ( .A1(n994), .A2(n616), .ZN(G153) );
  XNOR2_X1 U632 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G868), .A2(G301), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n650), .A2(G54), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G92), .A2(n640), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G79), .A2(n643), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n657), .A2(G66), .ZN(n568) );
  NOR2_X1 U639 ( .A1(n569), .A2(n511), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X2 U641 ( .A(KEYINPUT15), .B(n572), .Z(n995) );
  INV_X1 U642 ( .A(G868), .ZN(n597) );
  NAND2_X1 U643 ( .A1(n995), .A2(n597), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(G284) );
  NAND2_X1 U645 ( .A1(n640), .A2(G89), .ZN(n575) );
  XNOR2_X1 U646 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G76), .A2(n643), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U649 ( .A(n578), .B(KEYINPUT5), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n650), .A2(G51), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G63), .A2(n657), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U653 ( .A(KEYINPUT6), .B(n581), .Z(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n584), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U656 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U657 ( .A1(n650), .A2(G53), .ZN(n586) );
  NAND2_X1 U658 ( .A1(G65), .A2(n657), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G91), .A2(n640), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G78), .A2(n643), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n887) );
  INV_X1 U664 ( .A(n887), .ZN(G299) );
  NOR2_X1 U665 ( .A1(G286), .A2(n597), .ZN(n591) );
  XOR2_X1 U666 ( .A(KEYINPUT75), .B(n591), .Z(n593) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U669 ( .A(KEYINPUT76), .B(n594), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n616), .A2(G559), .ZN(n595) );
  INV_X1 U671 ( .A(n995), .ZN(n614) );
  NAND2_X1 U672 ( .A1(n595), .A2(n614), .ZN(n596) );
  XNOR2_X1 U673 ( .A(n596), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(n995), .A2(n597), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT77), .ZN(n599) );
  NOR2_X1 U676 ( .A1(G559), .A2(n599), .ZN(n601) );
  NOR2_X1 U677 ( .A1(G868), .A2(n994), .ZN(n600) );
  NOR2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U679 ( .A(KEYINPUT78), .B(n602), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G99), .A2(n976), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT80), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G111), .A2(n972), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT79), .B(n604), .Z(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G123), .A2(n973), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U687 ( .A1(G135), .A2(n977), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n984) );
  XOR2_X1 U690 ( .A(G2096), .B(n984), .Z(n612) );
  NOR2_X1 U691 ( .A1(G2100), .A2(n612), .ZN(n613) );
  XNOR2_X1 U692 ( .A(KEYINPUT81), .B(n613), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G559), .A2(n614), .ZN(n615) );
  XOR2_X1 U694 ( .A(n994), .B(n615), .Z(n666) );
  NAND2_X1 U695 ( .A1(n616), .A2(n666), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n650), .A2(G55), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G67), .A2(n657), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U699 ( .A(KEYINPUT82), .B(n619), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G93), .A2(n640), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G80), .A2(n643), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n668) );
  XOR2_X1 U704 ( .A(n624), .B(n668), .Z(G145) );
  NAND2_X1 U705 ( .A1(n650), .A2(G50), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G62), .A2(n657), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U708 ( .A(KEYINPUT86), .B(n627), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G88), .A2(n640), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G75), .A2(n643), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U712 ( .A1(n631), .A2(n630), .ZN(G166) );
  NAND2_X1 U713 ( .A1(n640), .A2(G85), .ZN(n632) );
  XOR2_X1 U714 ( .A(KEYINPUT66), .B(n632), .Z(n637) );
  NAND2_X1 U715 ( .A1(n650), .A2(G47), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G60), .A2(n657), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U718 ( .A(KEYINPUT69), .B(n635), .Z(n636) );
  NOR2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n643), .A2(G72), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U722 ( .A1(G48), .A2(n650), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G86), .A2(n640), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G73), .A2(n643), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n644), .B(KEYINPUT85), .ZN(n645) );
  XNOR2_X1 U727 ( .A(n645), .B(KEYINPUT2), .ZN(n646) );
  NOR2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G61), .A2(n657), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G49), .A2(n650), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(KEYINPUT83), .B(n653), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n654), .A2(G87), .ZN(n655) );
  XOR2_X1 U736 ( .A(KEYINPUT84), .B(n655), .Z(n656) );
  NOR2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(G288) );
  XNOR2_X1 U739 ( .A(G166), .B(n668), .ZN(n663) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n661) );
  XNOR2_X1 U741 ( .A(G290), .B(n887), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n664), .B(G305), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(G288), .ZN(n997) );
  XNOR2_X1 U746 ( .A(n666), .B(n997), .ZN(n667) );
  NAND2_X1 U747 ( .A1(n667), .A2(G868), .ZN(n670) );
  OR2_X1 U748 ( .A1(G868), .A2(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U756 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n675) );
  XNOR2_X1 U758 ( .A(n675), .B(KEYINPUT22), .ZN(n676) );
  XNOR2_X1 U759 ( .A(n676), .B(KEYINPUT88), .ZN(n677) );
  NOR2_X1 U760 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G96), .A2(n678), .ZN(n943) );
  NAND2_X1 U762 ( .A1(n943), .A2(G2106), .ZN(n684) );
  NOR2_X1 U763 ( .A1(G235), .A2(G237), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G120), .A2(n679), .ZN(n680) );
  XNOR2_X1 U765 ( .A(KEYINPUT89), .B(n680), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n681), .A2(G108), .ZN(n682) );
  XNOR2_X1 U767 ( .A(KEYINPUT90), .B(n682), .ZN(n944) );
  NAND2_X1 U768 ( .A1(n944), .A2(G567), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n1008) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n685) );
  XOR2_X1 U771 ( .A(KEYINPUT91), .B(n685), .Z(n686) );
  NOR2_X1 U772 ( .A1(n1008), .A2(n686), .ZN(n821) );
  NAND2_X1 U773 ( .A1(n821), .A2(G36), .ZN(n687) );
  XNOR2_X1 U774 ( .A(KEYINPUT92), .B(n687), .ZN(G176) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n767) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n766) );
  INV_X1 U778 ( .A(n766), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n767), .A2(n688), .ZN(n706) );
  NOR2_X1 U780 ( .A1(G2084), .A2(n706), .ZN(n736) );
  NOR2_X1 U781 ( .A1(n739), .A2(n736), .ZN(n689) );
  NAND2_X1 U782 ( .A1(G8), .A2(n689), .ZN(n690) );
  XNOR2_X1 U783 ( .A(KEYINPUT30), .B(n690), .ZN(n691) );
  XOR2_X1 U784 ( .A(KEYINPUT101), .B(n691), .Z(n692) );
  NOR2_X1 U785 ( .A1(G168), .A2(n692), .ZN(n696) );
  INV_X1 U786 ( .A(n706), .ZN(n710) );
  OR2_X1 U787 ( .A1(n710), .A2(G1961), .ZN(n694) );
  XNOR2_X1 U788 ( .A(G2078), .B(KEYINPUT25), .ZN(n861) );
  NAND2_X1 U789 ( .A1(n710), .A2(n861), .ZN(n693) );
  NAND2_X1 U790 ( .A1(n694), .A2(n693), .ZN(n724) );
  NOR2_X1 U791 ( .A1(G171), .A2(n724), .ZN(n695) );
  NOR2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U793 ( .A(n698), .B(n697), .ZN(n727) );
  NAND2_X1 U794 ( .A1(n710), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U795 ( .A(KEYINPUT27), .B(n699), .ZN(n702) );
  NAND2_X1 U796 ( .A1(G1956), .A2(n706), .ZN(n700) );
  XOR2_X1 U797 ( .A(KEYINPUT98), .B(n700), .Z(n701) );
  NOR2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n718) );
  NOR2_X1 U799 ( .A1(n887), .A2(n718), .ZN(n704) );
  XNOR2_X1 U800 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n703) );
  XNOR2_X1 U801 ( .A(n704), .B(n703), .ZN(n722) );
  XNOR2_X1 U802 ( .A(G1996), .B(KEYINPUT100), .ZN(n862) );
  NAND2_X1 U803 ( .A1(n862), .A2(n710), .ZN(n705) );
  XNOR2_X1 U804 ( .A(n705), .B(KEYINPUT26), .ZN(n708) );
  BUF_X1 U805 ( .A(n706), .Z(n728) );
  NAND2_X1 U806 ( .A1(n728), .A2(G1341), .ZN(n707) );
  NAND2_X1 U807 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U808 ( .A1(n994), .A2(n709), .ZN(n714) );
  NAND2_X1 U809 ( .A1(G1348), .A2(n728), .ZN(n712) );
  NAND2_X1 U810 ( .A1(G2067), .A2(n710), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n995), .A2(n715), .ZN(n713) );
  OR2_X1 U813 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n995), .A2(n715), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U816 ( .A1(n887), .A2(n718), .ZN(n719) );
  NAND2_X1 U817 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U818 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U819 ( .A(n723), .B(KEYINPUT29), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n737) );
  NAND2_X1 U821 ( .A1(n737), .A2(G286), .ZN(n733) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n764), .ZN(n730) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n731), .A2(G303), .ZN(n732) );
  NAND2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n734), .A2(G8), .ZN(n735) );
  XNOR2_X1 U828 ( .A(n735), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U829 ( .A1(G8), .A2(n736), .ZN(n741) );
  INV_X1 U830 ( .A(n737), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n756) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n744) );
  OR2_X1 U836 ( .A1(n750), .A2(n744), .ZN(n905) );
  XOR2_X1 U837 ( .A(KEYINPUT102), .B(n905), .Z(n745) );
  NAND2_X1 U838 ( .A1(n756), .A2(n745), .ZN(n748) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n892) );
  NOR2_X1 U840 ( .A1(n764), .A2(n746), .ZN(n747) );
  NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n749), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n764), .A2(n751), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n897) );
  NAND2_X1 U846 ( .A1(n754), .A2(n897), .ZN(n760) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U848 ( .A1(G8), .A2(n755), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n758), .A2(n764), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U853 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n812) );
  NAND2_X1 U855 ( .A1(G104), .A2(n976), .ZN(n769) );
  NAND2_X1 U856 ( .A1(G140), .A2(n977), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U858 ( .A(KEYINPUT34), .B(n770), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n972), .A2(G116), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G128), .A2(n973), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT35), .B(n773), .Z(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U864 ( .A(KEYINPUT36), .B(n776), .ZN(n990) );
  XNOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NOR2_X1 U866 ( .A1(n990), .A2(n810), .ZN(n834) );
  NAND2_X1 U867 ( .A1(n812), .A2(n834), .ZN(n808) );
  NAND2_X1 U868 ( .A1(n972), .A2(G107), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G119), .A2(n973), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G95), .A2(n976), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G131), .A2(n977), .ZN(n779) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT94), .B(n783), .Z(n965) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n965), .ZN(n784) );
  XNOR2_X1 U877 ( .A(n784), .B(KEYINPUT95), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G105), .A2(n976), .ZN(n785) );
  XNOR2_X1 U879 ( .A(n785), .B(KEYINPUT38), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n977), .A2(G141), .ZN(n787) );
  NAND2_X1 U881 ( .A1(G129), .A2(n973), .ZN(n786) );
  NAND2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U883 ( .A1(n972), .A2(G117), .ZN(n788) );
  XOR2_X1 U884 ( .A(KEYINPUT96), .B(n788), .Z(n789) );
  NOR2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n986) );
  AND2_X1 U887 ( .A1(G1996), .A2(n986), .ZN(n793) );
  NOR2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n853) );
  INV_X1 U889 ( .A(n812), .ZN(n795) );
  NOR2_X1 U890 ( .A1(n853), .A2(n795), .ZN(n804) );
  INV_X1 U891 ( .A(n804), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n808), .A2(n796), .ZN(n797) );
  XOR2_X1 U893 ( .A(KEYINPUT97), .B(n797), .Z(n798) );
  NOR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n801) );
  XNOR2_X1 U895 ( .A(G1986), .B(G290), .ZN(n904) );
  NAND2_X1 U896 ( .A1(n904), .A2(n812), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n815) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n986), .ZN(n831) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n965), .ZN(n840) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n840), .A2(n802), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U903 ( .A(n805), .B(KEYINPUT104), .ZN(n806) );
  NOR2_X1 U904 ( .A1(n831), .A2(n806), .ZN(n807) );
  XNOR2_X1 U905 ( .A(KEYINPUT39), .B(n807), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n990), .A2(n810), .ZN(n837) );
  NAND2_X1 U908 ( .A1(n811), .A2(n837), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n817) );
  XOR2_X1 U911 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n816) );
  XNOR2_X1 U912 ( .A(n817), .B(n816), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U915 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(G188) );
  XOR2_X1 U918 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  NAND2_X1 U920 ( .A1(G112), .A2(n972), .ZN(n823) );
  NAND2_X1 U921 ( .A1(G100), .A2(n976), .ZN(n822) );
  NAND2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n973), .A2(G124), .ZN(n824) );
  XNOR2_X1 U924 ( .A(n824), .B(KEYINPUT110), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n825), .B(KEYINPUT44), .ZN(n827) );
  NAND2_X1 U926 ( .A1(G136), .A2(n977), .ZN(n826) );
  NAND2_X1 U927 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U928 ( .A1(n829), .A2(n828), .ZN(G162) );
  XOR2_X1 U929 ( .A(G2090), .B(G162), .Z(n830) );
  NOR2_X1 U930 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n832), .B(KEYINPUT51), .ZN(n833) );
  NOR2_X1 U932 ( .A1(n834), .A2(n833), .ZN(n842) );
  XNOR2_X1 U933 ( .A(G2084), .B(G160), .ZN(n835) );
  XNOR2_X1 U934 ( .A(KEYINPUT115), .B(n835), .ZN(n836) );
  NOR2_X1 U935 ( .A1(n984), .A2(n836), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U937 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n856) );
  NAND2_X1 U939 ( .A1(G103), .A2(n976), .ZN(n844) );
  NAND2_X1 U940 ( .A1(G139), .A2(n977), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n849) );
  NAND2_X1 U942 ( .A1(n972), .A2(G115), .ZN(n846) );
  NAND2_X1 U943 ( .A1(G127), .A2(n973), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(KEYINPUT47), .B(n847), .Z(n848) );
  NOR2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n968) );
  XOR2_X1 U947 ( .A(G2072), .B(n968), .Z(n851) );
  XOR2_X1 U948 ( .A(G164), .B(G2078), .Z(n850) );
  NOR2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U950 ( .A(KEYINPUT50), .B(n852), .ZN(n854) );
  NAND2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U952 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U953 ( .A(KEYINPUT52), .B(n857), .ZN(n858) );
  INV_X1 U954 ( .A(KEYINPUT55), .ZN(n883) );
  NAND2_X1 U955 ( .A1(n858), .A2(n883), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n859), .A2(G29), .ZN(n941) );
  XNOR2_X1 U957 ( .A(G1991), .B(G25), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n860), .B(KEYINPUT116), .ZN(n872) );
  XNOR2_X1 U959 ( .A(G27), .B(n861), .ZN(n866) );
  XNOR2_X1 U960 ( .A(n862), .B(G32), .ZN(n864) );
  XNOR2_X1 U961 ( .A(G26), .B(G2067), .ZN(n863) );
  NOR2_X1 U962 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n869) );
  XOR2_X1 U964 ( .A(KEYINPUT117), .B(G2072), .Z(n867) );
  XNOR2_X1 U965 ( .A(G33), .B(n867), .ZN(n868) );
  NOR2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U967 ( .A(KEYINPUT118), .B(n870), .Z(n871) );
  NOR2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G28), .A2(n873), .ZN(n876) );
  XOR2_X1 U970 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n874) );
  XNOR2_X1 U971 ( .A(KEYINPUT53), .B(n874), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n876), .B(n875), .ZN(n881) );
  XNOR2_X1 U973 ( .A(G2084), .B(G34), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n877), .B(KEYINPUT54), .ZN(n879) );
  XNOR2_X1 U975 ( .A(G35), .B(G2090), .ZN(n878) );
  NOR2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n883), .B(n882), .ZN(n885) );
  INV_X1 U979 ( .A(G29), .ZN(n884) );
  NAND2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G11), .A2(n886), .ZN(n939) );
  XNOR2_X1 U982 ( .A(G16), .B(KEYINPUT56), .ZN(n909) );
  XNOR2_X1 U983 ( .A(G1956), .B(n887), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G1971), .A2(G303), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U986 ( .A(G1341), .B(n994), .ZN(n890) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n903) );
  XOR2_X1 U989 ( .A(G171), .B(G1961), .Z(n895) );
  XNOR2_X1 U990 ( .A(n995), .B(G1348), .ZN(n894) );
  NOR2_X1 U991 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U992 ( .A(KEYINPUT121), .B(n896), .Z(n901) );
  XNOR2_X1 U993 ( .A(G1966), .B(G168), .ZN(n898) );
  NAND2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n899), .B(KEYINPUT57), .ZN(n900) );
  NAND2_X1 U996 ( .A1(n901), .A2(n900), .ZN(n902) );
  NOR2_X1 U997 ( .A1(n903), .A2(n902), .ZN(n907) );
  NOR2_X1 U998 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U999 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1000 ( .A1(n909), .A2(n908), .ZN(n937) );
  XOR2_X1 U1001 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n933) );
  XNOR2_X1 U1002 ( .A(G1961), .B(G5), .ZN(n923) );
  XOR2_X1 U1003 ( .A(G1956), .B(G20), .Z(n914) );
  XNOR2_X1 U1004 ( .A(G1981), .B(G6), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(G1341), .B(G19), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(KEYINPUT122), .B(n912), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n917) );
  XOR2_X1 U1009 ( .A(KEYINPUT59), .B(G1348), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G4), .B(n915), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1012 ( .A(KEYINPUT60), .B(n918), .Z(n920) );
  XNOR2_X1 U1013 ( .A(G1966), .B(G21), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(KEYINPUT123), .B(n921), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n931) );
  XOR2_X1 U1017 ( .A(G1976), .B(KEYINPUT124), .Z(n924) );
  XNOR2_X1 U1018 ( .A(G23), .B(n924), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(G1986), .B(G24), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(G1971), .B(G22), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1023 ( .A(KEYINPUT58), .B(n929), .Z(n930) );
  NAND2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1025 ( .A(n933), .B(n932), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(G16), .A2(n934), .ZN(n935) );
  XOR2_X1 U1027 ( .A(KEYINPUT126), .B(n935), .Z(n936) );
  NAND2_X1 U1028 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1030 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1031 ( .A(KEYINPUT62), .B(n942), .Z(G311) );
  XNOR2_X1 U1032 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1033 ( .A(G132), .ZN(G219) );
  INV_X1 U1034 ( .A(G108), .ZN(G238) );
  INV_X1 U1035 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(G325) );
  INV_X1 U1037 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1038 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n946) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G2072), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n946), .B(n945), .ZN(n950) );
  XOR2_X1 U1041 ( .A(G2678), .B(KEYINPUT107), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G2067), .B(KEYINPUT42), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n948), .B(n947), .ZN(n949) );
  XOR2_X1 U1044 ( .A(n950), .B(n949), .Z(n952) );
  XNOR2_X1 U1045 ( .A(G2096), .B(G2100), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n952), .B(n951), .ZN(n954) );
  XOR2_X1 U1047 ( .A(G2078), .B(G2084), .Z(n953) );
  XNOR2_X1 U1048 ( .A(n954), .B(n953), .ZN(G227) );
  XOR2_X1 U1049 ( .A(G1971), .B(G1956), .Z(n956) );
  XNOR2_X1 U1050 ( .A(G1996), .B(G1981), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n956), .B(n955), .ZN(n960) );
  XOR2_X1 U1052 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n958) );
  XNOR2_X1 U1053 ( .A(G1991), .B(G1961), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n958), .B(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(n960), .B(n959), .Z(n962) );
  XNOR2_X1 U1056 ( .A(G1976), .B(G2474), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n962), .B(n961), .ZN(n964) );
  XOR2_X1 U1058 ( .A(G1986), .B(G1966), .Z(n963) );
  XNOR2_X1 U1059 ( .A(n964), .B(n963), .ZN(G229) );
  XOR2_X1 U1060 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n967) );
  XNOR2_X1 U1061 ( .A(n965), .B(KEYINPUT48), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(n967), .B(n966), .ZN(n969) );
  XOR2_X1 U1063 ( .A(n969), .B(n968), .Z(n971) );
  XNOR2_X1 U1064 ( .A(G160), .B(G164), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n971), .B(n970), .ZN(n992) );
  NAND2_X1 U1066 ( .A1(n972), .A2(G118), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(G130), .A2(n973), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n983) );
  NAND2_X1 U1069 ( .A1(G106), .A2(n976), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(G142), .A2(n977), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(KEYINPUT111), .B(n980), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT45), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n985) );
  XOR2_X1 U1075 ( .A(n985), .B(n984), .Z(n988) );
  XOR2_X1 U1076 ( .A(n986), .B(G162), .Z(n987) );
  XNOR2_X1 U1077 ( .A(n988), .B(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(n992), .B(n991), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(G37), .A2(n993), .ZN(G395) );
  XNOR2_X1 U1081 ( .A(G286), .B(n994), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(n996), .B(n995), .ZN(n999) );
  XOR2_X1 U1083 ( .A(G171), .B(n997), .Z(n998) );
  XNOR2_X1 U1084 ( .A(n999), .B(n998), .ZN(n1000) );
  NOR2_X1 U1085 ( .A1(G37), .A2(n1000), .ZN(G397) );
  NOR2_X1 U1086 ( .A1(G401), .A2(n1008), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(KEYINPUT113), .B(n1001), .ZN(n1004) );
  NOR2_X1 U1088 ( .A1(G227), .A2(G229), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT49), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(KEYINPUT114), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1092 ( .A1(G395), .A2(G397), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(G225) );
  INV_X1 U1094 ( .A(G225), .ZN(G308) );
  INV_X1 U1095 ( .A(n1008), .ZN(G319) );
  INV_X1 U1096 ( .A(G96), .ZN(G221) );
endmodule

