

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585;

  NOR2_X1 U326 ( .A1(n464), .A2(n514), .ZN(n460) );
  XNOR2_X1 U327 ( .A(n318), .B(n317), .ZN(n319) );
  INV_X1 U328 ( .A(n527), .ZN(n528) );
  XNOR2_X1 U329 ( .A(n390), .B(n295), .ZN(n326) );
  XOR2_X1 U330 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n294) );
  XOR2_X1 U331 ( .A(n325), .B(n324), .Z(n295) );
  INV_X1 U332 ( .A(KEYINPUT96), .ZN(n379) );
  XNOR2_X1 U333 ( .A(n448), .B(n316), .ZN(n317) );
  XNOR2_X1 U334 ( .A(n373), .B(KEYINPUT48), .ZN(n527) );
  XNOR2_X1 U335 ( .A(n380), .B(n379), .ZN(n381) );
  NOR2_X1 U336 ( .A1(n579), .A2(n487), .ZN(n488) );
  XNOR2_X1 U337 ( .A(n430), .B(n381), .ZN(n382) );
  XNOR2_X1 U338 ( .A(n436), .B(KEYINPUT55), .ZN(n437) );
  XNOR2_X1 U339 ( .A(n452), .B(n387), .ZN(n388) );
  XNOR2_X1 U340 ( .A(n438), .B(n437), .ZN(n455) );
  XNOR2_X1 U341 ( .A(n327), .B(n326), .ZN(n364) );
  XNOR2_X1 U342 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U343 ( .A(n454), .B(n453), .Z(n520) );
  XNOR2_X1 U344 ( .A(n491), .B(KEYINPUT38), .ZN(n498) );
  XNOR2_X1 U345 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U346 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n297) );
  XNOR2_X1 U348 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U350 ( .A(G106GAT), .B(n298), .ZN(n302) );
  XOR2_X1 U351 ( .A(G162GAT), .B(G218GAT), .Z(n425) );
  XOR2_X1 U352 ( .A(G190GAT), .B(KEYINPUT77), .Z(n374) );
  XOR2_X1 U353 ( .A(n425), .B(n374), .Z(n300) );
  NAND2_X1 U354 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(n303), .B(KEYINPUT11), .Z(n305) );
  XOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .Z(n315) );
  XNOR2_X1 U359 ( .A(G92GAT), .B(n315), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U361 ( .A(G29GAT), .B(KEYINPUT7), .Z(n307) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G36GAT), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U364 ( .A(G50GAT), .B(KEYINPUT8), .Z(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n332) );
  XNOR2_X1 U366 ( .A(n310), .B(n332), .ZN(n556) );
  XOR2_X1 U367 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n312) );
  XNOR2_X1 U368 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U370 ( .A(G57GAT), .B(KEYINPUT13), .Z(n347) );
  XOR2_X1 U371 ( .A(n313), .B(n347), .Z(n320) );
  XNOR2_X1 U372 ( .A(G148GAT), .B(G106GAT), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n314), .B(G78GAT), .ZN(n431) );
  XOR2_X1 U374 ( .A(n315), .B(n431), .Z(n318) );
  XOR2_X1 U375 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  NAND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n327) );
  XOR2_X1 U378 ( .A(G92GAT), .B(G64GAT), .Z(n322) );
  XNOR2_X1 U379 ( .A(G176GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U381 ( .A(KEYINPUT73), .B(n323), .ZN(n390) );
  XOR2_X1 U382 ( .A(KEYINPUT71), .B(KEYINPUT75), .Z(n325) );
  XNOR2_X1 U383 ( .A(KEYINPUT74), .B(KEYINPUT72), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n364), .B(KEYINPUT41), .ZN(n560) );
  XOR2_X1 U385 ( .A(G169GAT), .B(G8GAT), .Z(n375) );
  XOR2_X1 U386 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n329) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U389 ( .A(n375), .B(n330), .Z(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U391 ( .A(G113GAT), .B(G197GAT), .Z(n334) );
  XNOR2_X1 U392 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U394 ( .A(n336), .B(n335), .Z(n338) );
  XOR2_X1 U395 ( .A(G15GAT), .B(G1GAT), .Z(n348) );
  XOR2_X1 U396 ( .A(G141GAT), .B(G22GAT), .Z(n421) );
  XNOR2_X1 U397 ( .A(n348), .B(n421), .ZN(n337) );
  XOR2_X1 U398 ( .A(n338), .B(n337), .Z(n571) );
  INV_X1 U399 ( .A(n571), .ZN(n547) );
  NOR2_X1 U400 ( .A1(n560), .A2(n547), .ZN(n340) );
  XOR2_X1 U401 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n360) );
  XOR2_X1 U403 ( .A(G78GAT), .B(G71GAT), .Z(n342) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(G8GAT), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U406 ( .A(KEYINPUT15), .B(G211GAT), .Z(n344) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(G127GAT), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U409 ( .A(n346), .B(n345), .Z(n350) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U412 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n352) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U415 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n356) );
  XNOR2_X1 U417 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U419 ( .A(G155GAT), .B(n357), .ZN(n358) );
  XOR2_X1 U420 ( .A(n359), .B(n358), .Z(n566) );
  INV_X1 U421 ( .A(n566), .ZN(n579) );
  NOR2_X1 U422 ( .A1(n360), .A2(n579), .ZN(n361) );
  AND2_X1 U423 ( .A1(n556), .A2(n361), .ZN(n363) );
  INV_X1 U424 ( .A(KEYINPUT47), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n371) );
  XOR2_X1 U426 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n367) );
  XNOR2_X1 U427 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n556), .B(n365), .ZN(n582) );
  NAND2_X1 U429 ( .A1(n579), .A2(n582), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n571), .B(KEYINPUT69), .ZN(n558) );
  NAND2_X1 U432 ( .A1(n368), .A2(n558), .ZN(n369) );
  NOR2_X1 U433 ( .A1(n364), .A2(n369), .ZN(n370) );
  NOR2_X1 U434 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n372), .B(KEYINPUT64), .ZN(n373) );
  XOR2_X1 U436 ( .A(KEYINPUT95), .B(KEYINPUT78), .Z(n377) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n383) );
  XNOR2_X1 U439 ( .A(G197GAT), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n294), .B(n378), .ZN(n430) );
  NAND2_X1 U441 ( .A1(G226GAT), .A2(G233GAT), .ZN(n380) );
  XOR2_X1 U442 ( .A(n383), .B(n382), .Z(n389) );
  XOR2_X1 U443 ( .A(KEYINPUT17), .B(G183GAT), .Z(n385) );
  XNOR2_X1 U444 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(KEYINPUT85), .B(n386), .Z(n452) );
  XNOR2_X1 U447 ( .A(G36GAT), .B(G218GAT), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n517) );
  NOR2_X1 U449 ( .A1(n527), .A2(n517), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n392), .B(KEYINPUT54), .ZN(n414) );
  XOR2_X1 U451 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n394) );
  XNOR2_X1 U452 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n424) );
  XOR2_X1 U454 ( .A(G162GAT), .B(n424), .Z(n396) );
  NAND2_X1 U455 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(n397), .ZN(n413) );
  XOR2_X1 U458 ( .A(G148GAT), .B(G85GAT), .Z(n399) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(G141GAT), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U461 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n401) );
  XNOR2_X1 U462 ( .A(G120GAT), .B(G57GAT), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U464 ( .A(n403), .B(n402), .Z(n411) );
  XOR2_X1 U465 ( .A(G134GAT), .B(KEYINPUT0), .Z(n405) );
  XNOR2_X1 U466 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U468 ( .A(G127GAT), .B(n406), .ZN(n453) );
  XOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n408) );
  XNOR2_X1 U470 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U472 ( .A(n453), .B(n409), .Z(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n514) );
  NAND2_X1 U475 ( .A1(n414), .A2(n514), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n415), .B(KEYINPUT65), .ZN(n568) );
  XOR2_X1 U477 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n417) );
  XNOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT91), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n435) );
  XOR2_X1 U480 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n419) );
  XNOR2_X1 U481 ( .A(KEYINPUT86), .B(KEYINPUT90), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U483 ( .A(n420), .B(G204GAT), .Z(n423) );
  XNOR2_X1 U484 ( .A(G50GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n429) );
  XOR2_X1 U486 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U489 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U492 ( .A(n435), .B(n434), .Z(n466) );
  NAND2_X1 U493 ( .A1(n568), .A2(n466), .ZN(n438) );
  XOR2_X1 U494 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n436) );
  XOR2_X1 U495 ( .A(G99GAT), .B(G190GAT), .Z(n440) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(G43GAT), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U498 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n442) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(G176GAT), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U501 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n446) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n454) );
  INV_X1 U508 ( .A(n520), .ZN(n531) );
  NAND2_X1 U509 ( .A1(n455), .A2(n531), .ZN(n565) );
  NOR2_X1 U510 ( .A1(n556), .A2(n565), .ZN(n459) );
  XNOR2_X1 U511 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n457) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n456) );
  NOR2_X1 U513 ( .A1(n558), .A2(n364), .ZN(n490) );
  XNOR2_X1 U514 ( .A(n517), .B(KEYINPUT27), .ZN(n464) );
  XOR2_X1 U515 ( .A(KEYINPUT97), .B(n460), .Z(n529) );
  XNOR2_X1 U516 ( .A(n466), .B(KEYINPUT28), .ZN(n523) );
  INV_X1 U517 ( .A(n523), .ZN(n530) );
  NOR2_X1 U518 ( .A1(n530), .A2(n531), .ZN(n461) );
  NAND2_X1 U519 ( .A1(n529), .A2(n461), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT98), .ZN(n474) );
  NOR2_X1 U521 ( .A1(n531), .A2(n466), .ZN(n463) );
  XOR2_X1 U522 ( .A(n463), .B(KEYINPUT26), .Z(n569) );
  OR2_X1 U523 ( .A1(n464), .A2(n569), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n520), .A2(n517), .ZN(n465) );
  XNOR2_X1 U525 ( .A(KEYINPUT99), .B(n465), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(KEYINPUT100), .Z(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n472), .A2(n514), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n486) );
  NAND2_X1 U532 ( .A1(n556), .A2(n579), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  AND2_X1 U534 ( .A1(n486), .A2(n476), .ZN(n502) );
  NAND2_X1 U535 ( .A1(n490), .A2(n502), .ZN(n484) );
  NOR2_X1 U536 ( .A1(n514), .A2(n484), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n517), .A2(n484), .ZN(n480) );
  XOR2_X1 U541 ( .A(G8GAT), .B(n480), .Z(G1325GAT) );
  NOR2_X1 U542 ( .A1(n520), .A2(n484), .ZN(n482) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n523), .A2(n484), .ZN(n485) );
  XOR2_X1 U547 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  NAND2_X1 U548 ( .A1(n582), .A2(n486), .ZN(n487) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n488), .Z(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(n489), .ZN(n512) );
  NAND2_X1 U551 ( .A1(n512), .A2(n490), .ZN(n491) );
  NOR2_X1 U552 ( .A1(n514), .A2(n498), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n498), .A2(n517), .ZN(n494) );
  XOR2_X1 U556 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U557 ( .A1(n520), .A2(n498), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n498), .A2(n523), .ZN(n500) );
  XNOR2_X1 U562 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  NOR2_X1 U565 ( .A1(n571), .A2(n560), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n513), .A2(n502), .ZN(n509) );
  NOR2_X1 U567 ( .A1(n514), .A2(n509), .ZN(n503) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n503), .Z(n504) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n517), .A2(n509), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(n505), .Z(n506) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n520), .A2(n509), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n522) );
  NOR2_X1 U580 ( .A1(n514), .A2(n522), .ZN(n515) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n515), .Z(n516) );
  XNOR2_X1 U582 ( .A(KEYINPUT110), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n522), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n522), .ZN(n521) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U591 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n545) );
  NOR2_X1 U593 ( .A1(n530), .A2(n545), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(n533), .ZN(n542) );
  NOR2_X1 U596 ( .A1(n558), .A2(n542), .ZN(n534) );
  XOR2_X1 U597 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  NOR2_X1 U598 ( .A1(n542), .A2(n560), .ZN(n536) );
  XNOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n539) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n542), .A2(n566), .ZN(n540) );
  XOR2_X1 U606 ( .A(n541), .B(n540), .Z(G1342GAT) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n544) );
  NOR2_X1 U608 ( .A1(n556), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n549) );
  NOR2_X1 U611 ( .A1(n569), .A2(n545), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(n546), .Z(n555) );
  NOR2_X1 U613 ( .A1(n547), .A2(n555), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n551) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n555), .A2(n560), .ZN(n552) );
  XOR2_X1 U619 ( .A(n553), .B(n552), .Z(G1345GAT) );
  NOR2_X1 U620 ( .A1(n555), .A2(n566), .ZN(n554) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n554), .Z(G1346GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  NOR2_X1 U624 ( .A1(n565), .A2(n558), .ZN(n559) );
  XOR2_X1 U625 ( .A(G169GAT), .B(n559), .Z(G1348GAT) );
  NOR2_X1 U626 ( .A1(n565), .A2(n560), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  INV_X1 U633 ( .A(n568), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n583) );
  AND2_X1 U635 ( .A1(n583), .A2(n571), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n577) );
  NAND2_X1 U641 ( .A1(n583), .A2(n364), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n583), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

