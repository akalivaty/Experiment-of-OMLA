

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792;

  XNOR2_X1 U380 ( .A(n627), .B(n628), .ZN(n699) );
  XNOR2_X1 U381 ( .A(n358), .B(n773), .ZN(n494) );
  XNOR2_X1 U382 ( .A(n492), .B(n491), .ZN(n358) );
  NOR2_X1 U383 ( .A1(n699), .A2(n629), .ZN(n631) );
  XNOR2_X2 U384 ( .A(n432), .B(KEYINPUT19), .ZN(n598) );
  NAND2_X1 U385 ( .A1(n671), .A2(n383), .ZN(n582) );
  XNOR2_X2 U386 ( .A(n574), .B(n573), .ZN(n671) );
  NOR2_X2 U387 ( .A1(n705), .A2(n687), .ZN(n561) );
  XNOR2_X2 U388 ( .A(n440), .B(KEYINPUT90), .ZN(n775) );
  XOR2_X1 U389 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n490) );
  INV_X2 U390 ( .A(G953), .ZN(n778) );
  AND2_X2 U391 ( .A1(n455), .A2(n368), .ZN(n457) );
  AND2_X2 U392 ( .A1(n404), .A2(KEYINPUT1), .ZN(n386) );
  OR2_X2 U393 ( .A1(n681), .A2(n452), .ZN(n411) );
  XNOR2_X1 U394 ( .A(n360), .B(n361), .ZN(n577) );
  NOR2_X1 U395 ( .A1(n568), .A2(n363), .ZN(n360) );
  NAND2_X1 U396 ( .A1(n604), .A2(n433), .ZN(n432) );
  AND2_X1 U397 ( .A1(n396), .A2(n395), .ZN(n394) );
  NOR2_X1 U398 ( .A1(n577), .A2(n389), .ZN(n382) );
  NOR2_X1 U399 ( .A1(n752), .A2(n621), .ZN(n622) );
  NAND2_X1 U400 ( .A1(n576), .A2(n390), .ZN(n389) );
  NOR2_X1 U401 ( .A1(n577), .A2(n530), .ZN(n531) );
  XOR2_X1 U402 ( .A(KEYINPUT41), .B(n618), .Z(n752) );
  XOR2_X1 U403 ( .A(n642), .B(KEYINPUT38), .Z(n721) );
  XNOR2_X1 U404 ( .A(n501), .B(n500), .ZN(n571) );
  INV_X1 U405 ( .A(KEYINPUT32), .ZN(n381) );
  XOR2_X1 U406 ( .A(G101), .B(KEYINPUT65), .Z(n520) );
  BUF_X1 U407 ( .A(n639), .Z(n359) );
  XOR2_X1 U408 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n361) );
  AND2_X1 U409 ( .A1(n788), .A2(n578), .ZN(n383) );
  XNOR2_X1 U410 ( .A(n766), .B(n465), .ZN(n518) );
  XNOR2_X1 U411 ( .A(n520), .B(KEYINPUT68), .ZN(n465) );
  AND2_X1 U412 ( .A1(n411), .A2(n409), .ZN(n406) );
  OR2_X1 U413 ( .A1(n660), .A2(G472), .ZN(n421) );
  XNOR2_X1 U414 ( .A(G104), .B(G122), .ZN(n489) );
  AND2_X1 U415 ( .A1(n650), .A2(n711), .ZN(n449) );
  NAND2_X1 U416 ( .A1(n649), .A2(n446), .ZN(n445) );
  NAND2_X1 U417 ( .A1(KEYINPUT64), .A2(KEYINPUT2), .ZN(n446) );
  AND2_X1 U418 ( .A1(n626), .A2(n400), .ZN(n399) );
  NAND2_X1 U419 ( .A1(n732), .A2(KEYINPUT81), .ZN(n400) );
  NOR2_X1 U420 ( .A1(G237), .A2(G953), .ZN(n495) );
  XNOR2_X1 U421 ( .A(n466), .B(G146), .ZN(n488) );
  INV_X1 U422 ( .A(G125), .ZN(n466) );
  XNOR2_X1 U423 ( .A(n427), .B(n426), .ZN(n538) );
  INV_X1 U424 ( .A(KEYINPUT8), .ZN(n426) );
  NAND2_X1 U425 ( .A1(n778), .A2(G234), .ZN(n427) );
  XOR2_X1 U426 ( .A(G146), .B(G140), .Z(n516) );
  XOR2_X1 U427 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n569) );
  NAND2_X1 U428 ( .A1(n639), .A2(n552), .ZN(n554) );
  AND2_X1 U429 ( .A1(n660), .A2(n420), .ZN(n419) );
  AND2_X1 U430 ( .A1(G472), .A2(n543), .ZN(n420) );
  NAND2_X1 U431 ( .A1(n543), .A2(n453), .ZN(n452) );
  INV_X1 U432 ( .A(G469), .ZN(n453) );
  XNOR2_X1 U433 ( .A(KEYINPUT4), .B(G137), .ZN(n512) );
  XNOR2_X1 U434 ( .A(n439), .B(n438), .ZN(n525) );
  XNOR2_X1 U435 ( .A(KEYINPUT3), .B(KEYINPUT84), .ZN(n438) );
  NAND2_X1 U436 ( .A1(n462), .A2(n463), .ZN(n439) );
  XNOR2_X1 U437 ( .A(n437), .B(G122), .ZN(n504) );
  INV_X1 U438 ( .A(G116), .ZN(n437) );
  XNOR2_X1 U439 ( .A(KEYINPUT75), .B(G110), .ZN(n464) );
  XOR2_X1 U440 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n503) );
  INV_X1 U441 ( .A(KEYINPUT98), .ZN(n430) );
  AND2_X2 U442 ( .A1(n422), .A2(n647), .ZN(n777) );
  XNOR2_X1 U443 ( .A(n423), .B(n372), .ZN(n422) );
  XNOR2_X1 U444 ( .A(n413), .B(KEYINPUT39), .ZN(n645) );
  INV_X1 U445 ( .A(n721), .ZN(n414) );
  INV_X1 U446 ( .A(n735), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n507), .B(n425), .ZN(n560) );
  INV_X1 U448 ( .A(G478), .ZN(n425) );
  NAND2_X1 U449 ( .A1(n374), .A2(n365), .ZN(n578) );
  INV_X1 U450 ( .A(KEYINPUT70), .ZN(n583) );
  INV_X1 U451 ( .A(KEYINPUT1), .ZN(n409) );
  NOR2_X1 U452 ( .A1(n411), .A2(n409), .ZN(n408) );
  INV_X1 U453 ( .A(G113), .ZN(n461) );
  XNOR2_X1 U454 ( .A(KEYINPUT66), .B(G131), .ZN(n513) );
  XOR2_X1 U455 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n491) );
  NAND2_X1 U456 ( .A1(n447), .A2(n445), .ZN(n444) );
  NAND2_X1 U457 ( .A1(n508), .A2(KEYINPUT64), .ZN(n447) );
  NAND2_X1 U458 ( .A1(n398), .A2(KEYINPUT81), .ZN(n395) );
  NAND2_X1 U459 ( .A1(n631), .A2(n630), .ZN(n637) );
  AND2_X1 U460 ( .A1(n417), .A2(n421), .ZN(n605) );
  OR2_X1 U461 ( .A1(n720), .A2(n367), .ZN(n418) );
  XOR2_X1 U462 ( .A(G128), .B(G137), .Z(n459) );
  XOR2_X1 U463 ( .A(G110), .B(G119), .Z(n537) );
  XNOR2_X1 U464 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n532) );
  XNOR2_X1 U465 ( .A(n488), .B(n388), .ZN(n773) );
  XNOR2_X1 U466 ( .A(G140), .B(KEYINPUT10), .ZN(n388) );
  XNOR2_X1 U467 ( .A(n775), .B(n519), .ZN(n681) );
  NAND2_X1 U468 ( .A1(n450), .A2(n366), .ZN(n714) );
  XNOR2_X1 U469 ( .A(n637), .B(n387), .ZN(n633) );
  INV_X1 U470 ( .A(KEYINPUT110), .ZN(n387) );
  NAND2_X1 U471 ( .A1(n416), .A2(n421), .ZN(n738) );
  OR2_X1 U472 ( .A1(n588), .A2(n551), .ZN(n731) );
  XNOR2_X1 U473 ( .A(n588), .B(n548), .ZN(n735) );
  XNOR2_X1 U474 ( .A(n527), .B(n528), .ZN(n660) );
  XNOR2_X1 U475 ( .A(n525), .B(n434), .ZN(n768) );
  XNOR2_X1 U476 ( .A(n504), .B(n435), .ZN(n434) );
  XNOR2_X1 U477 ( .A(n436), .B(KEYINPUT16), .ZN(n435) );
  INV_X1 U478 ( .A(KEYINPUT73), .ZN(n436) );
  XNOR2_X1 U479 ( .A(n431), .B(n428), .ZN(n676) );
  XNOR2_X1 U480 ( .A(n505), .B(n429), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n503), .B(n430), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n412), .B(n624), .ZN(n786) );
  INV_X1 U483 ( .A(KEYINPUT35), .ZN(n573) );
  INV_X1 U484 ( .A(n578), .ZN(n692) );
  AND2_X1 U485 ( .A1(n378), .A2(n714), .ZN(n379) );
  XOR2_X1 U486 ( .A(G104), .B(G107), .Z(n362) );
  NAND2_X1 U487 ( .A1(n722), .A2(n734), .ZN(n363) );
  NAND2_X1 U488 ( .A1(G902), .A2(G469), .ZN(n364) );
  AND2_X1 U489 ( .A1(n738), .A2(n588), .ZN(n365) );
  AND2_X1 U490 ( .A1(n777), .A2(KEYINPUT2), .ZN(n366) );
  AND2_X1 U491 ( .A1(G902), .A2(n659), .ZN(n367) );
  AND2_X1 U492 ( .A1(n458), .A2(n610), .ZN(n368) );
  NOR2_X1 U493 ( .A1(n568), .A2(n569), .ZN(n369) );
  AND2_X1 U494 ( .A1(n403), .A2(n359), .ZN(n370) );
  INV_X1 U495 ( .A(KEYINPUT81), .ZN(n402) );
  XOR2_X1 U496 ( .A(n634), .B(KEYINPUT111), .Z(n371) );
  INV_X1 U497 ( .A(n508), .ZN(n649) );
  XOR2_X1 U498 ( .A(n636), .B(KEYINPUT67), .Z(n372) );
  AND2_X1 U499 ( .A1(n649), .A2(KEYINPUT64), .ZN(n373) );
  NAND2_X1 U500 ( .A1(n454), .A2(n364), .ZN(n404) );
  NAND2_X1 U501 ( .A1(n407), .A2(n405), .ZN(n639) );
  NOR2_X1 U502 ( .A1(n408), .A2(n386), .ZN(n407) );
  NOR2_X1 U503 ( .A1(n577), .A2(n359), .ZN(n374) );
  XNOR2_X1 U504 ( .A(n382), .B(n381), .ZN(n788) );
  XNOR2_X1 U505 ( .A(n385), .B(KEYINPUT45), .ZN(n760) );
  NOR2_X1 U506 ( .A1(G902), .A2(n665), .ZN(n501) );
  BUF_X1 U507 ( .A(n681), .Z(n375) );
  BUF_X1 U508 ( .A(n775), .Z(n376) );
  INV_X1 U509 ( .A(n712), .ZN(n450) );
  NAND2_X1 U510 ( .A1(n378), .A2(n377), .ZN(n667) );
  AND2_X1 U511 ( .A1(n714), .A2(G475), .ZN(n377) );
  NAND2_X1 U512 ( .A1(n443), .A2(n441), .ZN(n378) );
  NAND2_X1 U513 ( .A1(n443), .A2(n441), .ZN(n451) );
  NAND2_X1 U514 ( .A1(n442), .A2(n373), .ZN(n441) );
  NAND2_X1 U515 ( .A1(n451), .A2(n714), .ZN(n380) );
  NAND2_X1 U516 ( .A1(n760), .A2(n777), .ZN(n648) );
  XNOR2_X2 U517 ( .A(n555), .B(KEYINPUT31), .ZN(n705) );
  XNOR2_X2 U518 ( .A(n487), .B(KEYINPUT0), .ZN(n568) );
  NAND2_X1 U519 ( .A1(n384), .A2(n369), .ZN(n456) );
  INV_X1 U520 ( .A(n719), .ZN(n384) );
  XNOR2_X2 U521 ( .A(n567), .B(n566), .ZN(n719) );
  NAND2_X1 U522 ( .A1(n586), .A2(n585), .ZN(n385) );
  NAND2_X1 U523 ( .A1(n681), .A2(G469), .ZN(n454) );
  XNOR2_X1 U524 ( .A(n471), .B(n472), .ZN(n473) );
  NAND2_X1 U525 ( .A1(n394), .A2(n397), .ZN(n423) );
  NOR2_X2 U526 ( .A1(n582), .A2(KEYINPUT44), .ZN(n584) );
  XNOR2_X1 U527 ( .A(n391), .B(n474), .ZN(n652) );
  XNOR2_X1 U528 ( .A(n473), .B(n518), .ZN(n391) );
  XNOR2_X2 U529 ( .A(n392), .B(n514), .ZN(n440) );
  XNOR2_X1 U530 ( .A(n392), .B(n502), .ZN(n431) );
  XNOR2_X2 U531 ( .A(n506), .B(G134), .ZN(n392) );
  AND2_X1 U532 ( .A1(n393), .A2(n399), .ZN(n396) );
  NAND2_X1 U533 ( .A1(n403), .A2(n401), .ZN(n393) );
  XNOR2_X2 U534 ( .A(n635), .B(n371), .ZN(n403) );
  XNOR2_X1 U535 ( .A(n625), .B(KEYINPUT46), .ZN(n397) );
  INV_X1 U536 ( .A(n403), .ZN(n398) );
  AND2_X1 U537 ( .A1(n359), .A2(n402), .ZN(n401) );
  INV_X1 U538 ( .A(n404), .ZN(n410) );
  NAND2_X1 U539 ( .A1(n410), .A2(n411), .ZN(n619) );
  NAND2_X1 U540 ( .A1(n410), .A2(n406), .ZN(n405) );
  NAND2_X1 U541 ( .A1(n645), .A2(n627), .ZN(n412) );
  NAND2_X1 U542 ( .A1(n415), .A2(n414), .ZN(n413) );
  INV_X1 U543 ( .A(n623), .ZN(n415) );
  NOR2_X1 U544 ( .A1(n419), .A2(n367), .ZN(n416) );
  NOR2_X1 U545 ( .A1(n419), .A2(n418), .ZN(n417) );
  INV_X1 U546 ( .A(n560), .ZN(n570) );
  XNOR2_X2 U547 ( .A(n424), .B(KEYINPUT99), .ZN(n627) );
  NAND2_X1 U548 ( .A1(n571), .A2(n560), .ZN(n424) );
  INV_X1 U549 ( .A(n613), .ZN(n642) );
  INV_X1 U550 ( .A(n432), .ZN(n632) );
  NAND2_X1 U551 ( .A1(n598), .A2(n486), .ZN(n487) );
  INV_X1 U552 ( .A(n720), .ZN(n433) );
  XNOR2_X1 U553 ( .A(n440), .B(n526), .ZN(n527) );
  INV_X1 U554 ( .A(n648), .ZN(n442) );
  AND2_X2 U555 ( .A1(n448), .A2(n444), .ZN(n443) );
  NAND2_X1 U556 ( .A1(n648), .A2(n449), .ZN(n448) );
  NAND2_X1 U557 ( .A1(n719), .A2(n569), .ZN(n455) );
  NAND2_X2 U558 ( .A1(n457), .A2(n456), .ZN(n574) );
  NAND2_X1 U559 ( .A1(n568), .A2(n569), .ZN(n458) );
  AND2_X1 U560 ( .A1(n619), .A2(n607), .ZN(n608) );
  AND2_X1 U561 ( .A1(n359), .A2(n575), .ZN(n576) );
  INV_X1 U562 ( .A(KEYINPUT48), .ZN(n636) );
  BUF_X1 U563 ( .A(n719), .Z(n751) );
  INV_X1 U564 ( .A(KEYINPUT36), .ZN(n634) );
  XNOR2_X1 U565 ( .A(n535), .B(n534), .ZN(n536) );
  OR2_X1 U566 ( .A1(n778), .A2(G952), .ZN(n674) );
  INV_X1 U567 ( .A(G119), .ZN(n460) );
  NAND2_X1 U568 ( .A1(G113), .A2(n460), .ZN(n463) );
  NAND2_X1 U569 ( .A1(n461), .A2(G119), .ZN(n462) );
  XNOR2_X1 U570 ( .A(KEYINPUT4), .B(n768), .ZN(n474) );
  XNOR2_X1 U571 ( .A(n362), .B(n464), .ZN(n766) );
  XOR2_X1 U572 ( .A(n488), .B(KEYINPUT17), .Z(n472) );
  XNOR2_X2 U573 ( .A(G128), .B(KEYINPUT77), .ZN(n468) );
  INV_X1 U574 ( .A(G143), .ZN(n467) );
  XNOR2_X2 U575 ( .A(n468), .B(n467), .ZN(n506) );
  NAND2_X1 U576 ( .A1(G224), .A2(n778), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n469), .B(KEYINPUT18), .ZN(n470) );
  XNOR2_X1 U578 ( .A(n506), .B(n470), .ZN(n471) );
  XNOR2_X1 U579 ( .A(G902), .B(KEYINPUT15), .ZN(n508) );
  NOR2_X1 U580 ( .A1(n652), .A2(n649), .ZN(n476) );
  OR2_X1 U581 ( .A1(G237), .A2(G902), .ZN(n477) );
  NAND2_X1 U582 ( .A1(G210), .A2(n477), .ZN(n475) );
  XNOR2_X1 U583 ( .A(n476), .B(n475), .ZN(n604) );
  NAND2_X1 U584 ( .A1(G214), .A2(n477), .ZN(n478) );
  XNOR2_X1 U585 ( .A(KEYINPUT85), .B(n478), .ZN(n720) );
  NAND2_X1 U586 ( .A1(G234), .A2(G237), .ZN(n479) );
  XNOR2_X1 U587 ( .A(n479), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U588 ( .A1(G952), .A2(n481), .ZN(n750) );
  NOR2_X1 U589 ( .A1(G953), .A2(n750), .ZN(n480) );
  XNOR2_X1 U590 ( .A(KEYINPUT86), .B(n480), .ZN(n589) );
  NAND2_X1 U591 ( .A1(n481), .A2(G902), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n482), .B(KEYINPUT88), .ZN(n590) );
  NOR2_X1 U593 ( .A1(G898), .A2(n778), .ZN(n483) );
  XNOR2_X1 U594 ( .A(KEYINPUT87), .B(n483), .ZN(n769) );
  NOR2_X1 U595 ( .A1(n590), .A2(n769), .ZN(n484) );
  NOR2_X1 U596 ( .A1(n589), .A2(n484), .ZN(n485) );
  XNOR2_X1 U597 ( .A(KEYINPUT89), .B(n485), .ZN(n486) );
  XNOR2_X1 U598 ( .A(n490), .B(n489), .ZN(n492) );
  XOR2_X1 U599 ( .A(n494), .B(G113), .Z(n499) );
  XNOR2_X1 U600 ( .A(n495), .B(KEYINPUT76), .ZN(n521) );
  NAND2_X1 U601 ( .A1(n521), .A2(G214), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n513), .B(G143), .ZN(n496) );
  XNOR2_X1 U603 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U604 ( .A(n499), .B(n498), .ZN(n665) );
  XNOR2_X1 U605 ( .A(KEYINPUT13), .B(G475), .ZN(n500) );
  NAND2_X1 U606 ( .A1(G217), .A2(n538), .ZN(n502) );
  XNOR2_X1 U607 ( .A(G107), .B(n504), .ZN(n505) );
  INV_X1 U608 ( .A(G902), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n676), .A2(n543), .ZN(n507) );
  NOR2_X1 U610 ( .A1(n571), .A2(n570), .ZN(n722) );
  NAND2_X1 U611 ( .A1(G234), .A2(n508), .ZN(n509) );
  XNOR2_X1 U612 ( .A(KEYINPUT20), .B(n509), .ZN(n544) );
  NAND2_X1 U613 ( .A1(G221), .A2(n544), .ZN(n511) );
  XNOR2_X1 U614 ( .A(KEYINPUT21), .B(KEYINPUT95), .ZN(n510) );
  XNOR2_X1 U615 ( .A(n511), .B(n510), .ZN(n734) );
  INV_X1 U616 ( .A(n734), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U618 ( .A1(G227), .A2(n778), .ZN(n515) );
  XNOR2_X1 U619 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U621 ( .A(n520), .B(G116), .Z(n523) );
  NAND2_X1 U622 ( .A1(G210), .A2(n521), .ZN(n522) );
  XNOR2_X1 U623 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U624 ( .A(n524), .B(KEYINPUT5), .Z(n528) );
  XNOR2_X1 U625 ( .A(n525), .B(G146), .ZN(n526) );
  INV_X1 U626 ( .A(G472), .ZN(n659) );
  INV_X1 U627 ( .A(KEYINPUT6), .ZN(n529) );
  XNOR2_X1 U628 ( .A(n738), .B(n529), .ZN(n575) );
  INV_X1 U629 ( .A(n575), .ZN(n630) );
  OR2_X1 U630 ( .A1(n359), .A2(n630), .ZN(n530) );
  XNOR2_X1 U631 ( .A(n531), .B(KEYINPUT82), .ZN(n549) );
  XOR2_X1 U632 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n533) );
  XNOR2_X1 U633 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U634 ( .A(KEYINPUT91), .B(KEYINPUT94), .Z(n534) );
  XNOR2_X1 U635 ( .A(n773), .B(n536), .ZN(n542) );
  XNOR2_X1 U636 ( .A(n537), .B(n459), .ZN(n540) );
  NAND2_X1 U637 ( .A1(n538), .A2(G221), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U639 ( .A(n542), .B(n541), .ZN(n673) );
  NAND2_X1 U640 ( .A1(n673), .A2(n543), .ZN(n547) );
  NAND2_X1 U641 ( .A1(G217), .A2(n544), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n545), .B(KEYINPUT25), .ZN(n546) );
  XNOR2_X1 U643 ( .A(n547), .B(n546), .ZN(n588) );
  INV_X1 U644 ( .A(KEYINPUT102), .ZN(n548) );
  NAND2_X1 U645 ( .A1(n549), .A2(n735), .ZN(n550) );
  XNOR2_X1 U646 ( .A(n550), .B(KEYINPUT103), .ZN(n791) );
  INV_X1 U647 ( .A(n731), .ZN(n552) );
  INV_X1 U648 ( .A(KEYINPUT74), .ZN(n553) );
  XNOR2_X2 U649 ( .A(n554), .B(n553), .ZN(n564) );
  INV_X1 U650 ( .A(n738), .ZN(n556) );
  NAND2_X1 U651 ( .A1(n564), .A2(n556), .ZN(n741) );
  OR2_X1 U652 ( .A1(n568), .A2(n741), .ZN(n555) );
  NOR2_X1 U653 ( .A1(n556), .A2(n731), .ZN(n557) );
  NAND2_X1 U654 ( .A1(n557), .A2(n619), .ZN(n558) );
  NOR2_X1 U655 ( .A1(n568), .A2(n558), .ZN(n687) );
  NOR2_X1 U656 ( .A1(n571), .A2(n560), .ZN(n559) );
  XNOR2_X1 U657 ( .A(KEYINPUT100), .B(n559), .ZN(n706) );
  NOR2_X1 U658 ( .A1(n706), .A2(n627), .ZN(n587) );
  NOR2_X1 U659 ( .A1(n561), .A2(n587), .ZN(n562) );
  XOR2_X1 U660 ( .A(KEYINPUT101), .B(n562), .Z(n563) );
  NOR2_X1 U661 ( .A1(n791), .A2(n563), .ZN(n580) );
  XNOR2_X1 U662 ( .A(n564), .B(KEYINPUT104), .ZN(n565) );
  NAND2_X1 U663 ( .A1(n565), .A2(n630), .ZN(n567) );
  XNOR2_X1 U664 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n566) );
  NAND2_X1 U665 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U666 ( .A(n572), .B(KEYINPUT105), .ZN(n610) );
  NAND2_X1 U667 ( .A1(n582), .A2(KEYINPUT44), .ZN(n579) );
  NAND2_X1 U668 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U669 ( .A(n581), .B(KEYINPUT83), .ZN(n586) );
  XNOR2_X1 U670 ( .A(n584), .B(n583), .ZN(n585) );
  INV_X1 U671 ( .A(n587), .ZN(n724) );
  XOR2_X1 U672 ( .A(KEYINPUT47), .B(n724), .Z(n603) );
  INV_X1 U673 ( .A(KEYINPUT47), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT28), .B(KEYINPUT108), .ZN(n597) );
  AND2_X1 U675 ( .A1(n734), .A2(n588), .ZN(n595) );
  INV_X1 U676 ( .A(n589), .ZN(n593) );
  NOR2_X1 U677 ( .A1(n590), .A2(G900), .ZN(n591) );
  NAND2_X1 U678 ( .A1(G953), .A2(n591), .ZN(n592) );
  NAND2_X1 U679 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U680 ( .A(KEYINPUT78), .B(n594), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n595), .A2(n607), .ZN(n629) );
  NOR2_X1 U682 ( .A1(n629), .A2(n738), .ZN(n596) );
  XNOR2_X1 U683 ( .A(n597), .B(n596), .ZN(n620) );
  NAND2_X1 U684 ( .A1(n598), .A2(n620), .ZN(n600) );
  INV_X1 U685 ( .A(n619), .ZN(n599) );
  OR2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n698) );
  NAND2_X1 U687 ( .A1(n601), .A2(n698), .ZN(n602) );
  NAND2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n614) );
  BUF_X1 U689 ( .A(n604), .Z(n613) );
  XOR2_X1 U690 ( .A(KEYINPUT30), .B(n605), .Z(n606) );
  NOR2_X1 U691 ( .A1(n606), .A2(n731), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n623) );
  INV_X1 U693 ( .A(n610), .ZN(n611) );
  NOR2_X1 U694 ( .A1(n623), .A2(n611), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n697) );
  NAND2_X1 U696 ( .A1(n614), .A2(n697), .ZN(n617) );
  NAND2_X1 U697 ( .A1(KEYINPUT47), .A2(n698), .ZN(n615) );
  XNOR2_X1 U698 ( .A(KEYINPUT79), .B(n615), .ZN(n616) );
  NOR2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n720), .A2(n721), .ZN(n725) );
  NAND2_X1 U701 ( .A1(n725), .A2(n722), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U703 ( .A(KEYINPUT42), .B(n622), .ZN(n789) );
  XNOR2_X1 U704 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n624) );
  NOR2_X1 U705 ( .A1(n789), .A2(n786), .ZN(n625) );
  INV_X1 U706 ( .A(KEYINPUT106), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n635) );
  INV_X1 U708 ( .A(n359), .ZN(n732) );
  INV_X1 U709 ( .A(n637), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n638), .A2(n433), .ZN(n640) );
  OR2_X1 U711 ( .A1(n640), .A2(n359), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n641), .B(KEYINPUT43), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n644), .B(KEYINPUT107), .ZN(n787) );
  NAND2_X1 U715 ( .A1(n645), .A2(n706), .ZN(n710) );
  INV_X1 U716 ( .A(n710), .ZN(n646) );
  NOR2_X1 U717 ( .A1(n787), .A2(n646), .ZN(n647) );
  INV_X1 U718 ( .A(KEYINPUT2), .ZN(n711) );
  INV_X1 U719 ( .A(KEYINPUT64), .ZN(n650) );
  INV_X1 U720 ( .A(n760), .ZN(n712) );
  INV_X1 U721 ( .A(G210), .ZN(n651) );
  NOR2_X1 U722 ( .A1(n380), .A2(n651), .ZN(n655) );
  XOR2_X1 U723 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n653) );
  XNOR2_X1 U724 ( .A(n652), .B(n653), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n656), .A2(n674), .ZN(n658) );
  INV_X1 U727 ( .A(KEYINPUT56), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(G51) );
  NOR2_X1 U729 ( .A1(n380), .A2(n659), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT62), .B(n660), .Z(n661) );
  XNOR2_X1 U731 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n663), .A2(n674), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U734 ( .A(n665), .B(KEYINPUT59), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n668), .A2(n674), .ZN(n670) );
  INV_X1 U737 ( .A(KEYINPUT60), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n670), .B(n669), .ZN(G60) );
  XNOR2_X1 U739 ( .A(n671), .B(G122), .ZN(G24) );
  AND2_X1 U740 ( .A1(n379), .A2(G217), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n673), .B(n672), .ZN(n675) );
  INV_X1 U742 ( .A(n674), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n675), .A2(n684), .ZN(G66) );
  NAND2_X1 U744 ( .A1(n379), .A2(G478), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n676), .B(KEYINPUT121), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n679), .A2(n684), .ZN(G63) );
  NAND2_X1 U748 ( .A1(n379), .A2(G469), .ZN(n683) );
  XOR2_X1 U749 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n680) );
  XNOR2_X1 U750 ( .A(n375), .B(n680), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(n685) );
  NOR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(G54) );
  INV_X1 U753 ( .A(n699), .ZN(n702) );
  NAND2_X1 U754 ( .A1(n702), .A2(n687), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(G104), .ZN(G6) );
  XOR2_X1 U756 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U757 ( .A1(n687), .A2(n706), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n689), .B(n688), .ZN(n691) );
  XOR2_X1 U759 ( .A(G107), .B(KEYINPUT27), .Z(n690) );
  XNOR2_X1 U760 ( .A(n691), .B(n690), .ZN(G9) );
  XOR2_X1 U761 ( .A(G110), .B(n692), .Z(n693) );
  XNOR2_X1 U762 ( .A(KEYINPUT114), .B(n693), .ZN(G12) );
  INV_X1 U763 ( .A(n706), .ZN(n694) );
  NOR2_X1 U764 ( .A1(n694), .A2(n698), .ZN(n696) );
  XNOR2_X1 U765 ( .A(G128), .B(KEYINPUT29), .ZN(n695) );
  XNOR2_X1 U766 ( .A(n696), .B(n695), .ZN(G30) );
  XNOR2_X1 U767 ( .A(G143), .B(n697), .ZN(G45) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U769 ( .A(G146), .B(KEYINPUT115), .ZN(n700) );
  XNOR2_X1 U770 ( .A(n701), .B(n700), .ZN(G48) );
  NAND2_X1 U771 ( .A1(n702), .A2(n705), .ZN(n703) );
  XNOR2_X1 U772 ( .A(n703), .B(KEYINPUT116), .ZN(n704) );
  XNOR2_X1 U773 ( .A(G113), .B(n704), .ZN(G15) );
  NAND2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U775 ( .A(n707), .B(G116), .ZN(G18) );
  XNOR2_X1 U776 ( .A(n370), .B(G125), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n708), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U778 ( .A(G134), .B(KEYINPUT117), .Z(n709) );
  XNOR2_X1 U779 ( .A(n710), .B(n709), .ZN(G36) );
  NAND2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U781 ( .A(n713), .B(KEYINPUT80), .ZN(n718) );
  INV_X1 U782 ( .A(n714), .ZN(n716) );
  NOR2_X1 U783 ( .A1(n777), .A2(KEYINPUT2), .ZN(n715) );
  NOR2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n758) );
  NAND2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n728) );
  NAND2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U789 ( .A(KEYINPUT118), .B(n726), .ZN(n727) );
  NAND2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U791 ( .A1(n384), .A2(n729), .ZN(n730) );
  XNOR2_X1 U792 ( .A(n730), .B(KEYINPUT119), .ZN(n747) );
  NAND2_X1 U793 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U794 ( .A(KEYINPUT50), .B(n733), .Z(n740) );
  NOR2_X1 U795 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U796 ( .A(n736), .B(KEYINPUT49), .ZN(n737) );
  NAND2_X1 U797 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U798 ( .A1(n740), .A2(n739), .ZN(n743) );
  INV_X1 U799 ( .A(n741), .ZN(n742) );
  NOR2_X1 U800 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U801 ( .A(KEYINPUT51), .B(n744), .Z(n745) );
  NOR2_X1 U802 ( .A1(n752), .A2(n745), .ZN(n746) );
  NOR2_X1 U803 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U804 ( .A(n748), .B(KEYINPUT52), .ZN(n749) );
  NOR2_X1 U805 ( .A1(n750), .A2(n749), .ZN(n754) );
  NOR2_X1 U806 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U807 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U808 ( .A(KEYINPUT120), .B(n755), .Z(n756) );
  NOR2_X1 U809 ( .A1(G953), .A2(n756), .ZN(n757) );
  NAND2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U811 ( .A(KEYINPUT53), .B(n759), .Z(G75) );
  NAND2_X1 U812 ( .A1(n450), .A2(n778), .ZN(n765) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n761) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n761), .ZN(n762) );
  NAND2_X1 U815 ( .A1(n762), .A2(G898), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n763), .B(KEYINPUT122), .ZN(n764) );
  NAND2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n772) );
  XOR2_X1 U818 ( .A(G101), .B(n766), .Z(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(n770) );
  NAND2_X1 U820 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U821 ( .A(n772), .B(n771), .Z(G69) );
  XOR2_X1 U822 ( .A(n773), .B(KEYINPUT123), .Z(n774) );
  XNOR2_X1 U823 ( .A(n376), .B(n774), .ZN(n780) );
  XOR2_X1 U824 ( .A(KEYINPUT124), .B(n780), .Z(n776) );
  XNOR2_X1 U825 ( .A(n777), .B(n776), .ZN(n779) );
  NAND2_X1 U826 ( .A1(n779), .A2(n778), .ZN(n784) );
  XNOR2_X1 U827 ( .A(n780), .B(G227), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n781), .A2(G900), .ZN(n782) );
  NAND2_X1 U829 ( .A1(n782), .A2(G953), .ZN(n783) );
  NAND2_X1 U830 ( .A1(n784), .A2(n783), .ZN(G72) );
  XOR2_X1 U831 ( .A(G131), .B(KEYINPUT126), .Z(n785) );
  XNOR2_X1 U832 ( .A(n786), .B(n785), .ZN(G33) );
  XOR2_X1 U833 ( .A(G140), .B(n787), .Z(G42) );
  XNOR2_X1 U834 ( .A(n788), .B(G119), .ZN(G21) );
  XNOR2_X1 U835 ( .A(G137), .B(KEYINPUT125), .ZN(n790) );
  XNOR2_X1 U836 ( .A(n790), .B(n789), .ZN(G39) );
  XOR2_X1 U837 ( .A(n791), .B(G101), .Z(n792) );
  XNOR2_X1 U838 ( .A(KEYINPUT112), .B(n792), .ZN(G3) );
endmodule

