//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT86), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G43gat), .ZN(new_n207));
  AOI21_X1  g006(.A(G50gat), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT87), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G50gat), .ZN(new_n212));
  AOI21_X1  g011(.A(G43gat), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n203), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(G43gat), .A2(G50gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G43gat), .A2(G50gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT15), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(KEYINPUT85), .B(KEYINPUT15), .C1(new_n215), .C2(new_n216), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT14), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT88), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT88), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n214), .A2(new_n221), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n224), .A2(new_n226), .A3(new_n229), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n204), .A2(new_n209), .ZN(new_n235));
  NAND2_X1  g034(.A1(G43gat), .A2(G50gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n203), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n234), .A2(new_n237), .A3(KEYINPUT84), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT84), .B1(new_n234), .B2(new_n237), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G22gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G15gat), .ZN(new_n245));
  INV_X1    g044(.A(G15gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G22gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n245), .B2(new_n247), .ZN(new_n251));
  INV_X1    g050(.A(G1gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT16), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n250), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT89), .ZN(new_n257));
  AOI21_X1  g056(.A(G1gat), .B1(new_n257), .B2(new_n249), .ZN(new_n258));
  OAI21_X1  g057(.A(G8gat), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n252), .B1(new_n250), .B2(new_n251), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n257), .A2(new_n253), .A3(new_n249), .ZN(new_n261));
  INV_X1    g060(.A(G8gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n233), .A2(KEYINPUT17), .A3(new_n240), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n243), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G229gat), .A2(G233gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n259), .A2(new_n263), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT90), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n268), .A2(new_n241), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n268), .B2(new_n241), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n266), .B(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT92), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT18), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n272), .B2(new_n274), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n268), .A2(new_n241), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT90), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n268), .A2(new_n241), .A3(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(KEYINPUT18), .A3(new_n267), .A4(new_n266), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n270), .A2(new_n271), .B1(new_n241), .B2(new_n268), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n267), .B(KEYINPUT13), .Z(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G113gat), .B(G141gat), .ZN(new_n286));
  INV_X1    g085(.A(G197gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT11), .B(G169gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n290), .B(KEYINPUT12), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n282), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n202), .B1(new_n277), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n282), .A2(new_n285), .A3(new_n292), .ZN(new_n295));
  NOR4_X1   g094(.A1(new_n295), .A2(new_n275), .A3(new_n276), .A4(KEYINPUT93), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n274), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(new_n282), .A3(new_n285), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT91), .B1(new_n298), .B2(new_n291), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n298), .A2(KEYINPUT91), .A3(new_n291), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n294), .A2(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT94), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI221_X1 g102(.A(KEYINPUT94), .B1(new_n300), .B2(new_n299), .C1(new_n294), .C2(new_n296), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n307));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(G183gat), .A3(G190gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G183gat), .B(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n309), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT25), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n312), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(new_n316), .B2(new_n317), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT65), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n318), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n313), .B1(new_n312), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT64), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT64), .B(new_n313), .C1(new_n312), .C2(new_n327), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n325), .A2(KEYINPUT66), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT66), .B1(new_n325), .B2(new_n333), .ZN(new_n335));
  OAI221_X1 g134(.A(new_n321), .B1(new_n333), .B2(new_n325), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT28), .B1(new_n339), .B2(new_n338), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n339), .A2(KEYINPUT28), .A3(new_n338), .ZN(new_n341));
  OAI221_X1 g140(.A(new_n336), .B1(new_n337), .B2(new_n338), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n308), .B1(new_n332), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n332), .A2(new_n342), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n343), .B1(new_n346), .B2(new_n308), .ZN(new_n347));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348));
  AND2_X1   g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(KEYINPUT22), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G211gat), .B(G218gat), .Z(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT70), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n351), .A2(KEYINPUT69), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(KEYINPUT69), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(KEYINPUT71), .A3(new_n356), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n307), .B1(new_n347), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n343), .ZN(new_n363));
  INV_X1    g162(.A(new_n308), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n332), .B2(new_n342), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(new_n360), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(KEYINPUT72), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT73), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n365), .B2(new_n364), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n361), .B(new_n371), .C1(new_n347), .C2(new_n370), .ZN(new_n372));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  NAND3_X1  g174(.A1(new_n369), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT30), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n369), .A2(new_n378), .A3(new_n372), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n347), .A2(new_n361), .A3(new_n307), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT72), .B1(new_n366), .B2(new_n367), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n372), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT74), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n372), .ZN(new_n386));
  INV_X1    g185(.A(new_n375), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n389));
  XOR2_X1   g188(.A(G155gat), .B(G162gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G141gat), .B(G148gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(KEYINPUT2), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT75), .B(G162gat), .ZN(new_n395));
  INV_X1    g194(.A(G155gat), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT2), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n394), .B1(new_n393), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n392), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G127gat), .B(G134gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT67), .ZN(new_n403));
  NOR2_X1   g202(.A1(G113gat), .A2(G120gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(KEYINPUT1), .ZN(new_n405));
  NAND2_X1  g204(.A1(G113gat), .A2(G120gat), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n402), .A2(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT67), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n408), .A2(KEYINPUT67), .A3(new_n406), .A4(new_n405), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(new_n392), .C1(new_n399), .C2(new_n400), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n389), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n420), .A3(KEYINPUT4), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n413), .B1(new_n401), .B2(KEYINPUT3), .ZN(new_n422));
  INV_X1    g221(.A(new_n392), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n393), .A2(new_n397), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT76), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n425), .B2(new_n398), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT3), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n421), .B(new_n417), .C1(new_n422), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n415), .A2(KEYINPUT4), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n431), .A3(new_n412), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT77), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n419), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n412), .B1(new_n426), .B2(new_n427), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n427), .B2(new_n426), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n432), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n389), .A4(new_n417), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT0), .ZN(new_n441));
  XNOR2_X1  g240(.A(G57gat), .B(G85gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n434), .A2(new_n443), .A3(new_n438), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n380), .A2(new_n388), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT78), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT79), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n345), .B1(new_n401), .B2(KEYINPUT3), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n367), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n350), .A2(new_n351), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT29), .B1(new_n353), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n401), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT80), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n460), .A2(KEYINPUT80), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n454), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT3), .B1(new_n357), .B2(new_n345), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n457), .B(new_n465), .C1(new_n426), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT31), .B(G50gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n244), .ZN(new_n472));
  NAND2_X1  g271(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n471), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n468), .A2(new_n474), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n380), .A2(new_n388), .A3(KEYINPUT78), .A4(new_n450), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G15gat), .B(G43gat), .Z(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n344), .A2(new_n412), .ZN(new_n484));
  AND2_X1   g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n332), .A2(new_n413), .A3(new_n342), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT33), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n484), .B2(new_n486), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI211_X1 g291(.A(KEYINPUT34), .B(new_n485), .C1(new_n484), .C2(new_n486), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n496), .B1(new_n500), .B2(new_n494), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT36), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  AOI211_X1 g304(.A(KEYINPUT68), .B(new_n505), .C1(new_n499), .C2(new_n501), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n479), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT82), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n479), .A2(new_n507), .A3(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n380), .A2(new_n388), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n417), .B1(new_n436), .B2(new_n437), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT39), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n443), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT39), .B1(new_n416), .B2(new_n418), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  OR3_X1    g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n517), .B1(new_n516), .B2(new_n519), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n521), .A2(new_n445), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n512), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n475), .A2(new_n476), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n369), .A2(new_n525), .A3(new_n372), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n526), .A2(KEYINPUT38), .A3(new_n387), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n385), .A2(KEYINPUT37), .A3(new_n386), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n367), .B(new_n371), .C1(new_n347), .C2(new_n370), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n366), .B2(new_n361), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT83), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT83), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n526), .A2(new_n533), .A3(new_n387), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT38), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n527), .A2(new_n528), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n448), .A2(new_n449), .A3(new_n376), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n523), .B(new_n524), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n510), .A2(new_n511), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n451), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542));
  INV_X1    g341(.A(new_n502), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n524), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n499), .A3(new_n501), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n545), .B1(new_n453), .B2(new_n478), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n546), .B2(new_n542), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n306), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  OR2_X1    g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(KEYINPUT96), .A3(new_n549), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556));
  AND2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(KEYINPUT95), .A2(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(G64gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n552), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n554), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n554), .A3(new_n559), .A4(new_n555), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n553), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g372(.A(G127gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n268), .B1(new_n570), .B2(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n573), .B(G127gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(new_n396), .ZN(new_n583));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n577), .A2(new_n580), .A3(new_n585), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT8), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT99), .B(G92gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n591), .B(new_n593), .C1(G85gat), .C2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n594), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n592), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n591), .A4(new_n593), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n243), .A2(new_n265), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  AND2_X1   g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n605), .A2(new_n241), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G190gat), .B(G218gat), .Z(new_n609));
  AND2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT98), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n612), .A2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G230gat), .ZN(new_n621));
  INV_X1    g420(.A(G233gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n569), .A2(new_n603), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n565), .A2(new_n559), .A3(new_n555), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT97), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n567), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(new_n553), .A3(new_n597), .A4(new_n602), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n570), .A2(new_n605), .A3(KEYINPUT10), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n623), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n624), .A2(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n623), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n635), .A3(new_n639), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n589), .A2(new_n620), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n548), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n450), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT101), .B(G1gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1324gat));
  XNOR2_X1  g451(.A(KEYINPUT16), .B(G8gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n548), .A2(new_n512), .A3(new_n646), .A4(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n658));
  INV_X1    g457(.A(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(new_n661), .A3(new_n656), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n548), .A2(new_n512), .A3(new_n646), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G8gat), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n658), .A2(new_n660), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT103), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n659), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n663), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n662), .A4(new_n658), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(G1325gat));
  OAI21_X1  g469(.A(new_n246), .B1(new_n647), .B2(new_n502), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT104), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n647), .A2(new_n246), .A3(new_n507), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n647), .A2(new_n524), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n620), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n540), .B2(new_n547), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n539), .A2(new_n479), .A3(new_n507), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n547), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT44), .B1(new_n683), .B2(new_n619), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n589), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n644), .ZN(new_n687));
  INV_X1    g486(.A(new_n299), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n298), .A2(KEYINPUT91), .A3(new_n291), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n297), .A2(KEYINPUT92), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT93), .B1(new_n692), .B2(new_n295), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n277), .A2(new_n202), .A3(new_n293), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n688), .A2(new_n689), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n685), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n649), .ZN(new_n698));
  INV_X1    g497(.A(new_n649), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n687), .A2(new_n620), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n548), .A2(new_n222), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n698), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n698), .A2(KEYINPUT105), .A3(new_n703), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1328gat));
  AND2_X1   g508(.A1(new_n548), .A2(new_n700), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n223), .A3(new_n512), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n712));
  INV_X1    g511(.A(new_n512), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n697), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n205), .A2(new_n207), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n697), .B2(new_n507), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n717), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n710), .A2(new_n721), .A3(new_n543), .ZN(new_n722));
  INV_X1    g521(.A(new_n507), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n685), .A2(new_n723), .A3(new_n696), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n718), .B(new_n722), .C1(new_n719), .C2(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1330gat));
  NAND2_X1  g528(.A1(new_n210), .A2(new_n212), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n697), .B2(new_n524), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n524), .A2(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n710), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n731), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n731), .B2(new_n734), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  NAND3_X1  g537(.A1(new_n589), .A2(new_n620), .A3(new_n643), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n301), .B(new_n739), .C1(new_n547), .C2(new_n682), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n699), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n512), .B1(new_n743), .B2(new_n563), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n563), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n740), .A2(new_n749), .A3(new_n543), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n740), .A2(new_n723), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n749), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g552(.A1(new_n740), .A2(new_n477), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n589), .A2(new_n301), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n643), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n685), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n649), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n683), .A2(new_n619), .A3(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n619), .A4(new_n756), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n699), .A2(new_n599), .A3(new_n643), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  NAND2_X1  g567(.A1(new_n540), .A2(new_n547), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n679), .ZN(new_n770));
  INV_X1    g569(.A(new_n684), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n512), .A4(new_n758), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n594), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n713), .A2(G92gat), .A3(new_n644), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n765), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n774), .B(KEYINPUT109), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n765), .A2(new_n778), .ZN(new_n779));
  AOI211_X1 g578(.A(KEYINPUT110), .B(new_n777), .C1(new_n773), .C2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n681), .A2(new_n684), .A3(new_n713), .A4(new_n757), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n782), .B2(new_n598), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n781), .B1(new_n783), .B2(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n776), .B1(new_n780), .B2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n759), .B2(new_n507), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n502), .A2(G99gat), .A3(new_n644), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n766), .B2(new_n787), .ZN(G1338gat));
  NOR3_X1   g587(.A1(new_n524), .A2(G106gat), .A3(new_n644), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT111), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n765), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n685), .A2(new_n477), .A3(new_n758), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n793), .A2(G106gat), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT53), .B1(new_n799), .B2(new_n791), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1339gat));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n630), .A2(new_n631), .A3(new_n623), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n632), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n630), .A2(new_n631), .ZN(new_n807));
  INV_X1    g606(.A(new_n623), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n640), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n642), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n630), .A2(new_n631), .A3(new_n623), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n639), .B1(new_n632), .B2(new_n805), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT113), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n814), .A2(new_n815), .A3(new_n818), .A4(KEYINPUT55), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n812), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n281), .A2(new_n266), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n821), .A2(new_n267), .B1(new_n283), .B2(new_n284), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n290), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n693), .B2(new_n694), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n820), .B(new_n619), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n823), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n294), .B2(new_n296), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n301), .A2(new_n820), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n827), .B(new_n643), .C1(new_n294), .C2(new_n296), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n619), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n802), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n642), .A3(new_n811), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n695), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n620), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n825), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n619), .A4(new_n820), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n841), .A3(KEYINPUT115), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n834), .A2(new_n686), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n645), .A2(new_n301), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n649), .A2(new_n545), .A3(new_n512), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(G113gat), .A3(new_n695), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n301), .A2(new_n820), .B1(new_n824), .B2(new_n643), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n850), .A2(new_n619), .B1(new_n826), .B2(new_n829), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n589), .B1(new_n851), .B2(new_n802), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n844), .B1(new_n852), .B2(new_n842), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n853), .B2(new_n477), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n855), .A3(new_n524), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n649), .A2(new_n502), .A3(new_n512), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n305), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n849), .B1(new_n859), .B2(G113gat), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT117), .ZN(G1340gat));
  NOR3_X1   g660(.A1(new_n848), .A2(G120gat), .A3(new_n644), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n643), .A3(new_n858), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(G120gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT118), .ZN(G1341gat));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n857), .A2(new_n858), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n686), .A2(new_n574), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n858), .A4(new_n868), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n574), .B1(new_n848), .B2(new_n686), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1342gat));
  NOR3_X1   g672(.A1(new_n848), .A2(G134gat), .A3(new_n620), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n867), .B2(new_n620), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1343gat));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n846), .A2(new_n477), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n507), .A2(new_n699), .A3(new_n713), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(G141gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n305), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n524), .A2(new_n884), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n836), .B1(new_n303), .B2(new_n304), .ZN(new_n887));
  INV_X1    g686(.A(new_n832), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n620), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n589), .B1(new_n889), .B2(new_n841), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n890), .B2(new_n844), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n880), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n305), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n878), .B(new_n883), .C1(new_n893), .C2(new_n882), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n301), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n896), .A3(G141gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT58), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT120), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(G141gat), .B2(new_n895), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n894), .B1(new_n898), .B2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(G148gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n881), .A2(new_n902), .A3(new_n643), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n902), .C1(new_n892), .C2(new_n643), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n645), .A2(new_n305), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n477), .B1(new_n890), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n884), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  INV_X1    g708(.A(new_n886), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n853), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n846), .A2(KEYINPUT122), .A3(new_n886), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n880), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n643), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n905), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n903), .B1(new_n904), .B2(new_n916), .ZN(G1345gat));
  NAND3_X1  g716(.A1(new_n881), .A2(new_n396), .A3(new_n589), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n892), .A2(new_n589), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n396), .ZN(G1346gat));
  NAND3_X1  g719(.A1(new_n881), .A2(new_n395), .A3(new_n619), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n892), .A2(new_n619), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n395), .ZN(G1347gat));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n853), .B2(new_n699), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n846), .A2(new_n925), .A3(new_n649), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n545), .A2(new_n713), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n301), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n649), .A2(new_n512), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT124), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n543), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n932), .B1(new_n854), .B2(new_n856), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n306), .A2(new_n314), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n929), .A2(new_n314), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  AND2_X1   g734(.A1(new_n933), .A2(new_n643), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n927), .A2(new_n928), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n643), .A2(new_n315), .ZN(new_n938));
  OAI22_X1  g737(.A1(new_n936), .A2(new_n315), .B1(new_n937), .B2(new_n938), .ZN(G1349gat));
  NAND4_X1  g738(.A1(new_n927), .A2(new_n339), .A3(new_n589), .A4(new_n928), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n933), .A2(new_n589), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n337), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n944), .B(new_n940), .C1(new_n941), .C2(new_n337), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1350gat));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n933), .A2(new_n619), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(G190gat), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT61), .B(new_n338), .C1(new_n933), .C2(new_n619), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n619), .A2(new_n338), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n949), .A2(new_n950), .B1(new_n937), .B2(new_n951), .ZN(G1351gat));
  NOR3_X1   g751(.A1(new_n723), .A2(new_n524), .A3(new_n713), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n927), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n301), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n931), .A2(new_n507), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n913), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n959), .A2(new_n287), .A3(new_n306), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n955), .A2(new_n960), .ZN(G1352gat));
  INV_X1    g760(.A(G204gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n954), .A2(new_n962), .A3(new_n643), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n959), .B2(new_n644), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n913), .A2(new_n589), .A3(new_n958), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G211gat), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(KEYINPUT126), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n686), .A2(G211gat), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n974), .A2(new_n975), .B1(new_n954), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n973), .A2(new_n977), .ZN(G1354gat));
  OAI21_X1  g777(.A(G218gat), .B1(new_n959), .B2(new_n620), .ZN(new_n979));
  INV_X1    g778(.A(G218gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n954), .A2(new_n980), .A3(new_n619), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1355gat));
endmodule


