

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XNOR2_X1 U323 ( .A(n393), .B(n392), .ZN(n531) );
  XNOR2_X1 U324 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n392) );
  XNOR2_X1 U325 ( .A(n316), .B(n315), .ZN(n320) );
  XNOR2_X1 U326 ( .A(n440), .B(n314), .ZN(n315) );
  NOR2_X1 U327 ( .A1(n470), .A2(n571), .ZN(n433) );
  XNOR2_X1 U328 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n388) );
  XNOR2_X1 U329 ( .A(n318), .B(n317), .ZN(n352) );
  INV_X1 U330 ( .A(KEYINPUT67), .ZN(n321) );
  NAND2_X1 U331 ( .A1(n531), .A2(n467), .ZN(n412) );
  XNOR2_X1 U332 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U333 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U334 ( .A(n363), .B(n362), .ZN(n558) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(n566) );
  XOR2_X1 U336 ( .A(n470), .B(KEYINPUT28), .Z(n534) );
  XNOR2_X1 U337 ( .A(n456), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U338 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  INV_X1 U339 ( .A(KEYINPUT121), .ZN(n452) );
  XOR2_X1 U340 ( .A(G50GAT), .B(G162GAT), .Z(n336) );
  XNOR2_X1 U341 ( .A(G106GAT), .B(G204GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n291), .B(G148GAT), .ZN(n309) );
  XOR2_X1 U343 ( .A(n336), .B(n309), .Z(n293) );
  NAND2_X1 U344 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U346 ( .A(n294), .B(KEYINPUT88), .Z(n296) );
  XOR2_X1 U347 ( .A(G22GAT), .B(G155GAT), .Z(n349) );
  XNOR2_X1 U348 ( .A(n349), .B(KEYINPUT87), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U350 ( .A(G78GAT), .B(KEYINPUT24), .Z(n298) );
  XNOR2_X1 U351 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(n300), .B(n299), .Z(n306) );
  XOR2_X1 U354 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n302) );
  XNOR2_X1 U355 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n416) );
  XOR2_X1 U357 ( .A(G211GAT), .B(KEYINPUT21), .Z(n304) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(G218GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n400) );
  XNOR2_X1 U360 ( .A(n416), .B(n400), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n470) );
  XOR2_X1 U362 ( .A(KEYINPUT31), .B(KEYINPUT68), .Z(n308) );
  XNOR2_X1 U363 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n326) );
  NAND2_X1 U365 ( .A1(n309), .A2(KEYINPUT32), .ZN(n313) );
  INV_X1 U366 ( .A(n309), .ZN(n311) );
  INV_X1 U367 ( .A(KEYINPUT32), .ZN(n310) );
  NAND2_X1 U368 ( .A1(n311), .A2(n310), .ZN(n312) );
  NAND2_X1 U369 ( .A1(n313), .A2(n312), .ZN(n316) );
  XOR2_X1 U370 ( .A(G176GAT), .B(G120GAT), .Z(n440) );
  AND2_X1 U371 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XOR2_X1 U372 ( .A(KEYINPUT13), .B(G57GAT), .Z(n318) );
  XNOR2_X1 U373 ( .A(G71GAT), .B(G78GAT), .ZN(n317) );
  XOR2_X1 U374 ( .A(G99GAT), .B(G85GAT), .Z(n331) );
  XOR2_X1 U375 ( .A(n352), .B(n331), .Z(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U377 ( .A(G92GAT), .B(G64GAT), .Z(n405) );
  XNOR2_X1 U378 ( .A(n405), .B(KEYINPUT33), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n382) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n328) );
  XNOR2_X1 U381 ( .A(G218GAT), .B(G106GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n335) );
  XOR2_X1 U383 ( .A(G29GAT), .B(G36GAT), .Z(n330) );
  XNOR2_X1 U384 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n366) );
  XOR2_X1 U386 ( .A(n331), .B(n366), .Z(n333) );
  NAND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U389 ( .A(n335), .B(n334), .Z(n338) );
  XOR2_X1 U390 ( .A(G43GAT), .B(G134GAT), .Z(n446) );
  XNOR2_X1 U391 ( .A(n446), .B(n336), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U393 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n340) );
  XNOR2_X1 U394 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U396 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n342) );
  XNOR2_X1 U397 ( .A(G190GAT), .B(G92GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U399 ( .A(n344), .B(n343), .Z(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n562) );
  XNOR2_X1 U401 ( .A(KEYINPUT36), .B(n562), .ZN(n586) );
  XOR2_X1 U402 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n348) );
  XNOR2_X1 U403 ( .A(G1GAT), .B(KEYINPUT79), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n363) );
  XOR2_X1 U405 ( .A(G8GAT), .B(KEYINPUT75), .Z(n403) );
  XOR2_X1 U406 ( .A(n403), .B(n349), .Z(n351) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U409 ( .A(n352), .B(G64GAT), .Z(n354) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U412 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U413 ( .A(G15GAT), .B(G127GAT), .Z(n441) );
  XOR2_X1 U414 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n358) );
  XNOR2_X1 U415 ( .A(KEYINPUT14), .B(KEYINPUT78), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n441), .B(n359), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  NOR2_X1 U419 ( .A1(n586), .A2(n558), .ZN(n364) );
  XOR2_X1 U420 ( .A(KEYINPUT45), .B(n364), .Z(n365) );
  NOR2_X1 U421 ( .A1(n382), .A2(n365), .ZN(n381) );
  XOR2_X1 U422 ( .A(n366), .B(KEYINPUT29), .Z(n368) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U425 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n370) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G8GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U428 ( .A(n372), .B(n371), .Z(n380) );
  XOR2_X1 U429 ( .A(G15GAT), .B(G50GAT), .Z(n374) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(G43GAT), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U432 ( .A(G22GAT), .B(G197GAT), .Z(n376) );
  XNOR2_X1 U433 ( .A(G113GAT), .B(G141GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n564) );
  NAND2_X1 U437 ( .A1(n381), .A2(n564), .ZN(n391) );
  XNOR2_X1 U438 ( .A(n382), .B(KEYINPUT41), .ZN(n567) );
  NOR2_X1 U439 ( .A1(n564), .A2(n567), .ZN(n384) );
  XNOR2_X1 U440 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(KEYINPUT109), .B(n558), .ZN(n543) );
  NOR2_X1 U443 ( .A1(n385), .A2(n543), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n386), .B(KEYINPUT111), .ZN(n387) );
  INV_X1 U445 ( .A(n562), .ZN(n547) );
  NOR2_X1 U446 ( .A1(n387), .A2(n547), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  NAND2_X1 U448 ( .A1(n391), .A2(n390), .ZN(n393) );
  XOR2_X1 U449 ( .A(G183GAT), .B(KEYINPUT19), .Z(n395) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT18), .B(KEYINPUT82), .Z(n397) );
  XNOR2_X1 U453 ( .A(G190GAT), .B(KEYINPUT83), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n447) );
  XNOR2_X1 U456 ( .A(n447), .B(n400), .ZN(n409) );
  XOR2_X1 U457 ( .A(G204GAT), .B(G176GAT), .Z(n402) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U460 ( .A(n404), .B(n403), .Z(n407) );
  XNOR2_X1 U461 ( .A(G36GAT), .B(n405), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n467) );
  XNOR2_X1 U464 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n410), .B(KEYINPUT119), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n432) );
  XOR2_X1 U467 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n414) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n431) );
  XNOR2_X1 U470 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n415), .B(KEYINPUT80), .ZN(n434) );
  XNOR2_X1 U472 ( .A(n434), .B(n416), .ZN(n429) );
  XOR2_X1 U473 ( .A(G85GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G134GAT), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U476 ( .A(G148GAT), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U477 ( .A(G127GAT), .B(G120GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n427) );
  XOR2_X1 U480 ( .A(G57GAT), .B(KEYINPUT5), .Z(n424) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT4), .B(n425), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n529) );
  NAND2_X1 U487 ( .A1(n432), .A2(n529), .ZN(n571) );
  XOR2_X1 U488 ( .A(KEYINPUT55), .B(n433), .Z(n450) );
  XOR2_X1 U489 ( .A(KEYINPUT81), .B(n434), .Z(n439) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n436) );
  XNOR2_X1 U491 ( .A(G99GAT), .B(G71GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n437), .B(KEYINPUT85), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n445) );
  XOR2_X1 U495 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n460) );
  NAND2_X1 U501 ( .A1(n450), .A2(n460), .ZN(n451) );
  INV_X1 U502 ( .A(n566), .ZN(n455) );
  NAND2_X1 U503 ( .A1(n455), .A2(n543), .ZN(n454) );
  XNOR2_X1 U504 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(G1350GAT) );
  NAND2_X1 U506 ( .A1(n455), .A2(n547), .ZN(n458) );
  XOR2_X1 U507 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n456) );
  NOR2_X1 U508 ( .A1(n564), .A2(n382), .ZN(n491) );
  NOR2_X1 U509 ( .A1(n547), .A2(n558), .ZN(n459) );
  XNOR2_X1 U510 ( .A(KEYINPUT16), .B(n459), .ZN(n476) );
  INV_X1 U511 ( .A(n460), .ZN(n536) );
  INV_X1 U512 ( .A(n467), .ZN(n519) );
  NOR2_X1 U513 ( .A1(n536), .A2(n519), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n470), .A2(n461), .ZN(n462) );
  XNOR2_X1 U515 ( .A(KEYINPUT92), .B(n462), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(KEYINPUT25), .ZN(n464) );
  NAND2_X1 U517 ( .A1(n464), .A2(n529), .ZN(n469) );
  XOR2_X1 U518 ( .A(KEYINPUT91), .B(KEYINPUT26), .Z(n466) );
  NAND2_X1 U519 ( .A1(n470), .A2(n536), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n466), .B(n465), .ZN(n572) );
  XOR2_X1 U521 ( .A(n467), .B(KEYINPUT27), .Z(n530) );
  NOR2_X1 U522 ( .A1(n572), .A2(n530), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n475) );
  XNOR2_X1 U524 ( .A(KEYINPUT86), .B(n536), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n471), .A2(n534), .ZN(n472) );
  NOR2_X1 U526 ( .A1(n472), .A2(n530), .ZN(n473) );
  NOR2_X1 U527 ( .A1(n529), .A2(n473), .ZN(n474) );
  NOR2_X1 U528 ( .A1(n475), .A2(n474), .ZN(n489) );
  AND2_X1 U529 ( .A1(n476), .A2(n489), .ZN(n507) );
  NAND2_X1 U530 ( .A1(n491), .A2(n507), .ZN(n485) );
  NOR2_X1 U531 ( .A1(n529), .A2(n485), .ZN(n478) );
  XNOR2_X1 U532 ( .A(KEYINPUT34), .B(KEYINPUT93), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n519), .A2(n485), .ZN(n481) );
  XNOR2_X1 U536 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  NOR2_X1 U539 ( .A1(n536), .A2(n485), .ZN(n484) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n534), .A2(n485), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT96), .B(n486), .Z(n487) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(n487), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(KEYINPUT97), .Z(n493) );
  INV_X1 U546 ( .A(n558), .ZN(n580) );
  NOR2_X1 U547 ( .A1(n586), .A2(n580), .ZN(n488) );
  NAND2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n490), .ZN(n517) );
  NAND2_X1 U550 ( .A1(n491), .A2(n517), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n502) );
  NOR2_X1 U552 ( .A1(n502), .A2(n529), .ZN(n496) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT98), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n502), .A2(n519), .ZN(n498) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT99), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  NOR2_X1 U559 ( .A1(n502), .A2(n536), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U562 ( .A(G43GAT), .B(n501), .Z(G1330GAT) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n504) );
  NOR2_X1 U564 ( .A1(n534), .A2(n502), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT102), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n509) );
  INV_X1 U569 ( .A(n564), .ZN(n573) );
  NOR2_X1 U570 ( .A1(n567), .A2(n573), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n516), .A2(n507), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n529), .A2(n512), .ZN(n508) );
  XOR2_X1 U573 ( .A(n509), .B(n508), .Z(G1332GAT) );
  NOR2_X1 U574 ( .A1(n519), .A2(n512), .ZN(n510) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n536), .A2(n512), .ZN(n511) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n534), .A2(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n529), .A2(n526), .ZN(n518) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n526), .ZN(n520) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n536), .A2(n526), .ZN(n522) );
  XNOR2_X1 U588 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n525) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(KEYINPUT108), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n534), .A2(n526), .ZN(n527) );
  XOR2_X1 U595 ( .A(n528), .B(n527), .Z(G1339GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT113), .B(n533), .ZN(n552) );
  NAND2_X1 U599 ( .A1(n552), .A2(n534), .ZN(n535) );
  NOR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n548), .A2(n573), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT114), .B(n537), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n541) );
  INV_X1 U605 ( .A(n567), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n548), .A2(n539), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n542), .Z(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n545) );
  NAND2_X1 U610 ( .A1(n548), .A2(n543), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  INV_X1 U616 ( .A(n572), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n564), .A2(n561), .ZN(n553) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n561), .A2(n567), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n561), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT118), .B(n559), .Z(n560) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n566), .ZN(n565) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n570), .ZN(G1349GAT) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U637 ( .A1(n573), .A2(n584), .ZN(n577) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U643 ( .A1(n584), .A2(n382), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n584), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n583) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n588) );
  INV_X1 U650 ( .A(n584), .ZN(n585) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(n588), .B(n587), .Z(G1355GAT) );
endmodule

