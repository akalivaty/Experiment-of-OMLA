//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT65), .B1(new_n190), .B2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n188), .A3(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(new_n191), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT11), .A2(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT66), .A2(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT11), .A2(G134), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT11), .A2(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n210), .B2(new_n214), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n204), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n214), .A3(new_n211), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n203), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n224));
  INV_X1    g038(.A(G113), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n226), .A2(new_n227), .B1(KEYINPUT2), .B2(G113), .ZN(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT2), .A2(G113), .ZN(new_n232));
  AND4_X1   g046(.A1(KEYINPUT68), .A2(new_n231), .A3(new_n232), .A4(new_n229), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n207), .A2(new_n236), .A3(new_n209), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n211), .B1(G134), .B2(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n220), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n193), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n199), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n222), .A2(new_n235), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n187), .B1(new_n249), .B2(KEYINPUT28), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n194), .A2(new_n193), .B1(new_n199), .B2(new_n201), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n219), .A2(new_n220), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n251), .A2(new_n252), .B1(new_n240), .B2(new_n247), .ZN(new_n253));
  INV_X1    g067(.A(new_n235), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT28), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n215), .A2(new_n216), .A3(new_n204), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT69), .B1(new_n219), .B2(new_n220), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n251), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n240), .A2(new_n247), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(KEYINPUT71), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n264));
  NOR2_X1   g078(.A1(G237), .A2(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G210), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G101), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n250), .A2(new_n256), .A3(new_n263), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n222), .A2(new_n271), .A3(new_n248), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n273));
  OAI21_X1  g087(.A(new_n235), .B1(new_n253), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n261), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n269), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT29), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT72), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n261), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n249), .A2(KEYINPUT73), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n262), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n250), .A2(new_n263), .A3(KEYINPUT29), .A4(new_n269), .ZN(new_n286));
  OAI211_X1 g100(.A(KEYINPUT74), .B(new_n280), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n270), .A2(new_n277), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n250), .A2(new_n263), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n235), .B1(new_n222), .B2(new_n248), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n249), .B2(KEYINPUT73), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n261), .A2(new_n282), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT28), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n291), .A2(new_n295), .A3(KEYINPUT29), .A4(new_n269), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT74), .B1(new_n296), .B2(new_n280), .ZN(new_n297));
  OAI21_X1  g111(.A(G472), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT75), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n250), .A2(new_n256), .A3(new_n263), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n261), .B(new_n269), .C1(new_n272), .C2(new_n274), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n259), .A2(KEYINPUT30), .A3(new_n260), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n252), .A2(new_n251), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n260), .ZN(new_n306));
  INV_X1    g120(.A(new_n273), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n254), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n309), .A2(KEYINPUT31), .A3(new_n261), .A4(new_n269), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n276), .A2(new_n300), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G472), .A2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT32), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n300), .A2(new_n276), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n303), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT32), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n312), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n321), .B(G472), .C1(new_n290), .C2(new_n297), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n299), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G217), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(G234), .B2(new_n280), .ZN(new_n325));
  INV_X1    g139(.A(G953), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(G221), .A3(G234), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT78), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G140), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT16), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n336));
  OR3_X1    g150(.A1(new_n335), .A2(new_n188), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n188), .B1(new_n335), .B2(new_n336), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n241), .A2(G119), .ZN(new_n340));
  INV_X1    g154(.A(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G128), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT24), .B(G110), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT23), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n340), .A2(KEYINPUT76), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n349), .A3(new_n342), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n350), .B2(G110), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n344), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n350), .B2(G110), .ZN(new_n354));
  XNOR2_X1  g168(.A(G125), .B(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n188), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n337), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n352), .A2(new_n357), .A3(KEYINPUT77), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT77), .B1(new_n352), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n330), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n352), .A2(new_n357), .ZN(new_n361));
  INV_X1    g175(.A(new_n330), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT25), .B1(new_n364), .B2(new_n280), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  AOI211_X1 g180(.A(new_n366), .B(G902), .C1(new_n360), .C2(new_n363), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n325), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n325), .A2(G902), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT9), .B(G234), .ZN(new_n373));
  OAI21_X1  g187(.A(G221), .B1(new_n373), .B2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G110), .B(G140), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n326), .A2(G227), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT3), .B1(new_n380), .B2(G107), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n382));
  INV_X1    g196(.A(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(G104), .ZN(new_n384));
  INV_X1    g198(.A(G101), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(G107), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n381), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n380), .A2(G107), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n383), .A2(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(G101), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n247), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(KEYINPUT80), .B(KEYINPUT1), .C1(new_n190), .C2(G146), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G128), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT80), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n192), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT81), .B(new_n192), .C1(new_n394), .C2(new_n395), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n243), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n392), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT12), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n219), .B2(new_n220), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n217), .A2(new_n221), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n406), .B(new_n403), .C1(new_n401), .C2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n391), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n192), .A2(KEYINPUT1), .A3(new_n241), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n396), .B2(new_n397), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n407), .B1(new_n414), .B2(new_n392), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n406), .B1(new_n415), .B2(new_n403), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n405), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n400), .A2(new_n391), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n381), .A2(new_n384), .A3(new_n386), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(G101), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT4), .A4(G101), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n251), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n247), .A2(new_n391), .A3(KEYINPUT10), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n421), .A2(new_n408), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n379), .B1(new_n417), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n379), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n414), .A2(new_n419), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n430), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n407), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n432), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n403), .B1(new_n401), .B2(new_n408), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT83), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n442), .A2(new_n409), .B1(new_n402), .B2(new_n404), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n435), .A2(new_n436), .A3(new_n407), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n378), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n437), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT84), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G469), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n379), .B1(new_n431), .B2(new_n437), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n417), .B2(new_n434), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(G469), .A3(G902), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n280), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n375), .B1(new_n448), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G116), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G119), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT5), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n225), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n341), .A2(G116), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(G119), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT5), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n461), .A2(KEYINPUT86), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT86), .B1(new_n461), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n231), .A2(new_n232), .A3(new_n229), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n228), .A2(KEYINPUT68), .A3(new_n229), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n467), .A2(new_n472), .A3(new_n391), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n230), .B1(new_n426), .B2(new_n427), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n457), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n235), .A2(new_n428), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n467), .A2(new_n472), .A3(new_n391), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n456), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(new_n457), .C1(new_n473), .C2(new_n474), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n203), .A2(G125), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n243), .A2(new_n246), .A3(new_n333), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G224), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n484), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n243), .A2(new_n246), .A3(KEYINPUT88), .A4(new_n333), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n482), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(KEYINPUT7), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n478), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT87), .B(KEYINPUT8), .Z(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n456), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n461), .A2(new_n464), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n472), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n500), .B2(new_n391), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n467), .A2(new_n472), .A3(new_n411), .ZN(new_n502));
  INV_X1    g316(.A(new_n494), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(new_n502), .B1(new_n484), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n489), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n489), .A2(new_n505), .A3(new_n507), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G214), .B1(G237), .B2(G902), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT85), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(G234), .A2(G237), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(G952), .A3(new_n326), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(G902), .A3(G953), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT21), .B(G898), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n380), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n355), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT19), .B1(new_n355), .B2(KEYINPUT90), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n188), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n265), .A2(G143), .A3(G214), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(G143), .B1(new_n265), .B2(G214), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G237), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n326), .A3(G214), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n190), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n211), .A3(new_n529), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n528), .A2(new_n537), .A3(new_n337), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n332), .A2(new_n334), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G146), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n356), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n356), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n535), .A2(new_n529), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n545), .B1(new_n546), .B2(new_n211), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n535), .A2(KEYINPUT18), .A3(G131), .A4(new_n529), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n542), .A2(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n525), .B1(new_n538), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n542), .A2(new_n544), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n532), .A2(new_n554), .A3(new_n536), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n545), .A2(KEYINPUT17), .A3(G131), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n338), .A3(new_n337), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n524), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G475), .A2(G902), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT20), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT20), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n373), .A2(new_n324), .A3(G953), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n190), .A2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n241), .A2(G143), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n236), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n458), .A2(G122), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n458), .A2(G122), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n383), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n570), .A2(new_n571), .A3(G107), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT91), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(new_n568), .C1(new_n576), .C2(new_n567), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n579), .B2(G134), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n574), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n236), .B1(new_n567), .B2(new_n568), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n569), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT14), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n571), .B1(new_n570), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n458), .A2(G122), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT14), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n588), .B2(KEYINPUT14), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(G107), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n593), .B2(G107), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n582), .B(new_n585), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n566), .B1(new_n581), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n585), .A2(new_n582), .ZN(new_n600));
  INV_X1    g414(.A(new_n597), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(new_n595), .ZN(new_n602));
  INV_X1    g416(.A(new_n566), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n602), .A2(new_n580), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n280), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G478), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(KEYINPUT15), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(KEYINPUT15), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n603), .B1(new_n602), .B2(new_n580), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n581), .A2(new_n598), .A3(new_n566), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n558), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n524), .B1(new_n553), .B2(new_n557), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n280), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G475), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n565), .A2(new_n612), .A3(new_n617), .A4(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n515), .A2(new_n522), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n323), .A2(new_n372), .A3(new_n455), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n317), .A2(new_n280), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n626), .A2(G472), .B1(new_n317), .B2(new_n312), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n455), .A2(new_n372), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n509), .A2(KEYINPUT95), .A3(new_n510), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n489), .A2(new_n505), .A3(new_n630), .A4(new_n507), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n514), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT33), .B1(new_n599), .B2(new_n604), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n613), .A2(new_n614), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(G478), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n606), .A2(new_n280), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n615), .B2(new_n606), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n565), .A2(new_n621), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n633), .A2(new_n642), .A3(new_n522), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n628), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(new_n641), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n612), .A2(new_n617), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n633), .A2(new_n522), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n628), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n383), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  OR2_X1    g468(.A1(new_n358), .A2(new_n359), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n330), .A2(KEYINPUT36), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n370), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n368), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n455), .A2(new_n623), .A3(new_n627), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT97), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  XOR2_X1   g478(.A(KEYINPUT98), .B(G900), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n520), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n517), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n631), .A2(new_n514), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n489), .A2(new_n505), .A3(new_n507), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n507), .B1(new_n489), .B2(new_n505), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n670), .B1(new_n673), .B2(KEYINPUT95), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n669), .A2(new_n674), .A3(new_n660), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n322), .A2(new_n320), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT74), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n287), .A3(new_n279), .A4(new_n289), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n321), .B1(new_n680), .B2(G472), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n675), .B(new_n455), .C1(new_n676), .C2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n673), .A2(KEYINPUT38), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n511), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n565), .A2(new_n621), .B1(new_n612), .B2(new_n617), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n368), .A3(new_n514), .A4(new_n659), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n684), .B(new_n686), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n283), .A2(new_n284), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(new_n276), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n693), .B(new_n276), .C1(new_n293), .C2(new_n294), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n301), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n280), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT100), .B1(new_n320), .B2(new_n699), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n320), .A2(KEYINPUT100), .A3(new_n699), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n692), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT102), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n667), .B(KEYINPUT39), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n455), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n692), .B(new_n708), .C1(new_n700), .C2(new_n701), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n703), .A2(new_n706), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  AND4_X1   g525(.A1(new_n641), .A2(new_n637), .A3(new_n639), .A4(new_n667), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n368), .A2(new_n659), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n714), .A3(new_n633), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n455), .B(new_n715), .C1(new_n676), .C2(new_n681), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  OAI21_X1  g531(.A(G469), .B1(new_n450), .B2(G902), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n442), .A2(new_n409), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n433), .B1(new_n719), .B2(new_n405), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n452), .B(new_n280), .C1(new_n720), .C2(new_n449), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n374), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT103), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n323), .A2(new_n372), .A3(new_n643), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n323), .A2(new_n372), .A3(new_n650), .A4(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  AND3_X1   g542(.A1(new_n718), .A2(new_n374), .A3(new_n721), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n674), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n722), .B2(new_n633), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n714), .A2(new_n522), .A3(new_n622), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n323), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  XOR2_X1   g550(.A(KEYINPUT105), .B(G472), .Z(new_n737));
  NAND2_X1  g551(.A1(new_n626), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n269), .B1(new_n291), .B2(new_n295), .ZN(new_n739));
  INV_X1    g553(.A(new_n316), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n312), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n372), .ZN(new_n743));
  INV_X1    g557(.A(new_n522), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n641), .A2(new_n648), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n633), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(new_n723), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  AND4_X1   g562(.A1(new_n660), .A2(new_n738), .A3(new_n712), .A4(new_n741), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT104), .B1(new_n729), .B2(new_n674), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n722), .A2(new_n633), .A3(new_n731), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  INV_X1    g567(.A(new_n372), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n322), .A2(new_n320), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(new_n299), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n375), .A2(new_n513), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n673), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n453), .B(KEYINPUT106), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n451), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n445), .A2(KEYINPUT107), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n432), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n764), .A3(G469), .A4(new_n446), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n758), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n756), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n372), .B(new_n766), .C1(new_n676), .C2(new_n681), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n713), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  INV_X1    g586(.A(new_n669), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n236), .ZN(G36));
  NAND2_X1  g589(.A1(new_n640), .A2(new_n647), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n627), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n660), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT109), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n673), .A2(new_n514), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n780), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n439), .B1(new_n432), .B2(new_n438), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n445), .A2(KEYINPUT84), .A3(new_n446), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT45), .A4(new_n446), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(G469), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n759), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n760), .A2(new_n796), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n451), .B1(new_n794), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(KEYINPUT108), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT108), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n374), .B(new_n704), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n788), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT110), .B(G137), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G39));
  NAND2_X1  g620(.A1(new_n794), .A2(new_n798), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n721), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n808), .A2(new_n809), .B1(new_n796), .B2(new_n795), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n375), .B1(new_n810), .B2(new_n801), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT47), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n374), .B1(new_n800), .B2(new_n802), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n323), .A2(new_n372), .A3(new_n713), .A4(new_n783), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NAND2_X1  g633(.A1(new_n372), .A2(new_n757), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT111), .Z(new_n821));
  NAND2_X1  g635(.A1(new_n684), .A2(new_n686), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n718), .A2(new_n721), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT49), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n821), .A2(new_n823), .A3(new_n776), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n701), .A2(new_n700), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(KEYINPUT49), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n326), .A2(G952), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n743), .A2(new_n778), .A3(new_n518), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(new_n832), .B2(new_n733), .ZN(new_n833));
  INV_X1    g647(.A(new_n783), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n729), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n827), .A2(new_n372), .A3(new_n518), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n833), .B1(new_n642), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n518), .A3(new_n778), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT115), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(new_n756), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(KEYINPUT117), .A3(KEYINPUT48), .ZN(new_n842));
  XOR2_X1   g656(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n843));
  AOI211_X1 g657(.A(new_n838), .B(new_n842), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n742), .A2(new_n660), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT116), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n822), .A2(new_n729), .A3(new_n513), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n831), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n850), .A2(KEYINPUT50), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(KEYINPUT50), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n640), .A2(new_n641), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n851), .A2(new_n852), .B1(new_n837), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n824), .A2(new_n374), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n834), .B(new_n832), .C1(new_n816), .C2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n857), .B1(new_n856), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n844), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n624), .A2(new_n735), .A3(new_n747), .A4(new_n661), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n642), .A2(new_n649), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n522), .A3(new_n515), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n372), .A3(new_n455), .A4(new_n627), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n724), .A2(new_n727), .A3(new_n868), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n714), .A2(new_n783), .A3(new_n622), .A4(new_n668), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n870), .B(new_n455), .C1(new_n676), .C2(new_n681), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n749), .A2(new_n766), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n871), .B(new_n872), .C1(new_n769), .C2(new_n773), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n865), .A2(new_n771), .A3(new_n869), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n667), .A2(new_n374), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n633), .A2(new_n660), .A3(new_n745), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n761), .A2(new_n765), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n877), .B(new_n878), .C1(new_n701), .C2(new_n700), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n682), .A2(new_n716), .A3(new_n879), .A4(new_n752), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n323), .B(new_n455), .C1(new_n675), .C2(new_n715), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(KEYINPUT52), .A3(new_n752), .A4(new_n879), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n864), .B1(new_n875), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n884), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n624), .A2(new_n735), .A3(new_n747), .A4(new_n661), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n724), .A2(new_n727), .A3(new_n868), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n873), .B1(new_n770), .B2(new_n767), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n887), .A2(new_n890), .A3(new_n891), .A4(KEYINPUT53), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(KEYINPUT112), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n864), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(KEYINPUT54), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n886), .A2(new_n898), .A3(new_n892), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n894), .A2(KEYINPUT114), .A3(new_n864), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n863), .B(new_n897), .C1(new_n901), .C2(KEYINPUT54), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n897), .A2(new_n863), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n862), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n829), .B1(new_n904), .B2(new_n905), .ZN(G75));
  NAND3_X1  g720(.A1(new_n901), .A2(G210), .A3(G902), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n479), .A2(new_n481), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n488), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n907), .B2(new_n908), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n326), .A2(G952), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G51));
  XOR2_X1   g730(.A(new_n759), .B(KEYINPUT57), .Z(new_n917));
  AND3_X1   g731(.A1(new_n899), .A2(KEYINPUT54), .A3(new_n900), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT54), .B1(new_n899), .B2(new_n900), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n720), .B2(new_n449), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n794), .B(KEYINPUT119), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n901), .A2(G902), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n915), .B1(new_n921), .B2(new_n923), .ZN(G54));
  NAND2_X1  g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT120), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n901), .A2(G902), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n559), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n915), .ZN(G60));
  AND2_X1   g745(.A1(new_n634), .A2(new_n636), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n638), .B(KEYINPUT59), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n918), .B2(new_n919), .ZN(new_n935));
  INV_X1    g749(.A(new_n915), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n933), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n902), .A2(new_n903), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n939), .B2(new_n932), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  NAND3_X1  g756(.A1(new_n899), .A2(new_n900), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n364), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n657), .A2(new_n658), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n899), .A2(new_n946), .A3(new_n900), .A4(new_n942), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n936), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT61), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT61), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n521), .B2(new_n485), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n890), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n909), .B1(G898), .B2(new_n326), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  INV_X1    g771(.A(new_n804), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n818), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n866), .A2(new_n783), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n756), .A2(new_n455), .A3(new_n704), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n883), .A2(new_n752), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n710), .A2(KEYINPUT62), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT62), .B1(new_n710), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n326), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n304), .B1(new_n253), .B2(new_n273), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT123), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n526), .A2(new_n527), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n804), .B1(new_n816), .B2(new_n817), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n756), .A2(new_n746), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT125), .B1(new_n803), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n811), .A2(new_n977), .A3(new_n704), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n774), .B(new_n962), .C1(new_n770), .C2(new_n767), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n974), .A2(new_n326), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n971), .B1(G900), .B2(G953), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n972), .A2(new_n973), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n326), .B1(G227), .B2(G900), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n972), .A2(KEYINPUT126), .A3(new_n984), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n987), .ZN(new_n991));
  AOI22_X1  g805(.A1(new_n967), .A2(new_n971), .B1(new_n982), .B2(new_n983), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT126), .B1(new_n992), .B2(new_n973), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(new_n275), .A2(new_n269), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n959), .A2(new_n966), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n890), .ZN(new_n998));
  XOR2_X1   g812(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n996), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n974), .A2(new_n890), .A3(new_n980), .A4(new_n981), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n269), .B(new_n275), .C1(new_n1003), .C2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n893), .A2(new_n896), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n275), .A2(new_n276), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n301), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n1001), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n936), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1002), .A2(new_n1004), .A3(new_n1009), .ZN(G57));
endmodule


