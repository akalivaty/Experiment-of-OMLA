

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n766), .A2(n515), .ZN(n796) );
  XOR2_X2 U552 ( .A(KEYINPUT1), .B(n516), .Z(n590) );
  XNOR2_X1 U553 ( .A(n762), .B(KEYINPUT99), .ZN(n766) );
  XOR2_X1 U554 ( .A(KEYINPUT66), .B(n541), .Z(n514) );
  OR2_X1 U555 ( .A1(n765), .A2(n764), .ZN(n515) );
  XNOR2_X1 U556 ( .A(n687), .B(KEYINPUT90), .ZN(n697) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n705) );
  XNOR2_X1 U558 ( .A(KEYINPUT95), .B(KEYINPUT29), .ZN(n709) );
  XNOR2_X1 U559 ( .A(n710), .B(n709), .ZN(n715) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n783) );
  NOR2_X2 U561 ( .A1(n629), .A2(n520), .ZN(n643) );
  NOR2_X1 U562 ( .A1(G543), .A2(G651), .ZN(n640) );
  NOR2_X1 U563 ( .A1(n629), .A2(G651), .ZN(n646) );
  INV_X1 U564 ( .A(G651), .ZN(n520) );
  NOR2_X1 U565 ( .A1(G543), .A2(n520), .ZN(n516) );
  NAND2_X1 U566 ( .A1(G63), .A2(n590), .ZN(n518) );
  XOR2_X1 U567 ( .A(KEYINPUT0), .B(G543), .Z(n629) );
  NAND2_X1 U568 ( .A1(G51), .A2(n646), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U570 ( .A(KEYINPUT6), .B(n519), .Z(n528) );
  NAND2_X1 U571 ( .A1(G76), .A2(n643), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n522) );
  NAND2_X1 U573 ( .A1(G89), .A2(n640), .ZN(n521) );
  XNOR2_X1 U574 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U576 ( .A(n525), .B(KEYINPUT5), .ZN(n526) );
  XNOR2_X1 U577 ( .A(KEYINPUT76), .B(n526), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U579 ( .A(KEYINPUT7), .B(n529), .ZN(G168) );
  XOR2_X1 U580 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U581 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n534), .A2(G2104), .ZN(n530) );
  XNOR2_X2 U583 ( .A(n530), .B(KEYINPUT65), .ZN(n983) );
  NAND2_X1 U584 ( .A1(G102), .A2(n983), .ZN(n533) );
  NOR2_X2 U585 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  XOR2_X2 U586 ( .A(KEYINPUT17), .B(n531), .Z(n984) );
  NAND2_X1 U587 ( .A1(G138), .A2(n984), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n538) );
  AND2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n979) );
  NAND2_X1 U590 ( .A1(G114), .A2(n979), .ZN(n536) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n534), .ZN(n980) );
  NAND2_X1 U592 ( .A1(G126), .A2(n980), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U594 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U595 ( .A1(G137), .A2(n984), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G113), .A2(n979), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n980), .A2(G125), .ZN(n542) );
  AND2_X1 U599 ( .A1(n514), .A2(n542), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G101), .A2(n983), .ZN(n543) );
  XOR2_X1 U601 ( .A(KEYINPUT23), .B(n543), .Z(n544) );
  AND2_X2 U602 ( .A1(n545), .A2(n544), .ZN(G160) );
  NAND2_X1 U603 ( .A1(G72), .A2(n643), .ZN(n547) );
  NAND2_X1 U604 ( .A1(G85), .A2(n640), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G60), .A2(n590), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G47), .A2(n646), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U609 ( .A1(n551), .A2(n550), .ZN(G290) );
  NAND2_X1 U610 ( .A1(G64), .A2(n590), .ZN(n553) );
  NAND2_X1 U611 ( .A1(G52), .A2(n646), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n643), .A2(G77), .ZN(n554) );
  XOR2_X1 U614 ( .A(KEYINPUT67), .B(n554), .Z(n556) );
  NAND2_X1 U615 ( .A1(n640), .A2(G90), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U618 ( .A1(n559), .A2(n558), .ZN(G171) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U620 ( .A1(n983), .A2(G99), .ZN(n560) );
  XOR2_X1 U621 ( .A(KEYINPUT79), .B(n560), .Z(n562) );
  NAND2_X1 U622 ( .A1(n979), .A2(G111), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U624 ( .A(KEYINPUT80), .B(n563), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n980), .A2(G123), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT18), .B(n564), .Z(n565) );
  NOR2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n984), .A2(G135), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n1005) );
  XNOR2_X1 U630 ( .A(G2096), .B(n1005), .ZN(n569) );
  OR2_X1 U631 ( .A1(G2100), .A2(n569), .ZN(G156) );
  NAND2_X1 U632 ( .A1(G56), .A2(n590), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT14), .ZN(n571) );
  XNOR2_X1 U634 ( .A(KEYINPUT69), .B(n571), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n640), .A2(G81), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT12), .B(n572), .Z(n576) );
  INV_X1 U637 ( .A(KEYINPUT70), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n643), .A2(G68), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(n577), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n646), .A2(G43), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n680) );
  INV_X1 U645 ( .A(G860), .ZN(n617) );
  OR2_X1 U646 ( .A1(n680), .A2(n617), .ZN(G153) );
  NAND2_X1 U647 ( .A1(G65), .A2(n590), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G53), .A2(n646), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G78), .A2(n643), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G91), .A2(n640), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n703) );
  INV_X1 U654 ( .A(n703), .ZN(G299) );
  INV_X1 U655 ( .A(G57), .ZN(G237) );
  INV_X1 U656 ( .A(G82), .ZN(G220) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n588), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U659 ( .A(G223), .ZN(n814) );
  NAND2_X1 U660 ( .A1(n814), .A2(G567), .ZN(n589) );
  XOR2_X1 U661 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  INV_X1 U662 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G54), .A2(n646), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G66), .A2(n590), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G79), .A2(n643), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G92), .A2(n640), .ZN(n593) );
  XNOR2_X1 U669 ( .A(KEYINPUT71), .B(n593), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n598), .B(KEYINPUT15), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n600), .B(n599), .ZN(n1009) );
  INV_X1 U674 ( .A(G868), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n1009), .A2(n604), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT74), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(G284) );
  NOR2_X1 U679 ( .A1(G286), .A2(n604), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n617), .A2(G559), .ZN(n607) );
  INV_X1 U683 ( .A(n1009), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n607), .A2(n614), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n680), .ZN(n609) );
  XOR2_X1 U687 ( .A(KEYINPUT77), .B(n609), .Z(n612) );
  NAND2_X1 U688 ( .A1(G868), .A2(n614), .ZN(n610) );
  NOR2_X1 U689 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U691 ( .A(KEYINPUT78), .B(n613), .ZN(G282) );
  XNOR2_X1 U692 ( .A(n680), .B(KEYINPUT81), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n614), .A2(G559), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n616), .B(n615), .ZN(n657) );
  NAND2_X1 U695 ( .A1(n617), .A2(n657), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G67), .A2(n590), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G55), .A2(n646), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U699 ( .A(KEYINPUT82), .B(n620), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G80), .A2(n643), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G93), .A2(n640), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n659) );
  XOR2_X1 U704 ( .A(n625), .B(n659), .Z(G145) );
  NAND2_X1 U705 ( .A1(G49), .A2(n646), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n590), .A2(n628), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G87), .A2(n629), .ZN(n630) );
  XOR2_X1 U710 ( .A(KEYINPUT83), .B(n630), .Z(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U712 ( .A1(G61), .A2(n590), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G86), .A2(n640), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n643), .A2(G73), .ZN(n635) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n635), .Z(n636) );
  NOR2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n646), .A2(G48), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G88), .A2(n640), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT86), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n590), .A2(G62), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n642), .B(KEYINPUT84), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G75), .A2(n643), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G50), .A2(n646), .ZN(n647) );
  XNOR2_X1 U727 ( .A(KEYINPUT85), .B(n647), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(G303) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(G288), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n659), .B(G305), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n652), .B(G303), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n703), .B(n653), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n1008) );
  XNOR2_X1 U736 ( .A(n657), .B(n1008), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n658), .A2(G868), .ZN(n661) );
  OR2_X1 U738 ( .A1(G868), .A2(n659), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U746 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NOR2_X1 U747 ( .A1(G219), .A2(G220), .ZN(n666) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U749 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G96), .A2(n668), .ZN(n819) );
  NAND2_X1 U751 ( .A1(G2106), .A2(n819), .ZN(n669) );
  XOR2_X1 U752 ( .A(KEYINPUT87), .B(n669), .Z(n673) );
  NAND2_X1 U753 ( .A1(G69), .A2(G120), .ZN(n670) );
  NOR2_X1 U754 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U755 ( .A1(G108), .A2(n671), .ZN(n820) );
  NAND2_X1 U756 ( .A1(G567), .A2(n820), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n1014) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U759 ( .A1(n1014), .A2(n674), .ZN(n818) );
  NAND2_X1 U760 ( .A1(n818), .A2(G36), .ZN(G176) );
  AND2_X1 U761 ( .A1(n783), .A2(G40), .ZN(n678) );
  AND2_X1 U762 ( .A1(n678), .A2(G1996), .ZN(n675) );
  AND2_X1 U763 ( .A1(n675), .A2(G160), .ZN(n677) );
  XOR2_X1 U764 ( .A(KEYINPUT26), .B(KEYINPUT92), .Z(n676) );
  XNOR2_X1 U765 ( .A(n677), .B(n676), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G160), .A2(n678), .ZN(n687) );
  AND2_X1 U767 ( .A1(n687), .A2(G1341), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n682) );
  AND2_X1 U769 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U770 ( .A(KEYINPUT64), .B(n684), .Z(n692) );
  NOR2_X1 U771 ( .A1(n692), .A2(n1009), .ZN(n685) );
  XNOR2_X1 U772 ( .A(n685), .B(KEYINPUT93), .ZN(n691) );
  INV_X1 U773 ( .A(n697), .ZN(n711) );
  NAND2_X1 U774 ( .A1(G2067), .A2(n711), .ZN(n686) );
  XNOR2_X1 U775 ( .A(n686), .B(KEYINPUT94), .ZN(n689) );
  BUF_X1 U776 ( .A(n687), .Z(n725) );
  NAND2_X1 U777 ( .A1(G1348), .A2(n725), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U780 ( .A1(n692), .A2(n1009), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n702) );
  NAND2_X1 U782 ( .A1(G2072), .A2(n711), .ZN(n696) );
  INV_X1 U783 ( .A(KEYINPUT27), .ZN(n695) );
  XNOR2_X1 U784 ( .A(n696), .B(n695), .ZN(n699) );
  NAND2_X1 U785 ( .A1(G1956), .A2(n697), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U787 ( .A(n700), .B(KEYINPUT91), .ZN(n704) );
  NAND2_X1 U788 ( .A1(n703), .A2(n704), .ZN(n701) );
  NAND2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n708) );
  NOR2_X1 U790 ( .A1(n704), .A2(n703), .ZN(n706) );
  XNOR2_X1 U791 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U792 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U793 ( .A(G1961), .B(KEYINPUT89), .ZN(n909) );
  NAND2_X1 U794 ( .A1(n725), .A2(n909), .ZN(n713) );
  XNOR2_X1 U795 ( .A(G2078), .B(KEYINPUT25), .ZN(n868) );
  NAND2_X1 U796 ( .A1(n711), .A2(n868), .ZN(n712) );
  NAND2_X1 U797 ( .A1(n713), .A2(n712), .ZN(n719) );
  NAND2_X1 U798 ( .A1(G171), .A2(n719), .ZN(n714) );
  NAND2_X1 U799 ( .A1(n715), .A2(n714), .ZN(n724) );
  NAND2_X1 U800 ( .A1(G8), .A2(n725), .ZN(n765) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n765), .ZN(n736) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n725), .ZN(n733) );
  NOR2_X1 U803 ( .A1(n736), .A2(n733), .ZN(n716) );
  NAND2_X1 U804 ( .A1(G8), .A2(n716), .ZN(n717) );
  XNOR2_X1 U805 ( .A(KEYINPUT30), .B(n717), .ZN(n718) );
  NOR2_X1 U806 ( .A1(G168), .A2(n718), .ZN(n721) );
  NOR2_X1 U807 ( .A1(G171), .A2(n719), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U809 ( .A(KEYINPUT31), .B(n722), .Z(n723) );
  NAND2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n734) );
  NAND2_X1 U811 ( .A1(n734), .A2(G286), .ZN(n730) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n765), .ZN(n727) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n725), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n728), .A2(G303), .ZN(n729) );
  NAND2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U817 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U818 ( .A(n732), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U819 ( .A1(G8), .A2(n733), .ZN(n738) );
  INV_X1 U820 ( .A(n734), .ZN(n735) );
  NOR2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U822 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U823 ( .A1(n740), .A2(n739), .ZN(n758) );
  NOR2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n883) );
  INV_X1 U825 ( .A(n883), .ZN(n743) );
  NOR2_X1 U826 ( .A1(G1971), .A2(G303), .ZN(n882) );
  XOR2_X1 U827 ( .A(n882), .B(KEYINPUT96), .Z(n741) );
  INV_X1 U828 ( .A(KEYINPUT33), .ZN(n747) );
  AND2_X1 U829 ( .A1(n741), .A2(n747), .ZN(n742) );
  AND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n758), .A2(n744), .ZN(n749) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n884) );
  INV_X1 U833 ( .A(n765), .ZN(n745) );
  NAND2_X1 U834 ( .A1(n884), .A2(n745), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U837 ( .A(n750), .B(KEYINPUT97), .ZN(n754) );
  XNOR2_X1 U838 ( .A(G1981), .B(G305), .ZN(n900) );
  NAND2_X1 U839 ( .A1(n883), .A2(KEYINPUT33), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n765), .A2(n751), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n900), .A2(n752), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n761) );
  NOR2_X1 U843 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U844 ( .A1(G8), .A2(n755), .ZN(n756) );
  XNOR2_X1 U845 ( .A(KEYINPUT98), .B(n756), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n759), .A2(n765), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U850 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NAND2_X1 U851 ( .A1(G95), .A2(n983), .ZN(n768) );
  NAND2_X1 U852 ( .A1(G131), .A2(n984), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U854 ( .A1(G107), .A2(n979), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G119), .A2(n980), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n996) );
  INV_X1 U858 ( .A(G1991), .ZN(n862) );
  NOR2_X1 U859 ( .A1(n996), .A2(n862), .ZN(n781) );
  NAND2_X1 U860 ( .A1(G117), .A2(n979), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G129), .A2(n980), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n983), .A2(G105), .ZN(n775) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(n775), .Z(n776) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n984), .A2(G141), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n1000) );
  AND2_X1 U868 ( .A1(n1000), .A2(G1996), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n833) );
  NAND2_X1 U870 ( .A1(G160), .A2(G40), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n809) );
  INV_X1 U872 ( .A(n809), .ZN(n784) );
  NOR2_X1 U873 ( .A1(n833), .A2(n784), .ZN(n802) );
  XOR2_X1 U874 ( .A(KEYINPUT88), .B(n802), .Z(n794) );
  NAND2_X1 U875 ( .A1(G104), .A2(n983), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G140), .A2(n984), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n787), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G116), .A2(n979), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G128), .A2(n980), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT35), .B(n790), .Z(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U884 ( .A(KEYINPUT36), .B(n793), .ZN(n994) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n807) );
  NOR2_X1 U886 ( .A1(n994), .A2(n807), .ZN(n835) );
  NAND2_X1 U887 ( .A1(n809), .A2(n835), .ZN(n805) );
  NAND2_X1 U888 ( .A1(n794), .A2(n805), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n798) );
  XNOR2_X1 U890 ( .A(G1986), .B(G290), .ZN(n887) );
  NAND2_X1 U891 ( .A1(n887), .A2(n809), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n812) );
  NOR2_X1 U893 ( .A1(G1996), .A2(n1000), .ZN(n848) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n800) );
  AND2_X1 U895 ( .A1(n862), .A2(n996), .ZN(n799) );
  XNOR2_X1 U896 ( .A(KEYINPUT100), .B(n799), .ZN(n831) );
  NOR2_X1 U897 ( .A1(n800), .A2(n831), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n848), .A2(n803), .ZN(n804) );
  XNOR2_X1 U900 ( .A(n804), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n994), .A2(n807), .ZN(n829) );
  NAND2_X1 U903 ( .A1(n808), .A2(n829), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U906 ( .A(KEYINPUT40), .B(n813), .ZN(G329) );
  NAND2_X1 U907 ( .A1(n814), .A2(G2106), .ZN(n815) );
  XNOR2_X1 U908 ( .A(n815), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U910 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(G188) );
  NOR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(G325) );
  XNOR2_X1 U914 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  NAND2_X1 U916 ( .A1(G100), .A2(n983), .ZN(n822) );
  NAND2_X1 U917 ( .A1(G112), .A2(n979), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n823), .B(KEYINPUT109), .ZN(n825) );
  NAND2_X1 U920 ( .A1(G136), .A2(n984), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n980), .A2(G124), .ZN(n826) );
  XOR2_X1 U923 ( .A(KEYINPUT44), .B(n826), .Z(n827) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G162) );
  NAND2_X1 U925 ( .A1(n829), .A2(n1005), .ZN(n856) );
  XOR2_X1 U926 ( .A(G160), .B(G2084), .Z(n830) );
  NOR2_X1 U927 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n854) );
  NAND2_X1 U930 ( .A1(G103), .A2(n983), .ZN(n837) );
  NAND2_X1 U931 ( .A1(G139), .A2(n984), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n843) );
  NAND2_X1 U933 ( .A1(n980), .A2(G127), .ZN(n838) );
  XOR2_X1 U934 ( .A(KEYINPUT111), .B(n838), .Z(n840) );
  NAND2_X1 U935 ( .A1(n979), .A2(G115), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT47), .B(n841), .Z(n842) );
  NOR2_X1 U938 ( .A1(n843), .A2(n842), .ZN(n998) );
  XOR2_X1 U939 ( .A(G2072), .B(n998), .Z(n845) );
  XOR2_X1 U940 ( .A(G164), .B(G2078), .Z(n844) );
  NOR2_X1 U941 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U942 ( .A(KEYINPUT50), .B(n846), .Z(n852) );
  XOR2_X1 U943 ( .A(G2090), .B(G162), .Z(n847) );
  NOR2_X1 U944 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U945 ( .A(KEYINPUT116), .B(n849), .Z(n850) );
  XOR2_X1 U946 ( .A(KEYINPUT51), .B(n850), .Z(n851) );
  NOR2_X1 U947 ( .A1(n852), .A2(n851), .ZN(n853) );
  NAND2_X1 U948 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U949 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U950 ( .A(KEYINPUT52), .B(n857), .ZN(n858) );
  INV_X1 U951 ( .A(KEYINPUT55), .ZN(n878) );
  NAND2_X1 U952 ( .A1(n858), .A2(n878), .ZN(n859) );
  NAND2_X1 U953 ( .A1(n859), .A2(G29), .ZN(n943) );
  XNOR2_X1 U954 ( .A(G2090), .B(G35), .ZN(n873) );
  XNOR2_X1 U955 ( .A(G1996), .B(G32), .ZN(n861) );
  XNOR2_X1 U956 ( .A(G33), .B(G2072), .ZN(n860) );
  NOR2_X1 U957 ( .A1(n861), .A2(n860), .ZN(n867) );
  XNOR2_X1 U958 ( .A(G25), .B(n862), .ZN(n863) );
  NAND2_X1 U959 ( .A1(n863), .A2(G28), .ZN(n865) );
  XNOR2_X1 U960 ( .A(G26), .B(G2067), .ZN(n864) );
  NOR2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n866) );
  NAND2_X1 U962 ( .A1(n867), .A2(n866), .ZN(n870) );
  XOR2_X1 U963 ( .A(G27), .B(n868), .Z(n869) );
  NOR2_X1 U964 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U965 ( .A(KEYINPUT53), .B(n871), .ZN(n872) );
  NOR2_X1 U966 ( .A1(n873), .A2(n872), .ZN(n876) );
  XOR2_X1 U967 ( .A(G2084), .B(G34), .Z(n874) );
  XNOR2_X1 U968 ( .A(KEYINPUT54), .B(n874), .ZN(n875) );
  NAND2_X1 U969 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U970 ( .A(n878), .B(n877), .ZN(n880) );
  INV_X1 U971 ( .A(G29), .ZN(n879) );
  NAND2_X1 U972 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U973 ( .A1(G11), .A2(n881), .ZN(n941) );
  XNOR2_X1 U974 ( .A(G16), .B(KEYINPUT56), .ZN(n908) );
  XOR2_X1 U975 ( .A(G1348), .B(n1009), .Z(n893) );
  NOR2_X1 U976 ( .A1(n883), .A2(n882), .ZN(n885) );
  NAND2_X1 U977 ( .A1(n885), .A2(n884), .ZN(n891) );
  XNOR2_X1 U978 ( .A(G1956), .B(G299), .ZN(n886) );
  NOR2_X1 U979 ( .A1(n887), .A2(n886), .ZN(n889) );
  NAND2_X1 U980 ( .A1(G1971), .A2(G303), .ZN(n888) );
  NAND2_X1 U981 ( .A1(n889), .A2(n888), .ZN(n890) );
  NOR2_X1 U982 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U983 ( .A1(n893), .A2(n892), .ZN(n896) );
  XNOR2_X1 U984 ( .A(G1341), .B(n680), .ZN(n894) );
  XNOR2_X1 U985 ( .A(KEYINPUT120), .B(n894), .ZN(n895) );
  NOR2_X1 U986 ( .A1(n896), .A2(n895), .ZN(n906) );
  XNOR2_X1 U987 ( .A(G171), .B(G1961), .ZN(n897) );
  XNOR2_X1 U988 ( .A(n897), .B(KEYINPUT119), .ZN(n904) );
  XOR2_X1 U989 ( .A(KEYINPUT57), .B(KEYINPUT118), .Z(n902) );
  XNOR2_X1 U990 ( .A(G1966), .B(G168), .ZN(n898) );
  XNOR2_X1 U991 ( .A(n898), .B(KEYINPUT117), .ZN(n899) );
  NOR2_X1 U992 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U993 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U994 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U995 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U996 ( .A1(n908), .A2(n907), .ZN(n939) );
  INV_X1 U997 ( .A(G16), .ZN(n937) );
  XOR2_X1 U998 ( .A(G1966), .B(G21), .Z(n911) );
  XNOR2_X1 U999 ( .A(n909), .B(G5), .ZN(n910) );
  NAND2_X1 U1000 ( .A1(n911), .A2(n910), .ZN(n925) );
  XNOR2_X1 U1001 ( .A(KEYINPUT121), .B(G1956), .ZN(n912) );
  XNOR2_X1 U1002 ( .A(n912), .B(G20), .ZN(n916) );
  XOR2_X1 U1003 ( .A(G4), .B(KEYINPUT123), .Z(n914) );
  XNOR2_X1 U1004 ( .A(G1348), .B(KEYINPUT59), .ZN(n913) );
  XNOR2_X1 U1005 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1006 ( .A1(n916), .A2(n915), .ZN(n921) );
  XNOR2_X1 U1007 ( .A(G1981), .B(G6), .ZN(n918) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G19), .ZN(n917) );
  NOR2_X1 U1009 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1010 ( .A(n919), .B(KEYINPUT122), .Z(n920) );
  NOR2_X1 U1011 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1012 ( .A(KEYINPUT60), .B(n922), .Z(n923) );
  XNOR2_X1 U1013 ( .A(n923), .B(KEYINPUT124), .ZN(n924) );
  NOR2_X1 U1014 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1015 ( .A(KEYINPUT125), .B(n926), .ZN(n934) );
  XOR2_X1 U1016 ( .A(G1986), .B(G24), .Z(n930) );
  XNOR2_X1 U1017 ( .A(G1971), .B(G22), .ZN(n928) );
  XNOR2_X1 U1018 ( .A(G23), .B(G1976), .ZN(n927) );
  NOR2_X1 U1019 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1020 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1021 ( .A(KEYINPUT126), .B(n931), .ZN(n932) );
  XNOR2_X1 U1022 ( .A(KEYINPUT58), .B(n932), .ZN(n933) );
  NOR2_X1 U1023 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1024 ( .A(KEYINPUT61), .B(n935), .ZN(n936) );
  NAND2_X1 U1025 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1026 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1027 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1028 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1029 ( .A(KEYINPUT62), .B(n944), .Z(G311) );
  XNOR2_X1 U1030 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1031 ( .A(G120), .ZN(G236) );
  INV_X1 U1032 ( .A(G96), .ZN(G221) );
  INV_X1 U1033 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1034 ( .A(G2427), .B(G1348), .ZN(n954) );
  XOR2_X1 U1035 ( .A(G2451), .B(G2430), .Z(n946) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G2443), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n946), .B(n945), .ZN(n950) );
  XOR2_X1 U1038 ( .A(G2438), .B(KEYINPUT101), .Z(n948) );
  XNOR2_X1 U1039 ( .A(G2454), .B(G2435), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n948), .B(n947), .ZN(n949) );
  XOR2_X1 U1041 ( .A(n950), .B(n949), .Z(n952) );
  XNOR2_X1 U1042 ( .A(KEYINPUT102), .B(G2446), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(n952), .B(n951), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(n954), .B(n953), .ZN(n955) );
  NAND2_X1 U1045 ( .A1(n955), .A2(G14), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(KEYINPUT103), .B(n956), .ZN(G401) );
  XOR2_X1 U1047 ( .A(G2678), .B(G2084), .Z(n958) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G2078), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(n958), .B(n957), .ZN(n959) );
  XOR2_X1 U1050 ( .A(n959), .B(KEYINPUT107), .Z(n961) );
  XNOR2_X1 U1051 ( .A(G2072), .B(KEYINPUT42), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n961), .B(n960), .ZN(n965) );
  XOR2_X1 U1053 ( .A(G2100), .B(G2096), .Z(n963) );
  XNOR2_X1 U1054 ( .A(G2090), .B(KEYINPUT43), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n963), .B(n962), .ZN(n964) );
  XOR2_X1 U1056 ( .A(n965), .B(n964), .Z(G227) );
  XNOR2_X1 U1057 ( .A(G1986), .B(G1976), .ZN(n975) );
  XOR2_X1 U1058 ( .A(G1971), .B(G1956), .Z(n967) );
  XNOR2_X1 U1059 ( .A(G1996), .B(G1966), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n967), .B(n966), .ZN(n971) );
  XOR2_X1 U1061 ( .A(KEYINPUT108), .B(G2474), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G1991), .B(G1981), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1064 ( .A(n971), .B(n970), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G1961), .B(KEYINPUT41), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(G229) );
  XNOR2_X1 U1068 ( .A(G160), .B(G162), .ZN(n1004) );
  XOR2_X1 U1069 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(n977), .B(n976), .ZN(n978) );
  XOR2_X1 U1072 ( .A(n978), .B(KEYINPUT115), .Z(n993) );
  NAND2_X1 U1073 ( .A1(G118), .A2(n979), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(G130), .A2(n980), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(G106), .A2(n983), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(G142), .A2(n984), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT45), .B(n987), .Z(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT110), .B(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n991), .B(KEYINPUT114), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(n993), .B(n992), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(n994), .ZN(n997) );
  XOR2_X1 U1085 ( .A(n997), .B(n996), .Z(n999) );
  XOR2_X1 U1086 ( .A(n999), .B(n998), .Z(n1002) );
  XOR2_X1 U1087 ( .A(G164), .B(n1000), .Z(n1001) );
  XNOR2_X1 U1088 ( .A(n1002), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(n1004), .B(n1003), .ZN(n1006) );
  XOR2_X1 U1090 ( .A(n1006), .B(n1005), .Z(n1007) );
  NOR2_X1 U1091 ( .A1(G37), .A2(n1007), .ZN(G395) );
  XOR2_X1 U1092 ( .A(n1008), .B(G286), .Z(n1011) );
  XNOR2_X1 U1093 ( .A(n1009), .B(G171), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(n1012), .B(n680), .ZN(n1013) );
  NOR2_X1 U1096 ( .A1(G37), .A2(n1013), .ZN(G397) );
  XOR2_X1 U1097 ( .A(KEYINPUT106), .B(n1014), .Z(G319) );
  NOR2_X1 U1098 ( .A1(G227), .A2(G229), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(KEYINPUT49), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1100 ( .A1(G401), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1101 ( .A1(G395), .A2(G397), .ZN(n1017) );
  AND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(G319), .ZN(G225) );
  INV_X1 U1104 ( .A(G225), .ZN(G308) );
  INV_X1 U1105 ( .A(G303), .ZN(G166) );
  INV_X1 U1106 ( .A(G108), .ZN(G238) );
endmodule

