

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n703), .B(n702), .ZN(n709) );
  NOR2_X1 U552 ( .A1(n525), .A2(n524), .ZN(G160) );
  NOR2_X2 U553 ( .A1(n768), .A2(n767), .ZN(n769) );
  AND2_X4 U554 ( .A1(n521), .A2(G2104), .ZN(n561) );
  INV_X2 U555 ( .A(G2105), .ZN(n521) );
  AND2_X1 U556 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U557 ( .A1(n735), .A2(n945), .ZN(n679) );
  AND2_X1 U558 ( .A1(n978), .A2(n748), .ZN(n749) );
  NOR2_X2 U559 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XOR2_X2 U560 ( .A(KEYINPUT17), .B(n520), .Z(n875) );
  XOR2_X1 U561 ( .A(KEYINPUT13), .B(n588), .Z(n515) );
  XNOR2_X1 U562 ( .A(KEYINPUT30), .B(KEYINPUT95), .ZN(n715) );
  XNOR2_X1 U563 ( .A(n716), .B(n715), .ZN(n717) );
  INV_X1 U564 ( .A(KEYINPUT97), .ZN(n730) );
  INV_X1 U565 ( .A(n764), .ZN(n748) );
  INV_X1 U566 ( .A(n983), .ZN(n753) );
  OR2_X1 U567 ( .A1(n754), .A2(n753), .ZN(n755) );
  INV_X1 U568 ( .A(KEYINPUT73), .ZN(n596) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NOR2_X2 U570 ( .A1(G651), .A2(n626), .ZN(n644) );
  INV_X1 U571 ( .A(KEYINPUT23), .ZN(n516) );
  XNOR2_X1 U572 ( .A(n517), .B(n516), .ZN(n518) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U574 ( .A1(n879), .A2(G113), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n561), .A2(G101), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n519), .A2(n518), .ZN(n525) );
  NAND2_X1 U577 ( .A1(G137), .A2(n875), .ZN(n523) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n521), .ZN(n878) );
  NAND2_X1 U579 ( .A1(G125), .A2(n878), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n523), .A2(n522), .ZN(n524) );
  INV_X1 U581 ( .A(G651), .ZN(n531) );
  NOR2_X1 U582 ( .A1(G543), .A2(n531), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n526), .Z(n583) );
  BUF_X1 U584 ( .A(n583), .Z(n643) );
  NAND2_X1 U585 ( .A1(G63), .A2(n643), .ZN(n528) );
  NAND2_X1 U586 ( .A1(G51), .A2(n644), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U588 ( .A(KEYINPUT6), .B(n529), .ZN(n537) );
  NOR2_X2 U589 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U590 ( .A1(n639), .A2(G89), .ZN(n530) );
  XNOR2_X1 U591 ( .A(n530), .B(KEYINPUT4), .ZN(n533) );
  NOR2_X2 U592 ( .A1(n626), .A2(n531), .ZN(n640) );
  NAND2_X1 U593 ( .A1(G76), .A2(n640), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U595 ( .A(KEYINPUT74), .B(n534), .Z(n535) );
  XNOR2_X1 U596 ( .A(KEYINPUT5), .B(n535), .ZN(n536) );
  NOR2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U598 ( .A(KEYINPUT7), .B(n538), .Z(G168) );
  XOR2_X1 U599 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U600 ( .A1(G85), .A2(n639), .ZN(n540) );
  NAND2_X1 U601 ( .A1(G72), .A2(n640), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U603 ( .A1(G60), .A2(n643), .ZN(n542) );
  NAND2_X1 U604 ( .A1(G47), .A2(n644), .ZN(n541) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U606 ( .A1(n544), .A2(n543), .ZN(G290) );
  NAND2_X1 U607 ( .A1(G90), .A2(n639), .ZN(n546) );
  NAND2_X1 U608 ( .A1(G77), .A2(n640), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G64), .A2(n643), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n644), .A2(G52), .ZN(n550) );
  XOR2_X1 U614 ( .A(KEYINPUT64), .B(n550), .Z(n551) );
  NOR2_X1 U615 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U616 ( .A1(G135), .A2(n875), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G111), .A2(n879), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n878), .A2(G123), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT18), .B(n555), .Z(n556) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n561), .A2(G99), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n920) );
  XNOR2_X1 U624 ( .A(G2096), .B(n920), .ZN(n560) );
  OR2_X1 U625 ( .A1(G2100), .A2(n560), .ZN(G156) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  NAND2_X1 U628 ( .A1(n875), .A2(G138), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G102), .A2(n561), .ZN(n562) );
  XOR2_X1 U630 ( .A(KEYINPUT85), .B(n562), .Z(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G126), .A2(n878), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G114), .A2(n879), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(G164) );
  NAND2_X1 U636 ( .A1(G91), .A2(n639), .ZN(n570) );
  NAND2_X1 U637 ( .A1(G78), .A2(n640), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(KEYINPUT66), .B(n571), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G53), .A2(n644), .ZN(n572) );
  XNOR2_X1 U641 ( .A(KEYINPUT67), .B(n572), .ZN(n573) );
  NOR2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n643), .A2(G65), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U645 ( .A(KEYINPUT68), .B(n577), .ZN(G299) );
  NAND2_X1 U646 ( .A1(G94), .A2(G452), .ZN(n578) );
  XNOR2_X1 U647 ( .A(n578), .B(KEYINPUT65), .ZN(G173) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U649 ( .A(n579), .B(KEYINPUT10), .ZN(n580) );
  XNOR2_X1 U650 ( .A(KEYINPUT70), .B(n580), .ZN(G223) );
  INV_X1 U651 ( .A(G223), .ZN(n819) );
  NAND2_X1 U652 ( .A1(n819), .A2(G567), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n581), .B(KEYINPUT71), .ZN(n582) );
  XNOR2_X1 U654 ( .A(KEYINPUT11), .B(n582), .ZN(G234) );
  NAND2_X1 U655 ( .A1(G56), .A2(n583), .ZN(n584) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(n584), .Z(n589) );
  NAND2_X1 U657 ( .A1(n639), .A2(G81), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT12), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G68), .A2(n640), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n589), .A2(n515), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n644), .A2(G43), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n971) );
  INV_X1 U664 ( .A(G860), .ZN(n613) );
  OR2_X1 U665 ( .A1(n971), .A2(n613), .ZN(G153) );
  XOR2_X1 U666 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U668 ( .A1(G66), .A2(n643), .ZN(n593) );
  NAND2_X1 U669 ( .A1(G92), .A2(n639), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G54), .A2(n644), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G79), .A2(n640), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n597) );
  XNOR2_X1 U674 ( .A(n597), .B(n596), .ZN(n598) );
  NOR2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X2 U676 ( .A(KEYINPUT15), .B(n600), .Z(n892) );
  INV_X1 U677 ( .A(n892), .ZN(n964) );
  INV_X1 U678 ( .A(G868), .ZN(n659) );
  NAND2_X1 U679 ( .A1(n964), .A2(n659), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n602), .A2(n601), .ZN(G284) );
  NOR2_X1 U681 ( .A1(G286), .A2(n659), .ZN(n603) );
  XOR2_X1 U682 ( .A(KEYINPUT75), .B(n603), .Z(n605) );
  NOR2_X1 U683 ( .A1(G299), .A2(G868), .ZN(n604) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U685 ( .A1(G559), .A2(n613), .ZN(n606) );
  XNOR2_X1 U686 ( .A(KEYINPUT76), .B(n606), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n607), .A2(n892), .ZN(n608) );
  XNOR2_X1 U688 ( .A(KEYINPUT16), .B(n608), .ZN(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n971), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n892), .A2(G868), .ZN(n609) );
  NOR2_X1 U691 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U692 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G559), .A2(n892), .ZN(n612) );
  XOR2_X1 U694 ( .A(n971), .B(n612), .Z(n655) );
  NAND2_X1 U695 ( .A1(n613), .A2(n655), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G67), .A2(n643), .ZN(n615) );
  NAND2_X1 U697 ( .A1(G93), .A2(n639), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G80), .A2(n640), .ZN(n617) );
  NAND2_X1 U700 ( .A1(G55), .A2(n644), .ZN(n616) );
  NAND2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n658) );
  XOR2_X1 U703 ( .A(n620), .B(n658), .Z(G145) );
  NAND2_X1 U704 ( .A1(n644), .A2(G49), .ZN(n621) );
  XOR2_X1 U705 ( .A(KEYINPUT77), .B(n621), .Z(n623) );
  NAND2_X1 U706 ( .A1(G651), .A2(G74), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U708 ( .A1(n643), .A2(n624), .ZN(n625) );
  XNOR2_X1 U709 ( .A(n625), .B(KEYINPUT78), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n626), .A2(G87), .ZN(n627) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(n627), .Z(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n630), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G73), .A2(n640), .ZN(n631) );
  XNOR2_X1 U715 ( .A(n631), .B(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G86), .A2(n639), .ZN(n633) );
  NAND2_X1 U717 ( .A1(G48), .A2(n644), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G61), .A2(n643), .ZN(n634) );
  XNOR2_X1 U720 ( .A(KEYINPUT81), .B(n634), .ZN(n635) );
  NOR2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G88), .A2(n639), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G75), .A2(n640), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n648) );
  NAND2_X1 U726 ( .A1(G62), .A2(n643), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G50), .A2(n644), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U729 ( .A1(n648), .A2(n647), .ZN(G166) );
  XOR2_X1 U730 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n649) );
  XNOR2_X1 U731 ( .A(G305), .B(n649), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n658), .B(n650), .ZN(n652) );
  XNOR2_X1 U733 ( .A(G290), .B(G166), .ZN(n651) );
  XNOR2_X1 U734 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U735 ( .A(G288), .B(n653), .Z(n654) );
  XNOR2_X1 U736 ( .A(G299), .B(n654), .ZN(n895) );
  XOR2_X1 U737 ( .A(n655), .B(n895), .Z(n656) );
  XNOR2_X1 U738 ( .A(KEYINPUT83), .B(n656), .ZN(n657) );
  NOR2_X1 U739 ( .A1(n659), .A2(n657), .ZN(n661) );
  AND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U741 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U748 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U749 ( .A1(G219), .A2(G220), .ZN(n666) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U751 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(G96), .A2(n668), .ZN(n826) );
  NAND2_X1 U753 ( .A1(n826), .A2(G2106), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G120), .A2(G69), .ZN(n669) );
  NOR2_X1 U755 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U756 ( .A1(G108), .A2(n670), .ZN(n827) );
  NAND2_X1 U757 ( .A1(n827), .A2(G567), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n672), .A2(n671), .ZN(n849) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n673) );
  XNOR2_X1 U760 ( .A(KEYINPUT84), .B(n673), .ZN(n674) );
  NOR2_X1 U761 ( .A1(n849), .A2(n674), .ZN(n825) );
  NAND2_X1 U762 ( .A1(n825), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U765 ( .A(n770), .ZN(n676) );
  NOR2_X2 U766 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X2 U767 ( .A1(n676), .A2(n771), .ZN(n735) );
  AND2_X1 U768 ( .A1(n735), .A2(G1341), .ZN(n677) );
  NOR2_X1 U769 ( .A1(n971), .A2(n677), .ZN(n681) );
  INV_X1 U770 ( .A(G1996), .ZN(n945) );
  INV_X1 U771 ( .A(KEYINPUT26), .ZN(n678) );
  XNOR2_X1 U772 ( .A(n679), .B(n678), .ZN(n680) );
  AND2_X1 U773 ( .A1(n681), .A2(n680), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n687), .A2(n892), .ZN(n685) );
  INV_X1 U775 ( .A(n735), .ZN(n705) );
  NOR2_X1 U776 ( .A1(n705), .A2(G1348), .ZN(n683) );
  NOR2_X1 U777 ( .A1(G2067), .A2(n735), .ZN(n682) );
  NOR2_X1 U778 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U780 ( .A(KEYINPUT93), .B(n686), .Z(n689) );
  OR2_X1 U781 ( .A1(n892), .A2(n687), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n695) );
  XOR2_X1 U783 ( .A(KEYINPUT91), .B(KEYINPUT27), .Z(n691) );
  NAND2_X1 U784 ( .A1(G2072), .A2(n705), .ZN(n690) );
  XNOR2_X1 U785 ( .A(n691), .B(n690), .ZN(n693) );
  INV_X1 U786 ( .A(G1956), .ZN(n992) );
  NOR2_X1 U787 ( .A1(n705), .A2(n992), .ZN(n692) );
  NOR2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n697) );
  INV_X1 U789 ( .A(G299), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n701) );
  NOR2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n699) );
  XOR2_X1 U793 ( .A(KEYINPUT92), .B(KEYINPUT28), .Z(n698) );
  XNOR2_X1 U794 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n703) );
  XOR2_X1 U796 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n702) );
  XNOR2_X1 U797 ( .A(G1961), .B(KEYINPUT89), .ZN(n991) );
  NAND2_X1 U798 ( .A1(n735), .A2(n991), .ZN(n707) );
  XNOR2_X1 U799 ( .A(G2078), .B(KEYINPUT90), .ZN(n704) );
  XNOR2_X1 U800 ( .A(n704), .B(KEYINPUT25), .ZN(n949) );
  NAND2_X1 U801 ( .A1(n705), .A2(n949), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n718) );
  NAND2_X1 U803 ( .A1(n718), .A2(G171), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n723) );
  NOR2_X1 U805 ( .A1(n735), .A2(G2084), .ZN(n711) );
  INV_X1 U806 ( .A(KEYINPUT88), .ZN(n710) );
  XNOR2_X1 U807 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n712), .A2(G8), .ZN(n714) );
  NAND2_X1 U809 ( .A1(G8), .A2(n735), .ZN(n764) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n764), .ZN(n713) );
  NOR2_X1 U811 ( .A1(n714), .A2(n713), .ZN(n716) );
  NOR2_X1 U812 ( .A1(n717), .A2(G168), .ZN(n720) );
  NOR2_X1 U813 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U815 ( .A(n721), .B(KEYINPUT31), .Z(n722) );
  NAND2_X1 U816 ( .A1(n723), .A2(n722), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n740), .A2(G286), .ZN(n729) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n764), .ZN(n725) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n735), .ZN(n724) );
  NOR2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U821 ( .A(KEYINPUT96), .B(n726), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n727), .A2(G303), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n731) );
  XNOR2_X1 U824 ( .A(n731), .B(n730), .ZN(n732) );
  NAND2_X1 U825 ( .A1(n732), .A2(G8), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n733), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U827 ( .A1(KEYINPUT88), .A2(G1966), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n734), .A2(n735), .ZN(n738) );
  XOR2_X1 U829 ( .A(KEYINPUT88), .B(G2084), .Z(n736) );
  NAND2_X1 U830 ( .A1(n736), .A2(n705), .ZN(n737) );
  NAND2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n739), .A2(G8), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n759) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NOR2_X1 U836 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U837 ( .A1(n977), .A2(n744), .ZN(n745) );
  NAND2_X1 U838 ( .A1(n759), .A2(n745), .ZN(n746) );
  XNOR2_X1 U839 ( .A(n746), .B(KEYINPUT98), .ZN(n750) );
  NAND2_X1 U840 ( .A1(G288), .A2(G1976), .ZN(n747) );
  XOR2_X1 U841 ( .A(KEYINPUT99), .B(n747), .Z(n978) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n751), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n977), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n752), .A2(n764), .ZN(n754) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n983) );
  NOR2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n768) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n757) );
  XNOR2_X1 U848 ( .A(n757), .B(KEYINPUT100), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n758), .A2(G8), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n761), .A2(n764), .ZN(n766) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U853 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  OR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U856 ( .A(n769), .B(KEYINPUT101), .ZN(n801) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n815) );
  NAND2_X1 U858 ( .A1(G95), .A2(n561), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G119), .A2(n878), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G131), .A2(n875), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G107), .A2(n879), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U865 ( .A(n778), .B(KEYINPUT87), .ZN(n889) );
  NAND2_X1 U866 ( .A1(G1991), .A2(n889), .ZN(n787) );
  NAND2_X1 U867 ( .A1(G141), .A2(n875), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G117), .A2(n879), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n561), .A2(G105), .ZN(n781) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n878), .A2(G129), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n869) );
  NAND2_X1 U875 ( .A1(G1996), .A2(n869), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n923) );
  NAND2_X1 U877 ( .A1(n815), .A2(n923), .ZN(n805) );
  XNOR2_X1 U878 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U879 ( .A1(n815), .A2(n968), .ZN(n788) );
  AND2_X1 U880 ( .A1(n805), .A2(n788), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G104), .A2(n561), .ZN(n790) );
  NAND2_X1 U882 ( .A1(G140), .A2(n875), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n791), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G128), .A2(n878), .ZN(n793) );
  NAND2_X1 U886 ( .A1(G116), .A2(n879), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U888 ( .A(n794), .B(KEYINPUT35), .Z(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U890 ( .A(KEYINPUT36), .B(n797), .Z(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT86), .B(n798), .Z(n885) );
  XNOR2_X1 U892 ( .A(KEYINPUT37), .B(G2067), .ZN(n812) );
  NOR2_X1 U893 ( .A1(n885), .A2(n812), .ZN(n916) );
  NAND2_X1 U894 ( .A1(n815), .A2(n916), .ZN(n809) );
  AND2_X1 U895 ( .A1(n799), .A2(n809), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U897 ( .A(n802), .B(KEYINPUT102), .ZN(n817) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n889), .ZN(n919) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n919), .A2(n803), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n804), .B(KEYINPUT103), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U903 ( .A1(n869), .A2(G1996), .ZN(n930) );
  NAND2_X1 U904 ( .A1(n807), .A2(n930), .ZN(n808) );
  XOR2_X1 U905 ( .A(KEYINPUT39), .B(n808), .Z(n810) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(KEYINPUT104), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n885), .A2(n812), .ZN(n915) );
  NAND2_X1 U909 ( .A1(n813), .A2(n915), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(n819), .A2(G2106), .ZN(n820) );
  XOR2_X1 U914 ( .A(KEYINPUT105), .B(n820), .Z(G217) );
  INV_X1 U915 ( .A(G661), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G2), .A2(G15), .ZN(n821) );
  NOR2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U918 ( .A(KEYINPUT106), .B(n823), .Z(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XOR2_X1 U927 ( .A(G1981), .B(G1966), .Z(n829) );
  XNOR2_X1 U928 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U929 ( .A(n829), .B(n828), .ZN(n839) );
  XOR2_X1 U930 ( .A(KEYINPUT41), .B(G2474), .Z(n831) );
  XNOR2_X1 U931 ( .A(G1956), .B(KEYINPUT109), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U933 ( .A(G1976), .B(G1971), .Z(n833) );
  XNOR2_X1 U934 ( .A(G1986), .B(G1961), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U936 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U937 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U939 ( .A(n839), .B(n838), .Z(G229) );
  XOR2_X1 U940 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2067), .B(KEYINPUT108), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n842), .B(G2678), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2072), .B(G2090), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2100), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(G227) );
  INV_X1 U950 ( .A(n849), .ZN(G319) );
  NAND2_X1 U951 ( .A1(G124), .A2(n878), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n850), .B(KEYINPUT112), .ZN(n851) );
  XNOR2_X1 U953 ( .A(KEYINPUT44), .B(n851), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G136), .A2(n875), .ZN(n852) );
  XOR2_X1 U955 ( .A(KEYINPUT113), .B(n852), .Z(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G100), .A2(n561), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G112), .A2(n879), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U960 ( .A1(n858), .A2(n857), .ZN(G162) );
  NAND2_X1 U961 ( .A1(G130), .A2(n878), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G118), .A2(n879), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G106), .A2(n561), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G142), .A2(n875), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U967 ( .A(n863), .B(KEYINPUT45), .Z(n864) );
  NOR2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n866), .B(n920), .ZN(n874) );
  XOR2_X1 U970 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n867) );
  XNOR2_X1 U972 ( .A(n868), .B(n867), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n872) );
  XNOR2_X1 U974 ( .A(G164), .B(G160), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U976 ( .A(n874), .B(n873), .Z(n887) );
  NAND2_X1 U977 ( .A1(G103), .A2(n561), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G139), .A2(n875), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G127), .A2(n878), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G115), .A2(n879), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n926) );
  XNOR2_X1 U985 ( .A(n885), .B(n926), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(G162), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U989 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U990 ( .A(n971), .B(G286), .ZN(n894) );
  XNOR2_X1 U991 ( .A(G171), .B(n892), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G397) );
  NOR2_X1 U995 ( .A1(G229), .A2(G227), .ZN(n899) );
  XNOR2_X1 U996 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(KEYINPUT49), .B(n900), .Z(n911) );
  XOR2_X1 U999 ( .A(G2451), .B(G2430), .Z(n902) );
  XNOR2_X1 U1000 ( .A(G2438), .B(G2443), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n908) );
  XOR2_X1 U1002 ( .A(G2435), .B(G2454), .Z(n904) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1005 ( .A(G2446), .B(G2427), .Z(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1007 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1008 ( .A1(G14), .A2(n909), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n914), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n914), .ZN(G401) );
  INV_X1 U1016 ( .A(n915), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n925) );
  XOR2_X1 U1018 ( .A(G160), .B(G2084), .Z(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n936) );
  XOR2_X1 U1023 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT50), .B(n929), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G162), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT51), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n937), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n959) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n959), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n939), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1036 ( .A(KEYINPUT119), .B(G2090), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n940), .B(G35), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT120), .B(G34), .Z(n942) );
  XNOR2_X1 U1039 ( .A(G2084), .B(KEYINPUT54), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n942), .B(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n958) );
  XNOR2_X1 U1042 ( .A(G32), .B(n945), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n946), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1044 ( .A(G1991), .B(G25), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n953) );
  XOR2_X1 U1047 ( .A(n949), .B(G27), .Z(n951) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT53), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n960), .B(n959), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(G29), .A2(n961), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT121), .B(n962), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(G11), .ZN(n1019) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1059 ( .A(n964), .B(G1348), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G299), .B(G1956), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n976) );
  XNOR2_X1 U1062 ( .A(G171), .B(G1961), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G303), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n971), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT124), .B(n972), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(KEYINPUT123), .B(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1073 ( .A(KEYINPUT125), .B(n982), .Z(n988) );
  XNOR2_X1 U1074 ( .A(G168), .B(G1966), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n985), .B(KEYINPUT57), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(KEYINPUT122), .B(n986), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n1017) );
  INV_X1 U1080 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1081 ( .A(G5), .B(n991), .ZN(n1004) );
  XNOR2_X1 U1082 ( .A(G20), .B(n992), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G6), .B(G1981), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1087 ( .A(KEYINPUT59), .B(G1348), .Z(n997) );
  XNOR2_X1 U1088 ( .A(G4), .B(n997), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1000), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G1986), .B(KEYINPUT126), .Z(n1007) );
  XNOR2_X1 U1098 ( .A(G24), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT62), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(KEYINPUT127), .B(n1023), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

