//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT65), .B(G244), .Z(new_n209));
  AND2_X1   g0009(.A1(new_n209), .A2(G77), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G87), .A2(G250), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n205), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT64), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n220), .A2(G1), .A3(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n208), .B(new_n217), .C1(new_n224), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G97), .B(G107), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G223), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n246), .A2(new_n248), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G222), .A3(new_n250), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n249), .A2(G77), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n256), .B2(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(G1), .B(G13), .C1(new_n245), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT71), .B(G179), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n222), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G58), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(KEYINPUT8), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n278), .A2(KEYINPUT8), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(KEYINPUT69), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(KEYINPUT69), .B2(new_n280), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n245), .A2(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n202), .A2(G20), .B1(G150), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n277), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n262), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n277), .A2(new_n289), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G50), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n295), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n288), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n271), .B1(new_n257), .B2(new_n260), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G169), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n275), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  AOI211_X1 g0104(.A(KEYINPUT9), .B(new_n288), .C1(new_n297), .C2(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n304), .A2(new_n305), .B1(new_n306), .B2(new_n273), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT73), .B1(new_n273), .B2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n300), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n298), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n296), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT9), .B1(new_n315), .B2(new_n288), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n299), .A2(new_n303), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n316), .A2(new_n317), .B1(G190), .B2(new_n300), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n308), .A2(new_n311), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n302), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G232), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n249), .A2(new_n323), .A3(new_n250), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n246), .A2(new_n248), .A3(G226), .A4(new_n250), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G33), .A2(G97), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n258), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  INV_X1    g0129(.A(new_n269), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n265), .B1(new_n330), .B2(G238), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n329), .B1(new_n328), .B2(new_n331), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G190), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n334), .A2(new_n310), .ZN(new_n338));
  INV_X1    g0138(.A(new_n291), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n277), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT72), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n222), .A2(new_n276), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n291), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n342), .A2(new_n345), .B1(new_n262), .B2(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G68), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n286), .A2(G50), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  INV_X1    g0149(.A(new_n284), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n348), .B1(new_n223), .B2(G68), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n343), .ZN(new_n352));
  INV_X1    g0152(.A(G68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n291), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT12), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT11), .B1(new_n351), .B2(new_n343), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n338), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n336), .A2(new_n337), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT75), .B1(new_n334), .B2(G179), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n332), .A2(new_n333), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT14), .B1(new_n334), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(G169), .C1(new_n332), .C2(new_n333), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT76), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n368), .B(new_n370), .C1(new_n362), .C2(new_n365), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT76), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n359), .B(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n265), .B1(new_n330), .B2(new_n209), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n251), .A2(G238), .B1(G107), .B2(new_n249), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n253), .A2(G232), .A3(new_n250), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n379), .B1(new_n382), .B2(new_n259), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G200), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n306), .B2(new_n383), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n346), .A2(G77), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n281), .A2(new_n279), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n350), .B2(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n343), .B1(new_n349), .B2(new_n291), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n383), .A2(new_n274), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n383), .A2(new_n367), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n322), .A2(new_n361), .A3(new_n378), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n270), .A2(new_n250), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n246), .B(new_n400), .C1(new_n401), .C2(new_n245), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT80), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n247), .A2(KEYINPUT78), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G33), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(G223), .A3(new_n250), .A4(new_n246), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n409), .A2(KEYINPUT80), .A3(new_n246), .A4(new_n400), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n404), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n258), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n266), .B1(new_n269), .B2(new_n323), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT81), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n413), .B2(new_n258), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT81), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n367), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(G58), .B(G68), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(G20), .B1(G159), .B2(new_n286), .ZN(new_n424));
  INV_X1    g0224(.A(new_n246), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n408), .B2(G33), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT7), .B1(new_n426), .B2(G20), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G68), .ZN(new_n428));
  NOR2_X1   g0228(.A1(KEYINPUT7), .A2(G20), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n246), .B1(new_n401), .B2(new_n245), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT79), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n409), .A2(new_n433), .A3(new_n246), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(KEYINPUT16), .B(new_n424), .C1(new_n428), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n223), .A2(KEYINPUT7), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n401), .A2(new_n245), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(new_n248), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT7), .B1(new_n249), .B2(new_n223), .ZN(new_n440));
  OAI21_X1  g0240(.A(G68), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n424), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT16), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n436), .A2(new_n444), .A3(new_n343), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n293), .A2(new_n283), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n283), .B2(new_n291), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n419), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n422), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n422), .A2(new_n448), .A3(KEYINPUT18), .A4(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n445), .A2(new_n447), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n419), .A2(new_n420), .ZN(new_n459));
  AOI211_X1 g0259(.A(KEYINPUT81), .B(new_n415), .C1(new_n413), .C2(new_n258), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n459), .A2(new_n460), .A3(G200), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n417), .A2(G190), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n457), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n418), .A2(new_n310), .A3(new_n421), .ZN(new_n466));
  INV_X1    g0266(.A(new_n462), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n448), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n457), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n455), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n399), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n262), .A2(G33), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G116), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n345), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT20), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  INV_X1    g0281(.A(G97), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(new_n223), .C1(G33), .C2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n223), .B2(G116), .ZN(new_n484));
  OR3_X1    g0284(.A1(new_n277), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n480), .B1(new_n277), .B2(new_n484), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n291), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G257), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n250), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G264), .B2(new_n250), .ZN(new_n492));
  INV_X1    g0292(.A(G303), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n431), .A2(new_n492), .B1(new_n493), .B2(new_n253), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT89), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT89), .ZN(new_n496));
  OAI221_X1 g0296(.A(new_n496), .B1(new_n493), .B2(new_n253), .C1(new_n431), .C2(new_n492), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n258), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT5), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G41), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G1), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n267), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n264), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n505), .A2(new_n268), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G270), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n367), .B1(new_n498), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n489), .A2(new_n509), .A3(KEYINPUT91), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT91), .B1(new_n489), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n473), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n498), .A2(new_n508), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n489), .B1(G200), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n306), .B2(new_n513), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(KEYINPUT21), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n498), .A2(G179), .A3(new_n508), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT90), .B1(new_n518), .B2(new_n489), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT90), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n479), .A2(new_n488), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n516), .C2(new_n517), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n512), .B(new_n515), .C1(new_n519), .C2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G107), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n291), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n525), .B(KEYINPUT25), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n344), .A2(new_n474), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(G107), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT93), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT23), .B1(new_n223), .B2(G107), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT94), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n223), .A2(G87), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n249), .B2(new_n534), .ZN(new_n535));
  OR3_X1    g0335(.A1(new_n223), .A2(KEYINPUT23), .A3(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n409), .A2(KEYINPUT22), .A3(G87), .A4(new_n246), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n529), .B(new_n538), .C1(new_n541), .C2(G20), .ZN(new_n542));
  AOI21_X1  g0342(.A(G20), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT93), .B1(new_n543), .B2(new_n537), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT24), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n343), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT24), .B1(new_n542), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n528), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n506), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G250), .A2(G1698), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n490), .B2(G1698), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n426), .A2(new_n551), .B1(G33), .B2(G294), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(new_n259), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n505), .A2(G264), .A3(new_n268), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G169), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT95), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n554), .B(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n553), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n556), .B1(new_n560), .B2(new_n364), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n548), .A2(new_n561), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n555), .A2(G190), .B1(new_n559), .B2(G200), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n563), .B(new_n528), .C1(new_n546), .C2(new_n547), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n250), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n481), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n426), .A2(G244), .A3(new_n250), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n570), .A2(new_n259), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n507), .A2(G257), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n571), .A2(new_n449), .A3(new_n549), .A4(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n339), .A2(G97), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n527), .B2(G97), .ZN(new_n575));
  OAI21_X1  g0375(.A(G107), .B1(new_n439), .B2(new_n440), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n524), .A2(KEYINPUT6), .A3(G97), .ZN(new_n577));
  INV_X1    g0377(.A(new_n242), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(KEYINPUT6), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT83), .B1(new_n581), .B2(new_n343), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n583), .B(new_n277), .C1(new_n576), .C2(new_n580), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n575), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n549), .B(new_n572), .C1(new_n570), .C2(new_n259), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n367), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n573), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n586), .A2(new_n306), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n582), .A2(new_n584), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(G200), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n575), .A4(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n562), .A2(new_n564), .A3(new_n588), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT86), .ZN(new_n595));
  OAI211_X1 g0395(.A(G244), .B(new_n246), .C1(new_n401), .C2(new_n245), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n250), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n426), .A2(KEYINPUT86), .A3(G244), .A4(G1698), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n426), .A2(G238), .A3(new_n250), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n540), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n258), .ZN(new_n601));
  INV_X1    g0401(.A(G250), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n503), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n268), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT85), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n503), .B2(G274), .ZN(new_n606));
  NOR4_X1   g0406(.A1(new_n502), .A2(new_n264), .A3(KEYINPUT85), .A4(G1), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n594), .B1(new_n601), .B2(new_n609), .ZN(new_n610));
  AOI211_X1 g0410(.A(KEYINPUT87), .B(new_n608), .C1(new_n600), .C2(new_n258), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n449), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n390), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n527), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n223), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(KEYINPUT88), .A3(new_n223), .ZN(new_n619));
  INV_X1    g0419(.A(G87), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n482), .A3(new_n524), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n353), .A2(G20), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n246), .B(new_n623), .C1(new_n401), .C2(new_n245), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT19), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n350), .B2(new_n482), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n343), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n291), .A2(new_n390), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n614), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n601), .A2(new_n609), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT87), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n601), .A2(new_n594), .A3(new_n609), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n612), .B(new_n630), .C1(new_n634), .C2(G169), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(G200), .A3(new_n633), .ZN(new_n636));
  OAI21_X1  g0436(.A(G190), .B1(new_n610), .B2(new_n611), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n344), .A2(G87), .A3(new_n474), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n628), .A2(new_n629), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n523), .A2(new_n593), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n472), .A2(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n518), .A2(new_n489), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n562), .A2(new_n512), .A3(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n592), .A2(new_n564), .A3(new_n588), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n631), .A2(new_n367), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n612), .A2(new_n630), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n639), .A2(KEYINPUT96), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT96), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n628), .A2(new_n651), .A3(new_n629), .A4(new_n638), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n310), .B1(new_n601), .B2(new_n609), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n637), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n649), .A2(KEYINPUT97), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT97), .B1(new_n649), .B2(new_n656), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n646), .B(new_n647), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n573), .A2(new_n585), .A3(new_n587), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n660), .B(new_n661), .C1(new_n657), .C2(new_n658), .ZN(new_n662));
  INV_X1    g0462(.A(new_n649), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n635), .A2(new_n641), .A3(new_n661), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(KEYINPUT26), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n472), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n397), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n361), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n378), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n464), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n469), .B1(new_n468), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n463), .A2(new_n457), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n455), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n313), .A2(new_n321), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n302), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n667), .A2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n512), .A2(new_n645), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n290), .A2(G20), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n262), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n521), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n680), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n523), .B2(new_n689), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n562), .A2(new_n564), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n548), .A2(new_n687), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n562), .B2(new_n688), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n562), .A2(new_n687), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n519), .A2(new_n522), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n687), .B1(new_n699), .B2(new_n512), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n206), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n621), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n225), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n666), .A2(new_n710), .A3(new_n688), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n664), .A2(new_n660), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT100), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT26), .B(new_n661), .C1(new_n657), .C2(new_n658), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n664), .A2(KEYINPUT100), .A3(new_n660), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n512), .B(new_n562), .C1(new_n519), .C2(new_n522), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(new_n647), .C1(new_n658), .C2(new_n657), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n649), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n688), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n711), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n571), .A2(new_n559), .A3(new_n572), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT98), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n517), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n517), .A2(new_n724), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n634), .A2(new_n723), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n559), .A2(new_n274), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n513), .A3(new_n631), .A4(new_n586), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n727), .B2(new_n728), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n688), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n593), .A2(new_n642), .ZN(new_n736));
  INV_X1    g0536(.A(new_n523), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(new_n688), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n735), .B1(new_n738), .B2(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n687), .A2(KEYINPUT31), .ZN(new_n740));
  INV_X1    g0540(.A(new_n734), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n729), .B1(new_n741), .B2(KEYINPUT99), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT99), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n734), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n740), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(G330), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n722), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n709), .B1(new_n748), .B2(G1), .ZN(G364));
  AOI21_X1  g0549(.A(new_n262), .B1(new_n681), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n704), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n692), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n691), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n222), .B1(G20), .B2(new_n367), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n240), .A2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n432), .ZN(new_n762));
  INV_X1    g0562(.A(new_n434), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n703), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n761), .B(new_n765), .C1(G45), .C2(new_n225), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n703), .A2(new_n249), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G355), .B1(new_n487), .B2(new_n703), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n760), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n755), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n223), .A2(G179), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n310), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G190), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G283), .A2(new_n774), .B1(new_n777), .B2(G329), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n306), .A2(new_n310), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n771), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n249), .C1(new_n493), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n306), .A2(G200), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n223), .B1(new_n782), .B2(new_n364), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n781), .B1(G294), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n274), .A2(G20), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n782), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n779), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G322), .A2(new_n789), .B1(new_n791), .B2(G326), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n775), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n787), .A2(new_n772), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G311), .A2(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n785), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G58), .A2(new_n789), .B1(new_n794), .B2(G77), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n773), .A2(new_n524), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n253), .B1(new_n780), .B2(new_n620), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G97), .C2(new_n784), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n791), .A2(G50), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT32), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n776), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n777), .A2(KEYINPUT32), .A3(G159), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n796), .A2(G68), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n770), .B1(new_n799), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n752), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n769), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n758), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n691), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n754), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n393), .A2(new_n687), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n394), .A2(new_n397), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT104), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n397), .A2(new_n688), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n666), .B2(new_n688), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n666), .A2(new_n688), .A3(new_n820), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT105), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n666), .A2(KEYINPUT105), .A3(new_n688), .A4(new_n820), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n746), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT106), .ZN(new_n830));
  OR3_X1    g0630(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n828), .B2(new_n829), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n752), .B1(new_n828), .B2(new_n829), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n755), .A2(new_n756), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n752), .B1(new_n836), .B2(G77), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT102), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G116), .A2(new_n794), .B1(new_n791), .B2(G303), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G283), .A2(new_n796), .B1(new_n789), .B2(G294), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n249), .B1(new_n776), .B2(new_n841), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n780), .A2(new_n524), .B1(new_n773), .B2(new_n620), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n842), .B(new_n843), .C1(G97), .C2(new_n784), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n839), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G150), .A2(new_n796), .B1(new_n794), .B2(G159), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  INV_X1    g0647(.A(G143), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n847), .B2(new_n790), .C1(new_n848), .C2(new_n788), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n764), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G68), .A2(new_n774), .B1(new_n777), .B2(G132), .ZN(new_n853));
  INV_X1    g0653(.A(G50), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n854), .B2(new_n780), .C1(new_n278), .C2(new_n783), .ZN(new_n855));
  OR3_X1    g0655(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n849), .A2(new_n850), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(KEYINPUT103), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n755), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n838), .B1(new_n859), .B2(new_n861), .C1(new_n822), .C2(new_n757), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n834), .A2(new_n862), .ZN(G384));
  XNOR2_X1  g0663(.A(new_n579), .B(KEYINPUT107), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(new_n867), .A3(G116), .A4(new_n224), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  OAI211_X1 g0669(.A(new_n226), .B(G77), .C1(new_n278), .C2(new_n353), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n854), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n262), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G330), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n377), .B1(new_n374), .B2(KEYINPUT76), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n372), .B1(new_n366), .B2(new_n371), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT108), .B(new_n361), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT109), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n377), .A2(new_n687), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT109), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n378), .A2(KEYINPUT108), .A3(new_n880), .A4(new_n361), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n878), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n735), .A2(KEYINPUT31), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT31), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n643), .B2(new_n688), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n735), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n888), .A3(new_n822), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n424), .B1(new_n428), .B2(new_n435), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n443), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n343), .A3(new_n436), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n685), .B1(new_n895), .B2(new_n447), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n674), .B2(new_n455), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n466), .A2(new_n467), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n896), .B1(new_n900), .B2(new_n458), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n895), .A2(new_n447), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n422), .A3(new_n450), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n899), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n685), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n448), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n463), .A2(new_n899), .A3(new_n451), .A4(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n892), .B1(new_n898), .B2(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n672), .A2(new_n673), .B1(new_n453), .B2(new_n454), .ZN(new_n911));
  OAI221_X1 g0711(.A(KEYINPUT38), .B1(new_n904), .B2(new_n908), .C1(new_n911), .C2(new_n897), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n890), .A2(new_n891), .A3(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n898), .A2(new_n909), .A3(new_n892), .ZN(new_n915));
  INV_X1    g0715(.A(new_n906), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n471), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n451), .A2(new_n906), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT37), .B1(new_n918), .B2(new_n468), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n907), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT40), .B1(new_n889), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n874), .B1(new_n914), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n888), .A2(G330), .A3(new_n472), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n923), .ZN(new_n927));
  INV_X1    g0727(.A(new_n913), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n889), .A2(KEYINPUT40), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n888), .A2(new_n472), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n924), .A2(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n455), .A2(new_n905), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT110), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n910), .B(new_n912), .C1(new_n921), .C2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(KEYINPUT110), .A2(KEYINPUT39), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n936), .A2(KEYINPUT39), .B1(new_n922), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n378), .A2(new_n687), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n934), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n397), .A2(new_n687), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n826), .B2(new_n827), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n882), .A2(new_n883), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n943), .A2(new_n928), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n932), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n678), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n666), .A2(new_n710), .A3(new_n688), .ZN(new_n949));
  INV_X1    g0749(.A(new_n720), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n687), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n949), .B1(new_n952), .B2(new_n710), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n948), .B1(new_n953), .B2(new_n472), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n262), .B2(new_n681), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n947), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n873), .B1(new_n956), .B2(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n765), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n235), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n760), .B1(new_n703), .B2(new_n613), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G283), .A2(new_n794), .B1(new_n796), .B2(G294), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n493), .B2(new_n788), .C1(new_n841), .C2(new_n790), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n773), .A2(new_n482), .ZN(new_n965));
  XNOR2_X1  g0765(.A(KEYINPUT114), .B(G317), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(new_n777), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n780), .A2(new_n487), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(KEYINPUT46), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n524), .B2(new_n783), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n964), .A2(new_n764), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT115), .ZN(new_n973));
  AOI22_X1  g0773(.A1(G150), .A2(new_n789), .B1(new_n796), .B2(G159), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n854), .B2(new_n793), .C1(new_n848), .C2(new_n790), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n783), .A2(new_n353), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n253), .B1(new_n780), .B2(new_n278), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n774), .A2(G77), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n847), .B2(new_n776), .ZN(new_n979));
  NOR4_X1   g0779(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n982), .A2(KEYINPUT47), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n755), .B1(new_n982), .B2(KEYINPUT47), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n752), .B1(new_n960), .B2(new_n962), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n657), .A2(new_n658), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n653), .A2(new_n687), .ZN(new_n987));
  MUX2_X1   g0787(.A(new_n649), .B(new_n986), .S(new_n987), .Z(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n758), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT113), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n700), .A2(new_n693), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n585), .A2(new_n687), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n592), .A2(new_n588), .A3(new_n992), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n991), .A2(KEYINPUT42), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n588), .B1(new_n993), .B2(new_n562), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n688), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT42), .B1(new_n991), .B2(new_n993), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n988), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n1001));
  NAND2_X1  g0801(.A1(new_n988), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT112), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n998), .A2(KEYINPUT112), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n998), .A2(new_n1002), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n661), .A2(new_n687), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n993), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1008), .B1(new_n697), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n697), .A2(new_n1011), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1005), .A2(new_n1013), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT44), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n701), .A2(new_n1016), .A3(new_n1010), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n701), .B2(new_n1010), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n701), .A2(new_n1010), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n1010), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n692), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n991), .B1(new_n696), .B2(new_n700), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n697), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n748), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n704), .B(KEYINPUT41), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n751), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n990), .B1(new_n1015), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1033), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1035), .A2(KEYINPUT113), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n989), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(G387));
  INV_X1    g0838(.A(new_n1030), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n751), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n959), .B1(new_n232), .B2(G45), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n706), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n767), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT50), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n388), .B2(new_n854), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n387), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n706), .B(new_n502), .C1(new_n353), .C2(new_n349), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1043), .A2(new_n1048), .B1(G107), .B2(new_n206), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n812), .B1(new_n1049), .B2(new_n759), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n784), .A2(new_n613), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n788), .B2(new_n854), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT116), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G68), .A2(new_n794), .B1(new_n791), .B2(G159), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n796), .A2(new_n283), .ZN(new_n1055));
  INV_X1    g0855(.A(G150), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n776), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n780), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n965), .C1(G77), .C2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1053), .A2(new_n1060), .A3(new_n852), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G322), .A2(new_n791), .B1(new_n789), .B2(new_n966), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n493), .B2(new_n793), .C1(new_n841), .C2(new_n795), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT48), .ZN(new_n1064));
  INV_X1    g0864(.A(G283), .ZN(new_n1065));
  INV_X1    g0865(.A(G294), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n783), .C1(new_n1066), .C2(new_n780), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G116), .A2(new_n774), .B1(new_n777), .B2(G326), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n852), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1061), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1050), .B1(new_n696), .B2(new_n814), .C1(new_n1073), .C2(new_n770), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1040), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n748), .A2(new_n1039), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n704), .B1(new_n747), .B2(new_n1030), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT117), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT117), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(G393));
  NOR2_X1   g0881(.A1(new_n747), .A2(new_n1030), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n705), .B1(new_n1082), .B2(new_n1025), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1025), .B(new_n697), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n1082), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1011), .A2(new_n758), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n959), .A2(new_n243), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n759), .B1(new_n482), .B2(new_n206), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n752), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1056), .A2(new_n790), .B1(new_n788), .B2(new_n806), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT51), .Z(new_n1091));
  AOI22_X1  g0891(.A1(G50), .A2(new_n796), .B1(new_n794), .B2(new_n388), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n783), .A2(new_n349), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n780), .A2(new_n353), .B1(new_n773), .B2(new_n620), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G143), .C2(new_n777), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n764), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G283), .A2(new_n1058), .B1(new_n777), .B2(G322), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n249), .C1(new_n524), .C2(new_n773), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G116), .B2(new_n784), .ZN(new_n1099));
  INV_X1    g0899(.A(G317), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n841), .A2(new_n788), .B1(new_n790), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT52), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G294), .A2(new_n794), .B1(new_n796), .B2(G303), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1091), .A2(new_n1096), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1089), .B1(new_n1107), .B2(new_n755), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1084), .A2(new_n751), .B1(new_n1086), .B2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1085), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G390));
  INV_X1    g0911(.A(new_n472), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n678), .B(new_n925), .C1(new_n722), .C2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n822), .B(G330), .C1(new_n739), .C2(new_n745), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n944), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n884), .A2(new_n888), .A3(G330), .A4(new_n822), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n826), .A2(new_n827), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n942), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n888), .A2(G330), .A3(new_n822), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n944), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n739), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n745), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1126), .A2(new_n884), .A3(G330), .A4(new_n822), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n688), .B(new_n820), .C1(new_n717), .C2(new_n720), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1119), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1123), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1113), .B1(new_n1121), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n938), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n940), .B1(new_n915), .B2(new_n921), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1129), .B2(new_n884), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1116), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1114), .A2(new_n944), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1140), .B(new_n1137), .C1(new_n1134), .C2(new_n938), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n939), .B1(new_n1120), .B2(new_n884), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n920), .B1(new_n911), .B2(new_n906), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n935), .B1(new_n1144), .B2(new_n892), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT39), .B1(new_n913), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n892), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n912), .A3(new_n937), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1127), .B(new_n1138), .C1(new_n1143), .C2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1137), .B1(new_n1134), .B2(new_n938), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1132), .C1(new_n1151), .C2(new_n1116), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1142), .A2(new_n704), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n752), .B1(new_n836), .B2(new_n283), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n253), .B(new_n1093), .C1(G87), .C2(new_n1058), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n773), .A2(new_n353), .B1(new_n776), .B2(new_n1066), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT118), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(new_n487), .C2(new_n788), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G107), .A2(new_n796), .B1(new_n791), .B2(G283), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n482), .B2(new_n793), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT54), .B(G143), .Z(new_n1161));
  AOI22_X1  g0961(.A1(G132), .A2(new_n789), .B1(new_n794), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n790), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n796), .A2(G137), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT53), .B1(new_n780), .B2(new_n1056), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n780), .A2(KEYINPUT53), .A3(new_n1056), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G159), .B2(new_n784), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n253), .B1(new_n773), .B2(new_n854), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G125), .B2(new_n777), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1158), .A2(new_n1160), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1154), .B1(new_n1172), .B2(new_n755), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1149), .B2(new_n757), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT119), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n751), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1153), .A2(new_n1177), .ZN(G378));
  INV_X1    g0978(.A(new_n924), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n302), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n677), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT55), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n299), .A2(new_n685), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n322), .A2(KEYINPUT55), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1181), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1191), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n1180), .A3(new_n1189), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n941), .A2(new_n1196), .A3(new_n945), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n933), .B1(new_n1149), .B2(new_n939), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1120), .A2(new_n913), .A3(new_n884), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1179), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1196), .B1(new_n941), .B2(new_n945), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1195), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n924), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(new_n751), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n752), .B1(new_n836), .B2(G50), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G128), .A2(new_n789), .B1(new_n796), .B2(G132), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n847), .B2(new_n793), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n784), .A2(G150), .B1(new_n1058), .B2(new_n1161), .ZN(new_n1209));
  INV_X1    g1009(.A(G125), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n790), .ZN(new_n1211));
  OR3_X1    g1011(.A1(new_n1208), .A2(KEYINPUT59), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(KEYINPUT59), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n245), .B(new_n267), .C1(new_n773), .C2(new_n806), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G124), .B2(new_n777), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n764), .A2(G41), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G97), .A2(new_n796), .B1(new_n789), .B2(G107), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G116), .A2(new_n791), .B1(new_n794), .B2(new_n613), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n780), .A2(new_n349), .B1(new_n776), .B2(new_n1065), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n976), .B(new_n1220), .C1(G58), .C2(new_n774), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1217), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n854), .C1(G33), .C2(G41), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1216), .A2(new_n1224), .A3(new_n1225), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1206), .B1(new_n1228), .B2(new_n755), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1196), .B2(new_n757), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1205), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1121), .A2(new_n1131), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1113), .B1(new_n1176), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1201), .A2(KEYINPUT57), .A3(new_n1204), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n704), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1202), .A2(new_n1203), .A3(new_n924), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n924), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1113), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1152), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1231), .B1(new_n1235), .B2(new_n1241), .ZN(G375));
  NAND3_X1  g1042(.A1(new_n1121), .A2(new_n1131), .A3(new_n1113), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1133), .A2(new_n1032), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n764), .B1(new_n278), .B2(new_n773), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT121), .Z(new_n1246));
  AOI22_X1  g1046(.A1(G159), .A2(new_n1058), .B1(new_n777), .B2(G128), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n854), .B2(new_n783), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G150), .B2(new_n794), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n791), .A2(G132), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G137), .A2(new_n789), .B1(new_n796), .B2(new_n1161), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G97), .A2(new_n1058), .B1(new_n777), .B2(G303), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1253), .A2(new_n249), .A3(new_n978), .A4(new_n1051), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G107), .A2(new_n794), .B1(new_n791), .B2(G294), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G116), .A2(new_n796), .B1(new_n789), .B2(G283), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1246), .A2(new_n1252), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT122), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n755), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1258), .A2(KEYINPUT122), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n752), .B1(G68), .B2(new_n836), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n944), .B2(new_n756), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1232), .B2(new_n751), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1244), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(G381));
  OR2_X1    g1066(.A1(G375), .A2(G378), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1079), .A2(new_n1080), .A3(new_n816), .ZN(new_n1268));
  INV_X1    g1068(.A(G384), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1265), .A2(new_n1269), .A3(new_n1110), .ZN(new_n1270));
  OR3_X1    g1070(.A1(G387), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT123), .ZN(G407));
  OAI211_X1 g1073(.A(G407), .B(G213), .C1(G343), .C2(new_n1267), .ZN(G409));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1153), .A2(new_n1177), .A3(new_n1205), .A4(new_n1230), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1238), .A2(new_n1240), .A3(new_n1032), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G378), .B2(G375), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1243), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1121), .A2(new_n1131), .A3(KEYINPUT60), .A4(new_n1113), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(new_n1133), .A3(new_n704), .A4(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(G384), .A3(new_n1264), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1286), .B2(new_n1264), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT124), .B1(new_n1282), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT126), .B1(new_n1282), .B2(new_n1290), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n1275), .A2(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G375), .A2(G378), .ZN(new_n1295));
  AND4_X1   g1095(.A1(new_n1153), .A2(new_n1177), .A3(new_n1205), .A4(new_n1230), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1238), .A2(new_n1240), .A3(new_n1032), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1277), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(new_n1298), .A3(new_n1290), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(KEYINPUT126), .B(KEYINPUT63), .C1(new_n1300), .C2(KEYINPUT124), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G393), .A2(G396), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1268), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT125), .B1(new_n1037), .B2(G390), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1037), .A2(G390), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n989), .B(new_n1110), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n1304), .A2(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G387), .A2(new_n1110), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1037), .A2(G390), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(KEYINPUT125), .A3(new_n1310), .A4(new_n1303), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1277), .A2(G2897), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1286), .A2(new_n1264), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1269), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1287), .A3(new_n1313), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1312), .A2(new_n1320), .A3(KEYINPUT61), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1294), .A2(new_n1301), .A3(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT127), .B1(new_n1320), .B2(KEYINPUT61), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT127), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1324), .B(new_n1325), .C1(new_n1282), .C2(new_n1319), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1282), .A2(new_n1328), .A3(new_n1290), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1323), .A2(new_n1326), .A3(new_n1327), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1312), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1322), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1267), .A2(new_n1295), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1333), .B(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1290), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1312), .A2(new_n1334), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1267), .B2(new_n1295), .ZN(new_n1338));
  OAI22_X1  g1138(.A1(new_n1337), .A2(new_n1338), .B1(new_n1289), .B2(new_n1288), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(G402));
endmodule


