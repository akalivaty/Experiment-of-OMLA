//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT69), .B1(new_n203), .B2(G183gat), .ZN(new_n204));
  NOR3_X1   g003(.A1(new_n204), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT67), .B(G183gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n206), .C1(new_n203), .C2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n211), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n213), .A2(KEYINPUT70), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT26), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n214), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(KEYINPUT26), .B2(new_n218), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n215), .B1(new_n214), .B2(new_n220), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n208), .B(new_n212), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT65), .B1(new_n229), .B2(KEYINPUT23), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  NAND3_X1  g031(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n235), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n210), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT64), .A4(new_n233), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n229), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n231), .A2(new_n236), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  OAI211_X1 g044(.A(G183gat), .B(G190gat), .C1(new_n245), .C2(KEYINPUT24), .ZN(new_n246));
  NAND2_X1  g045(.A1(G183gat), .A2(G190gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(KEYINPUT66), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n238), .A2(KEYINPUT67), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G183gat), .ZN(new_n253));
  AOI21_X1  g052(.A(G190gat), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n256), .A2(new_n226), .A3(KEYINPUT25), .A4(new_n227), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT68), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n249), .B(new_n246), .C1(new_n207), .C2(G190gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n224), .B1(new_n244), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G113gat), .ZN(new_n266));
  INV_X1    g065(.A(G113gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G120gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n269), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G127gat), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G134gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n270), .ZN(new_n279));
  XNOR2_X1  g078(.A(G113gat), .B(G120gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(KEYINPUT1), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n273), .A2(new_n281), .A3(KEYINPUT73), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT73), .B1(new_n273), .B2(new_n281), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n242), .A2(new_n243), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(new_n258), .A3(new_n262), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n284), .A3(new_n224), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G227gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n202), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g094(.A(KEYINPUT34), .B(new_n293), .C1(new_n286), .C2(new_n289), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G15gat), .B(G43gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n293), .A3(new_n289), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT33), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n302), .A2(new_n305), .A3(KEYINPUT32), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(new_n302), .B2(KEYINPUT32), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT75), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n310), .B(new_n304), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n286), .A2(new_n293), .A3(new_n289), .ZN(new_n314));
  AOI211_X1 g113(.A(new_n313), .B(new_n314), .C1(KEYINPUT33), .C2(new_n300), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n297), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n297), .ZN(new_n318));
  AOI211_X1 g117(.A(new_n315), .B(new_n318), .C1(new_n309), .C2(new_n311), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G148gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT80), .B(G148gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  AND2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327));
  NOR2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G148gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G141gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n327), .ZN(new_n335));
  XNOR2_X1  g134(.A(G155gat), .B(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n273), .A2(new_n281), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n325), .A2(new_n330), .B1(new_n335), .B2(new_n337), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n273), .A3(new_n281), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n321), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n342), .B1(new_n282), .B2(new_n283), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n339), .A2(new_n340), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(G148gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n354));
  OAI21_X1  g153(.A(G141gat), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n329), .B1(new_n355), .B2(new_n323), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n336), .B1(new_n334), .B2(new_n327), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n331), .A2(new_n359), .A3(new_n338), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n360), .A3(new_n340), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n351), .B1(new_n361), .B2(KEYINPUT4), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n347), .B1(new_n350), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n349), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n351), .A2(KEYINPUT4), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n346), .A2(KEYINPUT5), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n369), .A2(new_n361), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n363), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT6), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n363), .A2(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(new_n368), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n363), .A2(KEYINPUT82), .A3(new_n368), .A4(new_n372), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT31), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(G50gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT76), .B(G197gat), .ZN(new_n387));
  INV_X1    g186(.A(G204gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(G211gat), .B(G218gat), .Z(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT77), .B(G211gat), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT22), .B1(new_n391), .B2(G218gat), .ZN(new_n392));
  OR3_X1    g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n389), .B2(new_n392), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n360), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(KEYINPUT29), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n394), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT29), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(KEYINPUT83), .A3(new_n394), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT3), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n398), .B(new_n399), .C1(new_n404), .C2(new_n342), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n359), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n339), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n399), .B1(new_n410), .B2(new_n398), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n406), .A2(new_n411), .A3(G22gat), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n398), .ZN(new_n414));
  INV_X1    g213(.A(new_n399), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n416), .B2(new_n405), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n386), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n405), .A3(new_n413), .ZN(new_n419));
  OAI21_X1  g218(.A(G22gat), .B1(new_n406), .B2(new_n411), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n385), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G226gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(new_n292), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(KEYINPUT29), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n264), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n264), .A2(KEYINPUT78), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT78), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n288), .A2(new_n429), .A3(new_n224), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n431), .B2(new_n425), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n396), .ZN(new_n433));
  XNOR2_X1  g232(.A(G8gat), .B(G36gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n428), .A2(new_n430), .A3(new_n426), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n288), .A2(new_n425), .A3(new_n224), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n395), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT30), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n433), .A2(new_n441), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n436), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n320), .A2(new_n382), .A3(new_n423), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n363), .A2(KEYINPUT86), .A3(new_n372), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT86), .B1(new_n363), .B2(new_n372), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(new_n368), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n373), .A2(new_n374), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n379), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT87), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n456), .A2(new_n368), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n454), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n379), .A4(new_n375), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n461), .A2(new_n465), .A3(new_n381), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n466), .A2(new_n450), .A3(KEYINPUT35), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n317), .A2(new_n319), .A3(new_n422), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT40), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n370), .A2(new_n361), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n345), .B1(new_n472), .B2(new_n369), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n377), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n476), .B2(KEYINPUT85), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(KEYINPUT85), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n471), .B1(new_n463), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n471), .B2(new_n479), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n422), .B1(new_n481), .B2(new_n450), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n433), .A2(new_n484), .A3(new_n441), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n436), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n433), .B2(new_n441), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT38), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT92), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(KEYINPUT38), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n485), .A2(new_n493), .A3(new_n436), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n432), .B2(new_n396), .ZN(new_n497));
  INV_X1    g296(.A(new_n425), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n428), .B2(new_n430), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT88), .B(new_n395), .C1(new_n499), .C2(new_n427), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n438), .A2(new_n396), .A3(new_n439), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n438), .A2(KEYINPUT89), .A3(new_n396), .A4(new_n439), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n497), .A2(new_n500), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n505), .A2(KEYINPUT90), .A3(KEYINPUT37), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT90), .B1(new_n505), .B2(KEYINPUT37), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n495), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n381), .A2(new_n461), .A3(new_n465), .A4(new_n442), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n492), .B1(new_n510), .B2(KEYINPUT91), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n483), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n419), .A2(new_n420), .A3(new_n385), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n385), .B1(new_n419), .B2(new_n420), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n418), .A2(KEYINPUT84), .A3(new_n421), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n445), .A2(new_n382), .A3(new_n447), .A4(new_n449), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n317), .A2(new_n319), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT74), .B1(new_n314), .B2(new_n313), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n302), .A2(new_n305), .A3(KEYINPUT32), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n310), .B1(new_n527), .B2(new_n304), .ZN(new_n528));
  INV_X1    g327(.A(new_n311), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n316), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n318), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n312), .A2(new_n316), .A3(new_n297), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT36), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n522), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n470), .B1(new_n514), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n382), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(G1gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT16), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n540), .B2(G1gat), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n537), .A3(new_n541), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT99), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT99), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G43gat), .B(G50gat), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT15), .B1(new_n550), .B2(KEYINPUT95), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(KEYINPUT95), .B2(new_n550), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n553));
  INV_X1    g352(.A(G29gat), .ZN(new_n554));
  INV_X1    g353(.A(G36gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI221_X1 g357(.A(new_n558), .B1(new_n554), .B2(new_n555), .C1(KEYINPUT15), .C2(new_n550), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(KEYINPUT96), .A3(new_n557), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n562), .B(new_n563), .C1(new_n554), .C2(new_n555), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n552), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT97), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n560), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n549), .B1(KEYINPUT17), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(new_n560), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT98), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT98), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n569), .A2(new_n576), .A3(KEYINPUT17), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n570), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n545), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n573), .A2(KEYINPUT98), .A3(new_n574), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n576), .B1(new_n569), .B2(KEYINPUT17), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n581), .B1(new_n588), .B2(new_n570), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(KEYINPUT18), .A3(new_n579), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n569), .B(new_n580), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n579), .B(KEYINPUT13), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n585), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n595));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT12), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n594), .A2(KEYINPUT94), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n594), .B2(KEYINPUT94), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(G71gat), .A2(G78gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  XOR2_X1   g407(.A(G57gat), .B(G64gat), .Z(new_n609));
  AOI211_X1 g408(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(KEYINPUT9), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n607), .B1(KEYINPUT9), .B2(new_n608), .ZN(new_n611));
  INV_X1    g410(.A(G64gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(G57gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT100), .B(G57gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(G64gat), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n611), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n545), .B1(KEYINPUT21), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT102), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n622));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT101), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n238), .ZN(new_n627));
  INV_X1    g426(.A(G211gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n624), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n621), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G99gat), .B(G106gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(KEYINPUT105), .A2(KEYINPUT7), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(G85gat), .A3(G92gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT106), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT7), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n639), .A2(new_n644), .A3(G85gat), .A4(G92gat), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G99gat), .A2(G106gat), .ZN(new_n647));
  INV_X1    g446(.A(G85gat), .ZN(new_n648));
  INV_X1    g447(.A(G92gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(KEYINPUT8), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n641), .A2(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n638), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n654), .A2(new_n637), .A3(new_n646), .A4(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n617), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n653), .A2(new_n655), .A3(new_n617), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n656), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n636), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n658), .A2(new_n660), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n636), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n664), .A2(KEYINPUT108), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n676), .B(new_n636), .C1(new_n661), .C2(new_n663), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n675), .A2(new_n677), .A3(new_n669), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n674), .B1(new_n678), .B2(new_n672), .ZN(new_n679));
  OAI221_X1 g478(.A(new_n656), .B1(new_n574), .B2(new_n573), .C1(new_n575), .C2(new_n577), .ZN(new_n680));
  NAND2_X1  g479(.A1(G232gat), .A2(G233gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n573), .A2(new_n662), .B1(KEYINPUT41), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(G190gat), .B(G218gat), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n683), .A2(KEYINPUT41), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G162gat), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT104), .B(G134gat), .Z(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n686), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n680), .A2(new_n692), .A3(new_n684), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n687), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n680), .A2(new_n692), .A3(new_n684), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n680), .B2(new_n684), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n634), .A2(new_n679), .A3(new_n694), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n606), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n535), .A2(new_n536), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g501(.A1(new_n535), .A2(new_n450), .A3(new_n700), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT110), .B(KEYINPUT16), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(new_n537), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT109), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n706), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n703), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT42), .B2(new_n706), .ZN(G1325gat));
  INV_X1    g507(.A(G15gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n535), .A2(new_n700), .ZN(new_n710));
  INV_X1    g509(.A(new_n320), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n524), .A2(new_n533), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G15gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT111), .Z(G1326gat));
  NAND3_X1  g515(.A1(new_n535), .A2(new_n520), .A3(new_n700), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT43), .B(G22gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  NAND2_X1  g518(.A1(new_n698), .A2(new_n694), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n505), .A2(KEYINPUT37), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT90), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n505), .A2(KEYINPUT90), .A3(KEYINPUT37), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n494), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n461), .A2(new_n465), .A3(new_n381), .A4(new_n442), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT91), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n492), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n513), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n534), .B1(new_n729), .B2(new_n482), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n452), .A2(KEYINPUT35), .B1(new_n468), .B2(new_n467), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n720), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n678), .A2(new_n672), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n666), .B2(new_n673), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n606), .A2(new_n634), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n382), .A2(G29gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n737), .A2(KEYINPUT112), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT112), .B1(new_n737), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n679), .B(KEYINPUT113), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n605), .A3(new_n633), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n748), .B(new_n720), .C1(new_n730), .C2(new_n731), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G29gat), .B1(new_n751), .B2(new_n382), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n740), .A2(KEYINPUT45), .A3(new_n741), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n744), .A2(new_n752), .A3(new_n753), .ZN(G1328gat));
  NOR3_X1   g553(.A1(new_n737), .A2(G36gat), .A3(new_n451), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT46), .ZN(new_n756));
  OAI21_X1  g555(.A(G36gat), .B1(new_n751), .B2(new_n451), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759));
  INV_X1    g558(.A(new_n713), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n760), .B(new_n746), .C1(new_n747), .C2(new_n749), .ZN(new_n761));
  INV_X1    g560(.A(G43gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n733), .A2(new_n762), .A3(new_n320), .A4(new_n736), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI221_X1 g566(.A(new_n764), .B1(new_n759), .B2(KEYINPUT47), .C1(new_n761), .C2(new_n762), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1330gat));
  INV_X1    g568(.A(new_n520), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n737), .A2(G50gat), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n520), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G50gat), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(G50gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n750), .B2(new_n422), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n773), .A2(KEYINPUT48), .B1(new_n775), .B2(new_n777), .ZN(G1331gat));
  NOR3_X1   g577(.A1(new_n745), .A2(new_n633), .A3(new_n720), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n535), .A2(new_n606), .A3(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n382), .B(KEYINPUT115), .Z(new_n781));
  OR2_X1    g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(new_n614), .Z(G1332gat));
  OR2_X1    g582(.A1(new_n780), .A2(new_n451), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT49), .B(G64gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1333gat));
  INV_X1    g586(.A(G71gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n780), .B2(new_n711), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n713), .A2(G71gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n780), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT50), .ZN(G1334gat));
  OR2_X1    g591(.A1(new_n780), .A2(new_n770), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g593(.A1(new_n605), .A2(new_n634), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n735), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n747), .B2(new_n749), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G85gat), .B1(new_n798), .B2(new_n382), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n720), .B(new_n795), .C1(new_n730), .C2(new_n731), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n535), .A2(KEYINPUT51), .A3(new_n720), .A4(new_n795), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n735), .A2(new_n648), .A3(new_n536), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n799), .B1(new_n805), .B2(new_n806), .ZN(G1336gat));
  AOI21_X1  g606(.A(new_n649), .B1(new_n797), .B2(new_n450), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  INV_X1    g610(.A(new_n745), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n804), .A2(new_n649), .A3(new_n450), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n649), .A3(new_n450), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n810), .B1(new_n805), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n816), .B2(new_n808), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(G1337gat));
  OAI21_X1  g617(.A(G99gat), .B1(new_n798), .B2(new_n760), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n711), .A2(G99gat), .A3(new_n679), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n805), .B2(new_n820), .ZN(G1338gat));
  NOR2_X1   g620(.A1(new_n423), .A2(G106gat), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n812), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT117), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n805), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(G106gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n797), .B2(new_n520), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT53), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n796), .ZN(new_n829));
  INV_X1    g628(.A(new_n749), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n748), .B1(new_n535), .B2(new_n720), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n422), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  INV_X1    g633(.A(new_n823), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n804), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n834), .B1(new_n833), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n828), .B1(new_n837), .B2(new_n838), .ZN(G1339gat));
  NAND4_X1  g638(.A1(new_n585), .A2(new_n590), .A3(new_n593), .A4(new_n601), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n589), .A2(new_n579), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n591), .A2(new_n592), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n599), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(KEYINPUT121), .A3(new_n843), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n675), .B2(new_n677), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n661), .A2(new_n636), .A3(new_n663), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT119), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n661), .A2(new_n663), .A3(new_n852), .A4(new_n636), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n849), .B(new_n672), .C1(new_n666), .C2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n674), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n846), .A2(new_n847), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n720), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n594), .A2(KEYINPUT94), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n600), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n858), .A3(new_n602), .A4(new_n857), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n840), .A2(new_n843), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n720), .B1(new_n864), .B2(new_n735), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n860), .A2(new_n866), .A3(new_n633), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n605), .A2(new_n699), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n320), .A3(new_n770), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n451), .A2(new_n536), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G113gat), .B1(new_n874), .B2(new_n606), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n634), .B1(new_n863), .B2(new_n865), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n868), .B1(new_n876), .B2(new_n860), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(new_n450), .A3(new_n781), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n468), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n267), .A3(new_n605), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n875), .A2(new_n880), .ZN(G1340gat));
  OAI21_X1  g680(.A(G120gat), .B1(new_n874), .B2(new_n745), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n265), .A3(new_n735), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1341gat));
  AOI21_X1  g683(.A(G127gat), .B1(new_n879), .B2(new_n634), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n633), .A2(new_n276), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n873), .B2(new_n886), .ZN(G1342gat));
  NAND3_X1  g686(.A1(new_n879), .A2(new_n274), .A3(new_n720), .ZN(new_n888));
  XNOR2_X1  g687(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  INV_X1    g690(.A(new_n720), .ZN(new_n892));
  OAI21_X1  g691(.A(G134gat), .B1(new_n874), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(G1343gat));
  NAND2_X1  g693(.A1(new_n870), .A2(new_n520), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT57), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n870), .A2(new_n897), .A3(new_n422), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n713), .A2(new_n872), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G141gat), .B1(new_n900), .B2(new_n606), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n878), .A2(new_n422), .A3(new_n760), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n322), .A3(new_n605), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g704(.A(new_n324), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n906), .A3(new_n735), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n713), .A2(new_n679), .A3(new_n872), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n895), .B2(new_n897), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n910), .B(new_n897), .C1(new_n877), .C2(new_n770), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n870), .A2(KEYINPUT57), .A3(new_n422), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n909), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n332), .B1(new_n915), .B2(KEYINPUT124), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n917), .B(new_n909), .C1(new_n911), .C2(new_n914), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n908), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n900), .ZN(new_n920));
  AOI211_X1 g719(.A(KEYINPUT59), .B(new_n906), .C1(new_n920), .C2(new_n735), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n907), .B1(new_n919), .B2(new_n921), .ZN(G1345gat));
  AOI21_X1  g721(.A(G155gat), .B1(new_n902), .B2(new_n634), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n634), .A2(G155gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n920), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n900), .B2(new_n892), .ZN(new_n926));
  INV_X1    g725(.A(G162gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n902), .A2(new_n927), .A3(new_n720), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n877), .A2(new_n536), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(new_n450), .A3(new_n468), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n216), .A3(new_n605), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n781), .A2(new_n450), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT125), .Z(new_n934));
  NOR3_X1   g733(.A1(new_n871), .A2(new_n606), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n216), .B2(new_n935), .ZN(G1348gat));
  AOI21_X1  g735(.A(G176gat), .B1(new_n931), .B2(new_n735), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n871), .A2(new_n934), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n745), .A2(new_n217), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G1349gat));
  NAND3_X1  g739(.A1(new_n931), .A2(new_n209), .A3(new_n634), .ZN(new_n941));
  INV_X1    g740(.A(new_n207), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n871), .A2(new_n633), .A3(new_n934), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n931), .A2(new_n210), .A3(new_n720), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n938), .A2(new_n720), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(G190gat), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT61), .B(new_n210), .C1(new_n938), .C2(new_n720), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT126), .B(new_n946), .C1(new_n949), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  OR3_X1    g754(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT127), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n934), .A2(new_n713), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT127), .B1(new_n911), .B2(new_n914), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n956), .A2(new_n605), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G197gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n713), .A2(new_n423), .A3(new_n451), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n930), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OR3_X1    g762(.A1(new_n963), .A2(G197gat), .A3(new_n606), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n964), .ZN(G1352gat));
  NAND4_X1  g764(.A1(new_n956), .A2(new_n812), .A3(new_n957), .A4(new_n958), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n962), .A2(new_n388), .A3(new_n735), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT62), .Z(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1353gat));
  OR3_X1    g769(.A1(new_n963), .A2(new_n391), .A3(new_n633), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n911), .A2(new_n914), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n934), .A2(new_n713), .A3(new_n633), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n976));
  AOI211_X1 g775(.A(new_n976), .B(new_n628), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n971), .B1(new_n975), .B2(new_n977), .ZN(G1354gat));
  INV_X1    g777(.A(G218gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n892), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n963), .B2(new_n892), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


