//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G101), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n196), .A2(new_n199), .A3(new_n203), .A4(new_n200), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n206), .A3(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT0), .A3(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n198), .A2(G104), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n195), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n204), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(new_n224), .A3(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(G128), .B1(new_n210), .B2(new_n212), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n224), .A2(new_n209), .A3(G143), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n208), .A2(new_n219), .B1(new_n229), .B2(KEYINPUT10), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT10), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n226), .B2(new_n227), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n209), .A2(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n236), .B(KEYINPUT66), .C1(new_n217), .C2(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n232), .B1(new_n238), .B2(new_n225), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n204), .A2(new_n222), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n204), .B2(new_n222), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n239), .A2(KEYINPUT76), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT76), .B1(new_n239), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n231), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT78), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G134), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G137), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT64), .B(KEYINPUT11), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n252), .B(new_n254), .C1(new_n255), .C2(new_n249), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n253), .A2(G137), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n250), .A2(KEYINPUT11), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n250), .A2(KEYINPUT11), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n248), .A2(G134), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n249), .B2(new_n251), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n258), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT78), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n231), .B(new_n268), .C1(new_n244), .C2(new_n245), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n247), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n231), .B(new_n266), .C1(new_n244), .C2(new_n245), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n194), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n213), .A2(KEYINPUT1), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(new_n234), .B2(new_n237), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n223), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT77), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n228), .A2(new_n225), .ZN(new_n278));
  INV_X1    g092(.A(new_n223), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n275), .A2(new_n277), .A3(new_n223), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n267), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n281), .A2(KEYINPUT12), .A3(new_n267), .A4(new_n282), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n271), .A2(new_n194), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n187), .B(new_n188), .C1(new_n272), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n194), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n211), .A2(G146), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n273), .B1(new_n292), .B2(new_n235), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT66), .B1(new_n293), .B2(new_n236), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n226), .A2(new_n233), .A3(new_n227), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n225), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n243), .A2(new_n296), .A3(KEYINPUT10), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n239), .A2(KEYINPUT76), .A3(new_n243), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n230), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n291), .B1(new_n301), .B2(new_n266), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n267), .B1(new_n301), .B2(new_n268), .ZN(new_n303));
  INV_X1    g117(.A(new_n269), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n271), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n291), .B1(new_n287), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n307), .A3(G469), .ZN(new_n308));
  NAND2_X1  g122(.A1(G469), .A2(G902), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n290), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(KEYINPUT67), .A2(G116), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT67), .A2(G116), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(G119), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G116), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(G119), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT2), .B(G113), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n321), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n316), .A3(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n262), .A2(new_n264), .A3(new_n258), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n254), .A2(KEYINPUT65), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n253), .A3(G137), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n330), .A3(new_n249), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G131), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n296), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n219), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n257), .B2(new_n265), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n332), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n275), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n256), .A2(G131), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n219), .B1(new_n339), .B2(new_n327), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n338), .A2(KEYINPUT30), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n325), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G237), .A2(G953), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G210), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT27), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G101), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n325), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n333), .A2(new_n335), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n342), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT31), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT30), .B1(new_n338), .B2(new_n340), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n335), .B(new_n326), .C1(new_n275), .C2(new_n337), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n338), .A2(new_n340), .A3(new_n325), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT31), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n347), .ZN(new_n358));
  INV_X1    g172(.A(new_n347), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n335), .B1(new_n275), .B2(new_n337), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT68), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n325), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n335), .B(KEYINPUT68), .C1(new_n275), .C2(new_n337), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT28), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n325), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(new_n349), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n359), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n351), .A2(new_n358), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G472), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n188), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT32), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n369), .A2(new_n373), .A3(new_n370), .A4(new_n188), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n361), .B1(new_n338), .B2(new_n340), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n363), .A3(new_n348), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n365), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n348), .B1(new_n333), .B2(new_n335), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT28), .B1(new_n379), .B2(new_n355), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n380), .A3(new_n347), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G902), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n381), .B(new_n382), .C1(new_n347), .C2(new_n356), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n370), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n375), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(G234), .A2(G237), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(G952), .A3(new_n190), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(G902), .A3(G953), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT21), .B(G898), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G214), .B1(G237), .B2(G902), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n325), .A2(new_n207), .A3(new_n205), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n223), .A2(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n316), .A2(KEYINPUT5), .A3(new_n319), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n318), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(G113), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n204), .A2(new_n222), .A3(new_n240), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n405), .A3(new_n324), .A4(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G122), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n400), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT6), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n400), .A2(new_n407), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n416));
  INV_X1    g230(.A(G125), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n275), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n219), .A2(G125), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(G224), .A3(new_n190), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n190), .A2(G224), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n415), .A2(new_n416), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT80), .A2(KEYINPUT7), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(new_n419), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n405), .A2(new_n324), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n279), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n405), .A2(new_n324), .A3(new_n223), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n408), .B(KEYINPUT8), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n427), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n418), .A2(new_n419), .A3(new_n434), .A4(new_n425), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n428), .A2(new_n409), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n188), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n399), .B1(new_n424), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G210), .B1(G237), .B2(G902), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n421), .A2(new_n423), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n409), .A2(KEYINPUT6), .B1(new_n411), .B2(new_n413), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n188), .A4(new_n436), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n440), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n444), .A2(new_n188), .A3(new_n436), .A4(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n398), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n417), .A2(G140), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT16), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n454));
  INV_X1    g268(.A(G140), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(G125), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n417), .A2(KEYINPUT71), .A3(G140), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n450), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n453), .B1(new_n458), .B2(new_n452), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G146), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n343), .A2(G143), .A3(G214), .ZN(new_n461));
  AOI21_X1  g275(.A(G143), .B1(new_n343), .B2(G214), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n464));
  INV_X1    g278(.A(G237), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n190), .A3(G214), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n211), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n343), .A2(G143), .A3(G214), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n258), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n209), .B(new_n453), .C1(new_n458), .C2(new_n452), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT17), .B(G131), .C1(new_n461), .C2(new_n462), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n460), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n417), .A2(G140), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n451), .A2(new_n474), .A3(new_n209), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n458), .B2(new_n209), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n467), .A2(KEYINPUT83), .A3(new_n468), .ZN(new_n477));
  NAND2_X1  g291(.A1(KEYINPUT18), .A2(G131), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G113), .B(G122), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n195), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n477), .B(new_n478), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n486), .B2(new_n476), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n463), .A2(new_n469), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT19), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n451), .A2(new_n474), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n458), .B2(new_n489), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n460), .B(new_n488), .C1(G146), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n485), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT84), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n482), .A2(new_n484), .B1(new_n487), .B2(new_n492), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n494), .A4(new_n495), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n485), .A2(new_n493), .A3(new_n495), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT20), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n484), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n482), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n482), .A2(new_n505), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n188), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G475), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n503), .A2(KEYINPUT86), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT86), .B1(new_n503), .B2(new_n509), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G217), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n311), .A2(new_n513), .A3(G953), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n273), .A2(G143), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n253), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G128), .B(G143), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT87), .B1(new_n317), .B2(G122), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n522));
  INV_X1    g336(.A(G122), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(G116), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n314), .A2(G122), .A3(new_n315), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n198), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n198), .B1(new_n525), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n520), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n519), .A2(G134), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n519), .A2(G134), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n314), .A2(new_n534), .A3(G122), .A4(new_n315), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n535), .A2(new_n525), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n198), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n530), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n515), .B1(new_n539), .B2(KEYINPUT88), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n538), .A2(new_n533), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n530), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(KEYINPUT88), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n541), .A3(new_n530), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n515), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n547), .A3(new_n188), .ZN(new_n548));
  INV_X1    g362(.A(G478), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n548), .B(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n449), .A2(new_n512), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n513), .B1(G234), .B2(new_n188), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT72), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n560));
  INV_X1    g374(.A(G119), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(G128), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT23), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT23), .B1(new_n273), .B2(G119), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT70), .B1(new_n273), .B2(G119), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G110), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT69), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n273), .B2(G119), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(KEYINPUT69), .A3(G128), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n571), .A2(new_n572), .B1(G119), .B2(new_n273), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT24), .B(G110), .Z(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n460), .B2(new_n471), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n568), .A2(G110), .B1(new_n573), .B2(new_n574), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n460), .A2(new_n578), .A3(new_n475), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n559), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n460), .A2(new_n471), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n460), .A2(new_n578), .A3(new_n475), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n558), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n585), .A3(new_n188), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT25), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n554), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n585), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n554), .A2(G902), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n313), .A2(new_n388), .A3(new_n553), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n540), .A2(new_n543), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n539), .A2(KEYINPUT88), .A3(new_n514), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n514), .A2(KEYINPUT90), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n539), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT33), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n549), .A2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n548), .A2(new_n549), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n511), .B2(new_n510), .ZN(new_n611));
  INV_X1    g425(.A(new_n397), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n440), .B1(new_n424), .B2(new_n437), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n448), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n396), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT89), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n370), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n369), .A2(new_n188), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n619), .B1(new_n369), .B2(new_n188), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n621), .A2(new_n622), .A3(new_n595), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n313), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NAND2_X1  g440(.A1(new_n502), .A2(new_n496), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n627), .A2(new_n509), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n615), .A2(new_n552), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n313), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  OAI21_X1  g447(.A(KEYINPUT91), .B1(new_n577), .B2(new_n579), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT91), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n583), .A2(new_n635), .A3(new_n584), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n634), .B2(new_n636), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n593), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT92), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(KEYINPUT92), .B(new_n593), .C1(new_n638), .C2(new_n639), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n590), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT93), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n357), .B1(new_n356), .B2(new_n347), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n347), .B1(new_n378), .B2(new_n380), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n354), .A2(KEYINPUT31), .A3(new_n359), .A4(new_n355), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n618), .B1(new_n649), .B2(G902), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT93), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n590), .A2(new_n642), .A3(new_n651), .A4(new_n643), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n620), .A2(new_n645), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n313), .A2(new_n653), .A3(new_n553), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND2_X1  g470(.A1(new_n645), .A2(new_n652), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n375), .B2(new_n387), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n313), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n548), .B(new_n550), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT94), .B(G900), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n390), .B1(new_n661), .B2(new_n392), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n628), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n613), .A2(new_n448), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n397), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT95), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT95), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n663), .B2(new_n665), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n659), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XNOR2_X1  g486(.A(new_n662), .B(KEYINPUT39), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n313), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n366), .A2(new_n349), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT96), .B1(new_n676), .B2(new_n359), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n676), .A2(KEYINPUT96), .A3(new_n359), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n677), .B(new_n678), .C1(new_n347), .C2(new_n356), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n679), .B2(G902), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n375), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT97), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n446), .A2(new_n448), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT38), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n660), .B1(new_n510), .B2(new_n511), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n686), .A2(new_n612), .A3(new_n644), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT98), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n675), .A2(new_n682), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n211), .ZN(G45));
  NAND2_X1  g507(.A1(new_n503), .A2(new_n509), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT86), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n503), .A2(KEYINPUT86), .A3(new_n509), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n610), .A3(new_n662), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n665), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n659), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  OAI21_X1  g516(.A(new_n271), .B1(new_n303), .B2(new_n304), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n289), .B1(new_n703), .B2(new_n291), .ZN(new_n704));
  OAI21_X1  g518(.A(G469), .B1(new_n704), .B2(G902), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n705), .A2(new_n312), .A3(new_n290), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n388), .A2(new_n596), .A3(new_n706), .A4(new_n616), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n388), .A2(new_n596), .A3(new_n706), .A4(new_n630), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NAND4_X1  g525(.A1(new_n705), .A2(new_n312), .A3(new_n290), .A4(new_n614), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT99), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n696), .A2(new_n697), .A3(new_n552), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n395), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n658), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT100), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n386), .B1(new_n372), .B2(new_n374), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n718), .A2(new_n657), .A3(new_n714), .A4(new_n395), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT99), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n712), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n712), .A2(new_n721), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n719), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n717), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OAI21_X1  g540(.A(G472), .B1(new_n649), .B2(G902), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n371), .A2(new_n727), .A3(new_n596), .A4(new_n396), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n698), .A2(KEYINPUT101), .A3(new_n660), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n665), .B1(new_n686), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(new_n706), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n371), .A3(new_n644), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n699), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n722), .B2(new_n723), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  AND2_X1   g551(.A1(new_n448), .A2(new_n397), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n446), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n446), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n312), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n308), .A2(KEYINPUT102), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT102), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n305), .A2(new_n307), .A3(new_n745), .A4(G469), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n290), .A2(new_n744), .A3(new_n309), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT104), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n742), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n741), .B1(new_n446), .B2(new_n738), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n290), .A2(new_n744), .A3(new_n309), .A4(new_n746), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n752), .A3(new_n312), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n388), .A2(new_n596), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n699), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n756), .B1(new_n748), .B2(new_n754), .ZN(new_n763));
  OR2_X1    g577(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n758), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  XOR2_X1   g581(.A(new_n663), .B(KEYINPUT106), .Z(new_n768));
  NAND2_X1  g582(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(new_n312), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n305), .A2(new_n307), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT45), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(G469), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n775), .B2(new_n309), .ZN(new_n776));
  INV_X1    g590(.A(new_n290), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n309), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n771), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n673), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n751), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n512), .A2(new_n610), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(KEYINPUT43), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n789), .B(new_n644), .C1(new_n621), .C2(new_n622), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n782), .B(new_n792), .C1(new_n791), .C2(new_n790), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  XNOR2_X1  g608(.A(new_n780), .B(KEYINPUT47), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n783), .A2(new_n388), .A3(new_n596), .A4(new_n699), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  AND2_X1   g612(.A1(new_n789), .A2(new_n391), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n727), .A2(new_n371), .A3(new_n596), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n706), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n801), .A2(new_n397), .A3(new_n685), .A4(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT50), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT50), .ZN(new_n805));
  INV_X1    g619(.A(new_n734), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n802), .A2(new_n783), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n801), .A2(new_n783), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n705), .A2(new_n290), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT109), .Z(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n312), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n810), .B1(new_n795), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n682), .A2(new_n596), .A3(new_n391), .A4(new_n807), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT116), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n606), .A2(new_n607), .B1(new_n549), .B2(new_n548), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n512), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n809), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  OAI211_X1 g636(.A(G952), .B(new_n190), .C1(new_n801), .C2(new_n713), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n808), .A2(new_n757), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT48), .Z(new_n825));
  INV_X1    g639(.A(new_n611), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n823), .B(new_n825), .C1(new_n826), .C2(new_n816), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n597), .A2(new_n707), .A3(new_n710), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n817), .B1(new_n510), .B2(new_n511), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n830), .A2(new_n714), .A3(new_n449), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n312), .A3(new_n310), .A4(new_n623), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n654), .A2(new_n732), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n552), .A2(new_n628), .A3(new_n662), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT110), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n783), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n755), .A2(new_n735), .B1(new_n659), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n725), .A2(new_n834), .A3(new_n838), .A4(new_n769), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n763), .A2(new_n758), .A3(new_n764), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n760), .B1(new_n763), .B2(new_n758), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n658), .B(new_n313), .C1(new_n670), .C2(new_n700), .ZN(new_n845));
  INV_X1    g659(.A(new_n644), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n312), .A3(new_n662), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n375), .B2(new_n680), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n729), .A3(new_n731), .A4(new_n753), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n736), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n736), .A2(new_n845), .A3(KEYINPUT52), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n850), .A2(new_n855), .A3(KEYINPUT52), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n844), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n725), .A2(new_n834), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n838), .A2(new_n769), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n864), .A4(new_n766), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n858), .B1(new_n854), .B2(new_n856), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT115), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n854), .A2(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n725), .A2(new_n834), .A3(new_n769), .A4(new_n838), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n852), .A2(KEYINPUT113), .A3(new_n853), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n871), .A2(new_n872), .A3(new_n766), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n843), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n874), .B2(new_n843), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n868), .B(new_n869), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n874), .A2(new_n843), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n766), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n866), .B1(new_n880), .B2(KEYINPUT111), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(KEYINPUT111), .B2(new_n880), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n882), .B2(new_n843), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n878), .B1(new_n883), .B2(new_n869), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n828), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n682), .A2(new_n684), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n784), .A2(new_n595), .A3(new_n771), .A4(new_n612), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT108), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n812), .B2(KEYINPUT49), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(KEYINPUT49), .B2(new_n812), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n885), .B1(new_n886), .B2(new_n890), .ZN(G75));
  NAND2_X1  g705(.A1(new_n415), .A2(new_n416), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n441), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n874), .A2(new_n843), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT114), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n874), .A2(new_n875), .A3(new_n843), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n898), .A2(new_n899), .B1(new_n867), .B2(new_n862), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n896), .B1(new_n900), .B2(new_n188), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n868), .B1(new_n876), .B2(new_n877), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(KEYINPUT117), .A3(G902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n895), .B1(new_n904), .B2(new_n447), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n190), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n900), .A2(new_n188), .A3(new_n447), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n894), .B1(new_n908), .B2(KEYINPUT56), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(G51));
  INV_X1    g724(.A(new_n775), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n901), .A2(new_n911), .A3(new_n903), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n878), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n309), .B(KEYINPUT57), .Z(new_n915));
  AOI21_X1  g729(.A(new_n704), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n907), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(KEYINPUT118), .B(new_n907), .C1(new_n912), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(G54));
  INV_X1    g735(.A(new_n498), .ZN(new_n922));
  NAND2_X1  g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n904), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n907), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n904), .A2(new_n922), .A3(new_n923), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(G60));
  XOR2_X1   g741(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n928));
  NOR2_X1   g742(.A1(new_n549), .A2(new_n188), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n914), .A2(new_n606), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n606), .B1(new_n884), .B2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n906), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n900), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n638), .B2(new_n639), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n907), .C1(new_n592), .C2(new_n936), .ZN(new_n938));
  XOR2_X1   g752(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G66));
  INV_X1    g754(.A(G224), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n394), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT121), .ZN(new_n943));
  INV_X1    g757(.A(new_n863), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n190), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n415), .B(new_n416), .C1(G898), .C2(new_n190), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(G69));
  AND2_X1   g761(.A1(new_n797), .A2(new_n793), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n736), .A2(new_n845), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT62), .B1(new_n692), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n751), .A2(new_n714), .A3(new_n830), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n674), .A2(new_n756), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT123), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n692), .A2(KEYINPUT62), .A3(new_n949), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n948), .A2(new_n950), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n190), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n352), .A2(new_n353), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n491), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n190), .A2(G900), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT124), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AND4_X1   g777(.A1(new_n757), .A2(new_n782), .A3(new_n729), .A4(new_n731), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n949), .B1(new_n763), .B2(new_n768), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n948), .A3(new_n766), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n963), .B1(new_n967), .B2(new_n190), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n960), .B1(new_n968), .B2(new_n958), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G72));
  INV_X1    g785(.A(new_n356), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n347), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  NOR2_X1   g790(.A1(new_n356), .A2(new_n359), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT126), .Z(new_n980));
  NOR2_X1   g794(.A1(new_n883), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n967), .B2(new_n944), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n973), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n976), .B1(new_n955), .B2(new_n944), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n906), .B1(new_n985), .B2(new_n977), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n982), .A2(new_n984), .A3(new_n986), .ZN(G57));
endmodule


