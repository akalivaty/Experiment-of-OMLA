//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G217));
  OR4_X1    g029(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g036(.A(G261), .ZN(G325));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n464), .B1(new_n457), .B2(G2106), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT69), .ZN(G319));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n472), .B(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n469), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G137), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n479), .A2(G136), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT71), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n469), .A2(new_n484), .ZN(new_n485));
  MUX2_X1   g060(.A(G100), .B(G112), .S(G2105), .Z(new_n486));
  AOI22_X1  g061(.A1(new_n485), .A2(G124), .B1(G2104), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n488), .B(new_n489), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(new_n476), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n493), .B2(new_n494), .ZN(new_n499));
  AND2_X1   g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n484), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n484), .C1(new_n467), .C2(new_n468), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT73), .Z(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n507), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(new_n520), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  XNOR2_X1  g100(.A(new_n508), .B(KEYINPUT75), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n528), .B(new_n530), .C1(new_n521), .C2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n526), .A2(G52), .B1(G90), .B2(new_n522), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n519), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AND2_X1   g113(.A1(new_n515), .A2(new_n516), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  INV_X1    g115(.A(G68), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n514), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI221_X1 g119(.A(KEYINPUT76), .B1(new_n541), .B2(new_n514), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G651), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n526), .A2(G43), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT77), .B(G81), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n522), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n508), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n508), .B2(new_n559), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n560), .A2(new_n561), .B1(new_n522), .B2(G91), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n515), .B2(new_n516), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  AND2_X1   g140(.A1(G78), .A2(G543), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G651), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n562), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n522), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n509), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(new_n517), .A2(G61), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT80), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n519), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n522), .A2(G86), .B1(G48), .B2(new_n509), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n526), .A2(G47), .B1(G85), .B2(new_n522), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n519), .B2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n522), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n526), .A2(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n519), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(new_n588), .ZN(G284));
  AOI21_X1  g172(.A(new_n589), .B1(new_n596), .B2(new_n588), .ZN(G321));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT82), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(G868), .B2(new_n601), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(G868), .B2(new_n601), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G860), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT83), .ZN(G148));
  NOR2_X1   g181(.A1(new_n550), .A2(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n595), .A2(G559), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n479), .A2(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT13), .B(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n479), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n485), .A2(G123), .ZN(new_n617));
  AND2_X1   g192(.A1(G111), .A2(G2105), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(G99), .B2(new_n484), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n476), .C2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  XOR2_X1   g201(.A(G2443), .B(G2446), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT15), .B(G2435), .Z(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT86), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n630), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT87), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT88), .Z(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  INV_X1    g225(.A(new_n646), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .A3(new_n644), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n644), .B1(new_n651), .B2(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n648), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n645), .A2(new_n648), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n655), .B2(KEYINPUT17), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n650), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(new_n621), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2100), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n662), .A2(new_n665), .A3(new_n670), .ZN(new_n672));
  NAND4_X1  g247(.A1(new_n668), .A2(new_n669), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G25), .ZN(new_n681));
  MUX2_X1   g256(.A(G95), .B(G107), .S(G2105), .Z(new_n682));
  AOI22_X1  g257(.A1(new_n485), .A2(G119), .B1(G2104), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G131), .ZN(new_n684));
  INV_X1    g259(.A(new_n479), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n681), .B1(new_n687), .B2(new_n680), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT35), .B(G1991), .Z(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  NAND2_X1  g265(.A1(G290), .A2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G24), .ZN(new_n692));
  OAI21_X1  g267(.A(KEYINPUT91), .B1(new_n692), .B2(G16), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n692), .A2(KEYINPUT91), .A3(G16), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  NOR2_X1   g271(.A1(G16), .A2(G23), .ZN(new_n697));
  INV_X1    g272(.A(G288), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT92), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT33), .B(G1976), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT93), .Z(new_n702));
  XOR2_X1   g277(.A(new_n700), .B(new_n702), .Z(new_n703));
  NOR2_X1   g278(.A1(G6), .A2(G16), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n583), .B2(G16), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G22), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G166), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1971), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n703), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n690), .B(new_n696), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT36), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n713), .A2(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n715), .B2(new_n716), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n713), .A2(KEYINPUT94), .A3(KEYINPUT36), .A4(new_n714), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G20), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT23), .Z(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G299), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1956), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n680), .A2(G33), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n477), .A2(G103), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT25), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(KEYINPUT25), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n727), .A2(new_n728), .B1(G139), .B2(new_n479), .ZN(new_n729));
  INV_X1    g304(.A(new_n469), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(new_n484), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G2072), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT97), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n620), .A2(new_n680), .ZN(new_n737));
  OR2_X1    g312(.A1(KEYINPUT30), .A2(G28), .ZN(new_n738));
  NAND2_X1  g313(.A1(KEYINPUT30), .A2(G28), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  NOR3_X1   g316(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n680), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT98), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n680), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n742), .B1(new_n743), .B2(new_n749), .C1(new_n733), .C2(new_n734), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n736), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G171), .A2(new_n720), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G5), .B2(new_n720), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n720), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n720), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1966), .ZN(new_n758));
  NOR2_X1   g333(.A1(G27), .A2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G164), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  AND4_X1   g337(.A1(new_n724), .A2(new_n751), .A3(new_n755), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G32), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n485), .A2(G129), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT99), .Z(new_n766));
  AND2_X1   g341(.A1(new_n477), .A2(G105), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n767), .B(new_n769), .C1(G141), .C2(new_n479), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n764), .B1(new_n772), .B2(G29), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT100), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT101), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n753), .A2(new_n754), .B1(new_n743), .B2(new_n749), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n774), .B2(new_n775), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT102), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n680), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n680), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT29), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n779), .A2(new_n780), .B1(G2090), .B2(new_n784), .ZN(new_n785));
  AND4_X1   g360(.A1(new_n763), .A2(new_n777), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n784), .A2(G2090), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT103), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n596), .A2(G16), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G4), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT95), .B(G1348), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G19), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n551), .B2(G16), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1341), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n790), .A2(new_n791), .ZN(new_n796));
  MUX2_X1   g371(.A(G104), .B(G116), .S(G2105), .Z(new_n797));
  AOI22_X1  g372(.A1(new_n485), .A2(G128), .B1(G2104), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G140), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n685), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n680), .A2(G26), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT28), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n792), .A2(new_n795), .A3(new_n796), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT96), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n788), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n718), .A2(new_n719), .A3(new_n786), .A4(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  INV_X1    g387(.A(G67), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n539), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n519), .B1(new_n814), .B2(KEYINPUT104), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(KEYINPUT104), .B2(new_n814), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n526), .A2(G55), .B1(G93), .B2(new_n522), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n550), .B(KEYINPUT105), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n818), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n595), .A2(new_n604), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n820), .B1(new_n829), .B2(new_n831), .ZN(G145));
  MUX2_X1   g407(.A(G106), .B(G118), .S(G2105), .Z(new_n833));
  AOI22_X1  g408(.A1(new_n485), .A2(G130), .B1(G2104), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G142), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n685), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n686), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n613), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n800), .B(new_n505), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n771), .B(new_n732), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(G162), .B(G160), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(new_n620), .Z(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n842), .A3(new_n843), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g427(.A(new_n824), .B(new_n608), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n595), .B(new_n601), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT41), .Z(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n854), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(new_n853), .ZN(new_n858));
  XNOR2_X1  g433(.A(G305), .B(G303), .ZN(new_n859));
  XNOR2_X1  g434(.A(G290), .B(G288), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n858), .A2(KEYINPUT107), .A3(new_n863), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n866), .B(new_n867), .C1(new_n863), .C2(new_n858), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n818), .A2(new_n588), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(G295));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n870), .ZN(G331));
  XNOR2_X1  g447(.A(G301), .B(KEYINPUT108), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G286), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n824), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(G168), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n822), .A3(new_n823), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n855), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n877), .A3(new_n854), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n861), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n849), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n861), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT43), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n849), .A4(new_n881), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT44), .Z(G397));
  NAND2_X1  g464(.A1(G160), .A2(G40), .ZN(new_n890));
  INV_X1    g465(.A(G1384), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n505), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT45), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G1996), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT109), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n800), .B(G2067), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n772), .B2(new_n897), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n899), .A2(new_n772), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT110), .Z(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n687), .A3(new_n689), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n800), .A2(G2067), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n896), .B1(new_n772), .B2(new_n901), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n899), .B2(KEYINPUT46), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(KEYINPUT46), .B2(new_n899), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT47), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n686), .B(new_n689), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n904), .B1(new_n896), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n896), .A2(G1986), .A3(G290), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT126), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT48), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n913), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n908), .A2(new_n909), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G40), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n748), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n891), .A3(new_n505), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT112), .B(G8), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT114), .B(G1981), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n583), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n582), .ZN(new_n929));
  OAI21_X1  g504(.A(G1981), .B1(new_n929), .B2(new_n579), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT49), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(new_n926), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT113), .B1(new_n698), .B2(G1976), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n698), .A2(G1976), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n937), .A2(new_n940), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n892), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n891), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n890), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G2090), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n891), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n894), .A2(new_n922), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1971), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n948), .A2(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT111), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n957), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n955), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n959), .B1(new_n924), .B2(new_n953), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n944), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n894), .A2(new_n950), .ZN(new_n967));
  INV_X1    g542(.A(G2078), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n922), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n891), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT50), .B1(new_n505), .B2(new_n891), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n922), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n969), .A2(new_n970), .B1(new_n754), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n970), .B2(new_n969), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G171), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n743), .B(new_n922), .C1(new_n971), .C2(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT115), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n946), .A2(new_n947), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n743), .A4(new_n922), .ZN(new_n981));
  INV_X1    g556(.A(G1966), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n951), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(G168), .A2(new_n924), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT121), .A3(KEYINPUT51), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT121), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n986), .B1(new_n984), .B2(G8), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n984), .A2(new_n925), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(new_n992), .A3(new_n987), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n989), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n984), .A2(new_n986), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(KEYINPUT62), .A3(new_n997), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n976), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT56), .B(G2072), .Z(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT118), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n894), .A2(new_n922), .A3(new_n950), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n948), .B2(G1956), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1007));
  NAND2_X1  g582(.A1(G299), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1007), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n562), .A2(new_n569), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n890), .A2(new_n892), .ZN(new_n1014));
  INV_X1    g589(.A(G1348), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n805), .A2(new_n1014), .B1(new_n973), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n595), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1011), .B(new_n1005), .C1(new_n948), .C2(G1956), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT120), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(KEYINPUT61), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT61), .ZN(new_n1022));
  AOI211_X1 g597(.A(KEYINPUT120), .B(new_n1022), .C1(new_n1013), .C2(new_n1018), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1016), .A2(new_n595), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1016), .A2(new_n595), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT60), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n967), .A2(new_n897), .A3(new_n922), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT58), .B(G1341), .Z(new_n1029));
  NAND2_X1  g604(.A1(new_n923), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n550), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(KEYINPUT119), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1031), .A2(new_n1033), .B1(new_n1016), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1027), .B(new_n1035), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1019), .B1(new_n1024), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(G301), .B(KEYINPUT54), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n922), .B(KEYINPUT122), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(KEYINPUT53), .A3(new_n968), .A4(new_n967), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1040), .A2(KEYINPUT123), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(KEYINPUT123), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1043), .A2(new_n974), .B1(new_n975), .B2(new_n1038), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1037), .A2(new_n998), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n966), .B1(new_n1002), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n963), .A2(new_n943), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n934), .A2(new_n1048), .A3(new_n698), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n928), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n935), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1053));
  NOR2_X1   g628(.A1(new_n994), .A2(G286), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1053), .B1(new_n965), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n959), .B1(new_n954), .B2(new_n953), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n963), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(KEYINPUT63), .A3(new_n944), .A4(new_n1054), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1052), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1046), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(G290), .B(G1986), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n915), .B1(new_n895), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT124), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n976), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n996), .A2(KEYINPUT62), .A3(new_n997), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT62), .B1(new_n996), .B2(new_n997), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1037), .A2(new_n998), .A3(new_n1044), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n965), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1051), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT124), .B(new_n1063), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n920), .B1(new_n1064), .B2(new_n1074), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g650(.A1(G319), .A2(new_n659), .ZN(new_n1077));
  NOR2_X1   g651(.A1(new_n1077), .A2(G229), .ZN(new_n1078));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n642), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g653(.A(new_n1079), .B1(new_n884), .B2(new_n887), .ZN(new_n1080));
  INV_X1    g654(.A(KEYINPUT127), .ZN(new_n1081));
  XNOR2_X1  g655(.A(new_n1080), .B(new_n1081), .ZN(G308));
  XNOR2_X1  g656(.A(new_n1080), .B(KEYINPUT127), .ZN(G225));
endmodule


