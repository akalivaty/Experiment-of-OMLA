//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  AOI22_X1  g003(.A1(new_n203), .A2(new_n204), .B1(G29gat), .B2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT84), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT84), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT14), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(KEYINPUT14), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n203), .A2(new_n204), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n214), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n202), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT88), .A4(KEYINPUT17), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT85), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT16), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(KEYINPUT16), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G8gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n227), .B(new_n228), .C1(G1gat), .C2(new_n222), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT87), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n227), .B(KEYINPUT86), .C1(G1gat), .C2(new_n222), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(G8gat), .C1(KEYINPUT86), .C2(new_n227), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT17), .B1(new_n215), .B2(new_n216), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n217), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n239), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n234), .A2(new_n217), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT89), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n239), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n238), .B(KEYINPUT13), .Z(new_n247));
  NAND3_X1  g046(.A1(new_n234), .A2(KEYINPUT89), .A3(new_n217), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G197gat), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT11), .B(G169gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT12), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n255), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n242), .A2(new_n249), .A3(new_n257), .A4(new_n243), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT27), .B(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT26), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT23), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n266), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n267), .B2(KEYINPUT23), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n265), .A2(KEYINPUT24), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(G183gat), .A3(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G183gat), .B2(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(new_n262), .A3(KEYINPUT65), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n274), .B1(new_n283), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n280), .A2(new_n282), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n284), .A2(new_n286), .B1(new_n290), .B2(new_n262), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n266), .A2(KEYINPUT67), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(G169gat), .A3(G176gat), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n277), .A2(new_n296), .A3(new_n298), .A4(KEYINPUT25), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n293), .A2(new_n300), .A3(KEYINPUT68), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(new_n274), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n280), .A2(new_n282), .ZN(new_n304));
  INV_X1    g103(.A(new_n278), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n290), .A2(KEYINPUT24), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n307), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n265), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n289), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n303), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n295), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n277), .A2(KEYINPUT25), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n312), .A2(new_n304), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n302), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n273), .B1(new_n301), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n323));
  INV_X1    g122(.A(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G127gat), .ZN(new_n325));
  INV_X1    g124(.A(G127gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G134gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n322), .A2(new_n323), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n327), .ZN(new_n329));
  XNOR2_X1  g128(.A(G113gat), .B(G120gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n323), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT70), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT70), .B1(new_n328), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT68), .B1(new_n293), .B2(new_n300), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n311), .A2(new_n302), .A3(new_n315), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n272), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n335), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G71gat), .B(G99gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT33), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(KEYINPUT32), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT71), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n343), .A2(new_n350), .A3(KEYINPUT32), .A4(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(KEYINPUT32), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n355), .A3(new_n346), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n338), .B1(new_n337), .B2(new_n342), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT34), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n358), .A2(new_n359), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  NAND2_X1  g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT2), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT77), .ZN(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G141gat), .B(G148gat), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n369), .A2(KEYINPUT2), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G141gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G148gat), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G141gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n370), .B(new_n380), .C1(new_n383), .C2(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n368), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n375), .C2(new_n384), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n367), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT22), .ZN(new_n390));
  INV_X1    g189(.A(G211gat), .ZN(new_n391));
  INV_X1    g190(.A(G218gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G197gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT73), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G197gat), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n395), .A2(new_n397), .A3(G204gat), .ZN(new_n398));
  AOI21_X1  g197(.A(G204gat), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G211gat), .B(G218gat), .Z(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n401), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n403), .B(new_n393), .C1(new_n398), .C2(new_n399), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n375), .A2(new_n384), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n402), .B2(new_n404), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(KEYINPUT3), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n366), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT74), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n402), .A2(KEYINPUT74), .A3(new_n404), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n389), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n366), .A2(new_n411), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n365), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G78gat), .B(G106gat), .Z(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT31), .B(G50gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n418), .A2(new_n412), .A3(new_n410), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n412), .B1(new_n407), .B2(new_n410), .ZN(new_n426));
  OAI21_X1  g225(.A(G22gat), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n366), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n418), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n420), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n421), .A2(new_n424), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  AND4_X1   g230(.A1(KEYINPUT80), .A2(new_n427), .A3(new_n430), .A4(new_n424), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n352), .A2(new_n362), .A3(new_n356), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n364), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n417), .ZN(new_n436));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n438));
  OAI22_X1  g237(.A1(new_n293), .A2(new_n300), .B1(new_n264), .B2(new_n271), .ZN(new_n439));
  INV_X1    g238(.A(new_n437), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT75), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(KEYINPUT75), .B(new_n437), .C1(new_n341), .C2(KEYINPUT29), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n436), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n341), .A2(new_n440), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n439), .A2(new_n367), .A3(new_n437), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n406), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g252(.A1(new_n445), .A2(new_n446), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n440), .B1(new_n317), .B2(new_n367), .ZN(new_n455));
  INV_X1    g254(.A(new_n442), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n444), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n417), .ZN(new_n458));
  INV_X1    g257(.A(new_n449), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n445), .A2(new_n449), .A3(new_n453), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(KEYINPUT30), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n328), .A2(new_n332), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n408), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n385), .A2(new_n328), .A3(new_n332), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G225gat), .A2(G233gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n465), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n375), .A2(new_n384), .A3(KEYINPUT3), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n473), .A2(new_n466), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n387), .B2(new_n388), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n470), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n466), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n385), .B1(new_n333), .B2(new_n334), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(KEYINPUT4), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n472), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n478), .B2(KEYINPUT4), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(new_n465), .A3(new_n475), .A4(new_n470), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(G1gat), .B(G29gat), .Z(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G57gat), .B(G85gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(KEYINPUT6), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(new_n484), .B2(new_n489), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n489), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n480), .A2(new_n493), .A3(new_n483), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n458), .A2(new_n459), .A3(new_n452), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT76), .A3(new_n446), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n461), .A2(new_n464), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT35), .B1(new_n435), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT83), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT83), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(KEYINPUT35), .C1(new_n435), .C2(new_n499), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n453), .B1(new_n445), .B2(new_n449), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n449), .B1(new_n457), .B2(new_n417), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n452), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT30), .B1(new_n505), .B2(new_n452), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n504), .B(new_n506), .C1(new_n507), .C2(KEYINPUT76), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n385), .B(new_n466), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT5), .B1(new_n510), .B2(new_n470), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT78), .B1(new_n408), .B2(KEYINPUT3), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n385), .A2(new_n368), .A3(new_n386), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n471), .B1(new_n514), .B2(new_n474), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n478), .A2(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(KEYINPUT4), .B2(new_n468), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n511), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AND4_X1   g317(.A1(new_n465), .A2(new_n482), .A3(new_n470), .A4(new_n475), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n489), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT81), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n494), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n490), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n491), .B2(new_n494), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n509), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n498), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n508), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n364), .A2(KEYINPUT82), .A3(new_n434), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT82), .ZN(new_n530));
  INV_X1    g329(.A(new_n434), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n362), .B1(new_n352), .B2(new_n356), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(new_n433), .A3(new_n529), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n501), .A2(new_n503), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n452), .B1(new_n505), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(new_n536), .B2(new_n505), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT38), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n447), .A2(new_n406), .A3(new_n448), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n457), .B2(new_n417), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT38), .B1(new_n541), .B2(KEYINPUT37), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n537), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n524), .A2(new_n525), .A3(new_n463), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n470), .B1(new_n482), .B2(new_n475), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n489), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT39), .B1(new_n469), .B2(new_n471), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n552), .A2(new_n520), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n508), .B2(new_n527), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n545), .A2(new_n555), .A3(new_n433), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n364), .A2(new_n434), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT72), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(KEYINPUT72), .A3(KEYINPUT36), .ZN(new_n561));
  INV_X1    g360(.A(new_n433), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n499), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n556), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n260), .B1(new_n535), .B2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G120gat), .B(G148gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT100), .ZN(new_n567));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G57gat), .B(G64gat), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G57gat), .B(G64gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n576), .B1(new_n574), .B2(KEYINPUT90), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n582));
  OAI221_X1 g381(.A(new_n581), .B1(KEYINPUT90), .B2(new_n576), .C1(new_n578), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT93), .Z(new_n585));
  XOR2_X1   g384(.A(KEYINPUT95), .B(G92gat), .Z(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  INV_X1    g389(.A(G99gat), .ZN(new_n591));
  INV_X1    g390(.A(G106gat), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT8), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G99gat), .B(G106gat), .Z(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT10), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n585), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(KEYINPUT98), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(new_n583), .A3(new_n580), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n584), .B1(KEYINPUT98), .B2(new_n594), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n594), .B(new_n595), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n599), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n596), .A2(new_n601), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n604), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(KEYINPUT99), .A3(new_n599), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n598), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n611), .A2(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n570), .B1(new_n618), .B2(KEYINPUT101), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n620), .B(new_n569), .C1(new_n616), .C2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G232gat), .ZN(new_n623));
  INV_X1    g422(.A(G233gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT94), .ZN(new_n627));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G134gat), .B(G162gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI211_X1 g433(.A(new_n235), .B(new_n596), .C1(new_n219), .C2(new_n220), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n217), .B2(new_n596), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n604), .B1(new_n216), .B2(new_n215), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT96), .B1(new_n640), .B2(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n629), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n634), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI221_X1 g444(.A(new_n633), .B1(new_n629), .B2(new_n628), .C1(new_n635), .C2(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n584), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G127gat), .B(G155gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT20), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G183gat), .B(G211gat), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n233), .B(new_n231), .C1(new_n585), .C2(new_n648), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n654), .A2(new_n656), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n657), .B2(new_n661), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n647), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n622), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n565), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n565), .A2(KEYINPUT102), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n496), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  INV_X1    g473(.A(new_n508), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n498), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n669), .B2(new_n670), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT103), .B1(new_n678), .B2(new_n228), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n678), .A2(KEYINPUT103), .A3(new_n228), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n679), .B(new_n680), .C1(new_n683), .C2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(new_n671), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n560), .A2(new_n561), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G15gat), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(G15gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n533), .A2(new_n529), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n671), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(G1326gat));
  OAI21_X1  g493(.A(KEYINPUT104), .B1(new_n686), .B2(new_n433), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n671), .A2(new_n696), .A3(new_n562), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n698), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(new_n622), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n662), .A2(new_n663), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n260), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n535), .A2(new_n564), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n535), .A2(new_n564), .A3(KEYINPUT105), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n710), .A2(new_n711), .A3(new_n647), .A4(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n647), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n535), .B2(new_n564), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT44), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n707), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n496), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n715), .A2(new_n206), .A3(new_n672), .A4(new_n706), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(G1328gat));
  OAI21_X1  g522(.A(G36gat), .B1(new_n719), .B2(new_n677), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n705), .A2(new_n714), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n565), .A2(new_n207), .A3(new_n676), .A4(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT106), .B(KEYINPUT46), .Z(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(G1329gat));
  NAND2_X1  g528(.A1(new_n718), .A2(new_n687), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n705), .A2(G43gat), .A3(new_n691), .A4(new_n714), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(G43gat), .B1(new_n565), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n562), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT107), .B1(new_n433), .B2(G50gat), .ZN(new_n735));
  OR3_X1    g534(.A1(new_n433), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n725), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n734), .A2(G50gat), .B1(new_n565), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g538(.A1(new_n535), .A2(KEYINPUT105), .A3(new_n564), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT105), .B1(new_n535), .B2(new_n564), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n703), .ZN(new_n743));
  NOR4_X1   g542(.A1(new_n622), .A2(new_n743), .A3(new_n259), .A4(new_n647), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n672), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g547(.A(new_n676), .B(KEYINPUT108), .Z(new_n749));
  NOR2_X1   g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n745), .B2(new_n688), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n691), .A2(G71gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n745), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n746), .A2(new_n562), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n259), .A2(new_n703), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n622), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n713), .B2(new_n717), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n496), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT51), .B1(new_n715), .B2(new_n762), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n715), .A2(KEYINPUT51), .A3(new_n762), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n622), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n587), .A3(new_n672), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n773), .ZN(G1336gat));
  INV_X1    g573(.A(new_n586), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n767), .B2(new_n749), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  AND4_X1   g576(.A1(KEYINPUT51), .A2(new_n708), .A3(new_n647), .A4(new_n762), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n749), .A2(G92gat), .A3(new_n622), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(KEYINPUT110), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(KEYINPUT110), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n778), .A2(new_n769), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n647), .A2(new_n711), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n740), .A2(new_n741), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n715), .A2(new_n711), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n676), .B(new_n764), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n775), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n782), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n789), .B2(KEYINPUT52), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n791), .B(new_n777), .C1(new_n788), .C2(new_n782), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n783), .B1(new_n790), .B2(new_n792), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n767), .B2(new_n688), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n772), .A2(new_n591), .A3(new_n692), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1338gat));
  AOI21_X1  g595(.A(new_n592), .B1(new_n766), .B2(new_n562), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n702), .A2(new_n592), .A3(new_n562), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n798), .A2(KEYINPUT113), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n778), .B2(new_n769), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n562), .B(new_n764), .C1(new_n785), .C2(new_n786), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n807), .A2(new_n808), .A3(new_n803), .A4(new_n802), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n806), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT112), .B1(new_n806), .B2(G106gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n799), .A2(new_n813), .A3(new_n800), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n799), .B2(new_n800), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n778), .B2(new_n769), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n816), .B(KEYINPUT115), .C1(new_n778), .C2(new_n769), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n811), .A2(new_n812), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n810), .B1(new_n822), .B2(new_n803), .ZN(G1339gat));
  OAI21_X1  g622(.A(KEYINPUT117), .B1(new_n665), .B2(new_n259), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n622), .A2(new_n260), .A3(new_n825), .A4(new_n664), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n613), .A2(new_n615), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT99), .B1(new_n611), .B2(new_n599), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n607), .B(KEYINPUT10), .C1(new_n609), .C2(new_n610), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n830), .A2(new_n831), .B1(new_n585), .B2(new_n597), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n614), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n829), .A2(new_n833), .A3(KEYINPUT54), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n570), .B1(new_n833), .B2(KEYINPUT54), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n238), .B1(new_n237), .B2(new_n239), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n254), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n647), .A2(new_n258), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n618), .A2(new_n569), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n569), .B1(new_n616), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n829), .A2(new_n833), .A3(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n845));
  AND4_X1   g644(.A1(new_n836), .A2(new_n840), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n836), .A2(new_n259), .A3(new_n841), .A4(new_n845), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n619), .A2(new_n258), .A3(new_n621), .A4(new_n839), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n849), .B2(new_n714), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n827), .B1(new_n850), .B2(new_n703), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT118), .ZN(new_n852));
  INV_X1    g651(.A(new_n435), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n827), .B(new_n854), .C1(new_n850), .C2(new_n703), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(new_n672), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n858), .A3(new_n749), .ZN(new_n859));
  INV_X1    g658(.A(new_n749), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT119), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n260), .A2(G113gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n852), .A2(new_n855), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n692), .A2(new_n433), .ZN(new_n866));
  NOR4_X1   g665(.A1(new_n865), .A2(new_n496), .A3(new_n866), .A4(new_n860), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n320), .B1(new_n867), .B2(new_n259), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(new_n869), .A3(KEYINPUT120), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  INV_X1    g670(.A(new_n863), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n859), .B2(new_n861), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n873), .B2(new_n868), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(G1340gat));
  NAND3_X1  g674(.A1(new_n862), .A2(new_n318), .A3(new_n702), .ZN(new_n876));
  INV_X1    g675(.A(new_n867), .ZN(new_n877));
  OAI21_X1  g676(.A(G120gat), .B1(new_n877), .B2(new_n622), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1341gat));
  OAI21_X1  g678(.A(G127gat), .B1(new_n877), .B2(new_n743), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n857), .A2(new_n326), .A3(new_n703), .A4(new_n749), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1342gat));
  OAI21_X1  g681(.A(G134gat), .B1(new_n877), .B2(new_n714), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n676), .A2(new_n714), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n857), .A2(new_n324), .A3(new_n884), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(G1343gat));
  XOR2_X1   g687(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n889));
  NAND3_X1  g688(.A1(new_n749), .A2(new_n672), .A3(new_n688), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n852), .A2(new_n562), .A3(new_n855), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n846), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n714), .B1(new_n849), .B2(KEYINPUT121), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n847), .B2(new_n848), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n743), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n827), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n433), .A2(new_n892), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n890), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n376), .B1(new_n903), .B2(new_n259), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n688), .A2(new_n562), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n865), .A2(new_n496), .A3(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n906), .A2(new_n376), .A3(new_n259), .A4(new_n749), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n889), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n889), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n260), .B(new_n890), .C1(new_n893), .C2(new_n902), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n910), .B(new_n907), .C1(new_n911), .C2(new_n376), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(G1344gat));
  NOR2_X1   g712(.A1(new_n622), .A2(G148gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n906), .A2(new_n749), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n898), .A2(new_n743), .B1(new_n260), .B2(new_n666), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n892), .B1(new_n919), .B2(new_n433), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n852), .A2(new_n855), .A3(new_n901), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n890), .A2(new_n622), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n918), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  AOI211_X1 g724(.A(KEYINPUT59), .B(new_n378), .C1(new_n903), .C2(new_n702), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(G1345gat));
  INV_X1    g726(.A(new_n903), .ZN(new_n928));
  OAI21_X1  g727(.A(G155gat), .B1(new_n928), .B2(new_n743), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n743), .A2(G155gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n906), .A2(new_n749), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1346gat));
  OAI21_X1  g731(.A(G162gat), .B1(new_n928), .B2(new_n714), .ZN(new_n933));
  INV_X1    g732(.A(G162gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n906), .A2(new_n934), .A3(new_n884), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n865), .A2(new_n866), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n677), .A2(new_n672), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n275), .A3(new_n260), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n865), .A2(new_n672), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n749), .A2(new_n435), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(KEYINPUT124), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n259), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n940), .B1(new_n946), .B2(new_n275), .ZN(G1348gat));
  NAND4_X1  g746(.A1(new_n944), .A2(new_n276), .A3(new_n702), .A4(new_n945), .ZN(new_n948));
  OAI21_X1  g747(.A(G176gat), .B1(new_n939), .B2(new_n622), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n939), .B2(new_n743), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n941), .A2(new_n261), .A3(new_n703), .A4(new_n942), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT60), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1350gat));
  NAND4_X1  g756(.A1(new_n944), .A2(new_n262), .A3(new_n647), .A4(new_n945), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n937), .A2(new_n647), .A3(new_n938), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n262), .B1(new_n959), .B2(KEYINPUT61), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(new_n960), .A3(new_n962), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n958), .B1(new_n963), .B2(new_n965), .ZN(G1351gat));
  NAND2_X1  g765(.A1(new_n688), .A2(new_n938), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n260), .B(new_n967), .C1(new_n920), .C2(new_n921), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT127), .ZN(new_n969));
  OAI21_X1  g768(.A(G197gat), .B1(new_n968), .B2(KEYINPUT127), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n905), .A2(new_n749), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n941), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n259), .A2(new_n394), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n972), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  OAI22_X1  g776(.A1(new_n969), .A2(new_n970), .B1(new_n975), .B2(new_n977), .ZN(G1352gat));
  AOI21_X1  g777(.A(new_n967), .B1(new_n920), .B2(new_n921), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(G204gat), .B1(new_n980), .B2(new_n622), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n622), .A2(G204gat), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(KEYINPUT62), .B1(new_n972), .B2(new_n983), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n972), .A2(KEYINPUT62), .A3(new_n983), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(G1353gat));
  INV_X1    g785(.A(new_n972), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(new_n391), .A3(new_n703), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n979), .A2(new_n703), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT63), .ZN(new_n991));
  AOI211_X1 g790(.A(new_n991), .B(new_n391), .C1(new_n979), .C2(new_n703), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n990), .B2(new_n992), .ZN(G1354gat));
  OAI21_X1  g792(.A(G218gat), .B1(new_n980), .B2(new_n714), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n987), .A2(new_n392), .A3(new_n647), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


