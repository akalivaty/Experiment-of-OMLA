//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT2), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(KEYINPUT73), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n222), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(KEYINPUT1), .B2(new_n220), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT73), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n226), .B1(new_n209), .B2(new_n211), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n217), .A3(new_n215), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n219), .A2(new_n223), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT4), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n216), .A2(new_n218), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n217), .B1(new_n227), .B2(new_n215), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(new_n225), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n236), .A3(new_n228), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n232), .B2(new_n233), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n219), .A2(KEYINPUT74), .A3(new_n228), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n235), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n231), .B(new_n238), .C1(new_n242), .C2(KEYINPUT4), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n244));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n243), .A2(KEYINPUT78), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT78), .B1(new_n243), .B2(new_n248), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n246), .B1(new_n229), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n238), .ZN(new_n255));
  AOI211_X1 g054(.A(new_n253), .B(new_n235), .C1(new_n240), .C2(new_n241), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n235), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n232), .A2(new_n233), .A3(new_n239), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT74), .B1(new_n219), .B2(new_n228), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT4), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(KEYINPUT75), .A3(new_n238), .A4(new_n254), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n228), .A2(new_n219), .B1(new_n223), .B2(new_n225), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n230), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n244), .B1(new_n265), .B2(new_n245), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT77), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT77), .ZN(new_n269));
  AOI211_X1 g068(.A(new_n269), .B(new_n266), .C1(new_n257), .C2(new_n262), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n207), .B(new_n251), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n206), .B(KEYINPUT81), .Z(new_n274));
  AND2_X1   g073(.A1(new_n254), .A2(new_n238), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT75), .B1(new_n275), .B2(new_n261), .ZN(new_n276));
  INV_X1    g075(.A(new_n262), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n267), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n269), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n263), .A2(KEYINPUT77), .A3(new_n267), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n281), .B2(new_n251), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT84), .B1(new_n273), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n251), .B1(new_n268), .B2(new_n270), .ZN(new_n284));
  INV_X1    g083(.A(new_n274), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT84), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n272), .A4(new_n271), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(KEYINPUT6), .A3(new_n206), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT79), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n284), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(new_n206), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295));
  AND2_X1   g094(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n297));
  INV_X1    g096(.A(G211gat), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n299), .B2(KEYINPUT22), .ZN(new_n300));
  INV_X1    g099(.A(new_n297), .ZN(new_n301));
  NAND2_X1  g100(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(G211gat), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT22), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G197gat), .B(G204gat), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n295), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n295), .ZN(new_n311));
  AOI211_X1 g110(.A(new_n308), .B(new_n311), .C1(new_n300), .C2(new_n306), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT23), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(G183gat), .B2(G190gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n321), .B(KEYINPUT25), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n326), .B2(new_n322), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n322), .A2(new_n326), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n320), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n325), .B1(new_n330), .B2(KEYINPUT25), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT66), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT27), .ZN(new_n333));
  INV_X1    g132(.A(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n336));
  AOI21_X1  g135(.A(G190gat), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n338));
  OAI21_X1  g137(.A(new_n332), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G190gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n336), .ZN(new_n341));
  NOR2_X1   g140(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(KEYINPUT66), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n337), .A2(KEYINPUT28), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n339), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n349), .A2(new_n350), .B1(G183gat), .B2(G190gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(KEYINPUT67), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT67), .B1(new_n347), .B2(new_n351), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n331), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(KEYINPUT29), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n347), .A2(new_n351), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n331), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(new_n356), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n313), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT71), .B1(new_n365), .B2(new_n356), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n367));
  INV_X1    g166(.A(new_n322), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT64), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n369), .A2(new_n328), .A3(new_n324), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n370), .B2(new_n320), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n371), .A2(new_n325), .B1(new_n347), .B2(new_n351), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n356), .B1(new_n372), .B2(KEYINPUT29), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n324), .A2(new_n322), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n374), .A2(new_n320), .A3(new_n367), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n327), .A2(new_n329), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n321), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n377), .B2(new_n367), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n380), .B2(new_n352), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n373), .B1(new_n381), .B2(new_n356), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n366), .B1(new_n382), .B2(KEYINPUT71), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n363), .B1(new_n383), .B2(new_n313), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT72), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n392));
  INV_X1    g191(.A(new_n366), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n313), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT37), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n362), .B1(new_n355), .B2(new_n358), .ZN(new_n396));
  INV_X1    g195(.A(new_n313), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT38), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n386), .A2(new_n391), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT71), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n355), .A2(new_n357), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n373), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n397), .B1(new_n403), .B2(new_n366), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n391), .B1(new_n404), .B2(new_n363), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT38), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n390), .B1(new_n384), .B2(new_n385), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(KEYINPUT37), .A3(new_n363), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n289), .A2(new_n294), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT31), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G50gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G228gat), .ZN(new_n418));
  INV_X1    g217(.A(G233gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n299), .A2(KEYINPUT70), .A3(KEYINPUT22), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n309), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n311), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n307), .A2(new_n309), .A3(new_n295), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n236), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n364), .B1(new_n310), .B2(new_n312), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n429), .A2(new_n431), .B1(new_n232), .B2(new_n233), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n237), .A2(new_n364), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n313), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n421), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n241), .B(new_n240), .C1(new_n427), .C2(KEYINPUT3), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n437), .A3(new_n421), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n436), .A2(G22gat), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G22gat), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT3), .B1(new_n430), .B2(KEYINPUT80), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n428), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n442), .A2(new_n443), .B1(new_n228), .B2(new_n219), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n420), .B1(new_n444), .B2(new_n434), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n445), .B2(new_n438), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n417), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(G22gat), .B1(new_n436), .B2(new_n439), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n441), .A3(new_n438), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n416), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n243), .A2(KEYINPUT82), .A3(new_n246), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT82), .B1(new_n243), .B2(new_n246), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n452), .B1(new_n265), .B2(new_n245), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n459), .A3(new_n274), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT40), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n460), .A2(KEYINPUT83), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n461), .A2(KEYINPUT83), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n462), .A2(new_n282), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n363), .B(new_n391), .C1(new_n383), .C2(new_n313), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT30), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(new_n405), .ZN(new_n468));
  AOI211_X1 g267(.A(KEYINPUT30), .B(new_n391), .C1(new_n404), .C2(new_n363), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n451), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n413), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(G15gat), .B(G43gat), .Z(new_n473));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(KEYINPUT33), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n355), .A2(new_n235), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n258), .B(new_n331), .C1(new_n353), .C2(new_n354), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G227gat), .A2(G233gat), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT32), .B(new_n478), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n475), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n484), .A2(KEYINPUT33), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n479), .A2(new_n482), .A3(new_n480), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT34), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n489), .B(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(new_n483), .C1(new_n487), .C2(new_n486), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n491), .A2(new_n494), .A3(KEYINPUT36), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT36), .B1(new_n491), .B2(new_n494), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n284), .A2(new_n206), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(new_n272), .A3(new_n271), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n292), .A2(new_n499), .A3(new_n293), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n468), .A2(new_n469), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n497), .B1(new_n502), .B2(new_n451), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n447), .A2(new_n450), .A3(new_n494), .A4(new_n491), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT35), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n506));
  NOR3_X1   g305(.A1(new_n504), .A2(new_n470), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n289), .A2(new_n294), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n472), .A2(new_n503), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT95), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(KEYINPUT41), .ZN(new_n514));
  XOR2_X1   g313(.A(G190gat), .B(G218gat), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n516), .A2(KEYINPUT97), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n514), .B(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT88), .ZN(new_n523));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n521), .B(new_n523), .C1(KEYINPUT15), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n525), .B(new_n526), .Z(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n525), .B(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT8), .ZN(new_n534));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G92gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n203), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n534), .A2(new_n537), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G99gat), .B(G106gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT8), .A2(new_n533), .B1(new_n203), .B2(new_n538), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n545), .A2(new_n542), .A3(new_n537), .A4(new_n540), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n529), .A2(new_n530), .A3(new_n532), .A4(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n513), .A2(KEYINPUT41), .B1(new_n516), .B2(KEYINPUT97), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n530), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n527), .B1(new_n528), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n548), .B(new_n549), .C1(new_n547), .C2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n518), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n518), .A3(new_n556), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n562));
  INV_X1    g361(.A(G1gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G8gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(G8gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  OR2_X1    g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT9), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(KEYINPUT91), .A2(G64gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(KEYINPUT92), .A3(G57gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n580));
  INV_X1    g379(.A(G64gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(G57gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n578), .B1(KEYINPUT92), .B2(G57gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n577), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n574), .B(new_n575), .C1(new_n586), .C2(new_n576), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n572), .B1(new_n573), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n591));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G127gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n213), .ZN(new_n599));
  OR3_X1    g398(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n594), .B2(new_n595), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G183gat), .B(G211gat), .Z(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n560), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n510), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n588), .A2(new_n547), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n585), .A2(new_n544), .A3(new_n587), .A4(new_n546), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT98), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n613), .A2(new_n618), .A3(new_n614), .A4(new_n615), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n615), .B2(new_n614), .ZN(new_n621));
  INV_X1    g420(.A(new_n588), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n622), .A2(new_n550), .A3(KEYINPUT99), .A4(KEYINPUT10), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n617), .A2(new_n619), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n613), .A2(new_n615), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n626), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n612), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n625), .B1(new_n624), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n619), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n623), .A2(new_n621), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n634), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT101), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n629), .ZN(new_n638));
  INV_X1    g437(.A(new_n612), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n629), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT102), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n644), .B(new_n641), .C1(new_n637), .C2(new_n629), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n631), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n529), .A2(new_n572), .A3(new_n532), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n571), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n569), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n527), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n647), .A2(KEYINPUT18), .A3(new_n648), .A4(new_n651), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT90), .B1(new_n527), .B2(new_n650), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT90), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n572), .A2(new_n657), .A3(new_n531), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n651), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n648), .B(KEYINPUT13), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n654), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(G113gat), .B(G141gat), .Z(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT87), .B(G197gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT11), .B(G169gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT12), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n654), .A2(new_n669), .A3(new_n662), .A4(new_n655), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n646), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n609), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n500), .B(KEYINPUT103), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n563), .ZN(G1324gat));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  INV_X1    g480(.A(new_n676), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n470), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT104), .Z(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n683), .A2(new_n681), .A3(new_n685), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n684), .B2(G8gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n497), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n676), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n491), .A2(new_n494), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n682), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n690), .B2(new_n694), .ZN(G1326gat));
  INV_X1    g494(.A(new_n451), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n676), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n472), .A2(new_n503), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n505), .A2(new_n509), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n560), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n606), .A2(new_n607), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n704), .A2(new_n674), .A3(new_n646), .A4(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G29gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n677), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n706), .B1(new_n704), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n702), .A2(KEYINPUT44), .A3(new_n703), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n675), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n678), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n710), .A2(new_n715), .ZN(G1328gat));
  INV_X1    g515(.A(G36gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n707), .A2(new_n717), .A3(new_n470), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(KEYINPUT105), .ZN(new_n720));
  OAI21_X1  g519(.A(G36gat), .B1(new_n714), .B2(new_n501), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(KEYINPUT105), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n723), .ZN(G1329gat));
  OAI21_X1  g523(.A(G43gat), .B1(new_n714), .B2(new_n691), .ZN(new_n725));
  INV_X1    g524(.A(G43gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n707), .A2(new_n726), .A3(new_n693), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g528(.A(G50gat), .B1(new_n714), .B2(new_n696), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n696), .A2(G50gat), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT106), .Z(new_n732));
  NAND2_X1  g531(.A1(new_n707), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g534(.A(new_n631), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n634), .A2(new_n635), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n624), .A2(new_n632), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n625), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n630), .B1(new_n740), .B2(KEYINPUT101), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n644), .B1(new_n741), .B2(new_n641), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n638), .A2(KEYINPUT102), .A3(new_n642), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n736), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n673), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n609), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n677), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT107), .B(G57gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n470), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT49), .B(G64gat), .Z(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT108), .ZN(G1333gat));
  AOI21_X1  g553(.A(G71gat), .B1(new_n746), .B2(new_n693), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n497), .A2(G71gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n746), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g557(.A1(new_n746), .A2(new_n451), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT109), .B(G78gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1335gat));
  OAI21_X1  g560(.A(new_n711), .B1(new_n510), .B2(new_n560), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(new_n713), .A3(new_n705), .A4(new_n745), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT110), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n678), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n706), .A2(new_n673), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n702), .A2(KEYINPUT51), .A3(new_n703), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT111), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n702), .A2(new_n703), .A3(new_n766), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n677), .A2(new_n203), .A3(new_n646), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n765), .B1(new_n772), .B2(new_n773), .ZN(G1336gat));
  INV_X1    g573(.A(new_n772), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n501), .A2(new_n744), .A3(G92gat), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G92gat), .B1(new_n763), .B2(new_n501), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n769), .A2(KEYINPUT112), .A3(new_n770), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT112), .B1(new_n769), .B2(new_n770), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n782), .B2(new_n768), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n713), .A4(new_n745), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n501), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n787), .B2(new_n538), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n788), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT113), .B1(new_n788), .B2(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n779), .B1(new_n789), .B2(new_n790), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n764), .B2(new_n691), .ZN(new_n792));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n693), .A2(new_n646), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n772), .B2(new_n794), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n796), .B(G106gat), .C1(new_n764), .C2(new_n696), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n696), .B1(new_n784), .B2(new_n786), .ZN(new_n798));
  INV_X1    g597(.A(G106gat), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT114), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n696), .A2(G106gat), .A3(new_n744), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n782), .B2(new_n768), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n775), .B2(new_n801), .ZN(new_n805));
  OAI21_X1  g604(.A(G106gat), .B1(new_n763), .B2(new_n696), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n659), .A2(new_n661), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n648), .B1(new_n647), .B2(new_n651), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n668), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n672), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n744), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n813), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT117), .B1(new_n646), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  OAI221_X1 g617(.A(KEYINPUT54), .B1(new_n625), .B2(new_n737), .C1(new_n633), .C2(new_n636), .ZN(new_n819));
  XOR2_X1   g618(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n820));
  AOI21_X1  g619(.A(new_n639), .B1(new_n627), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n643), .A2(new_n645), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT116), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  OAI221_X1 g624(.A(new_n825), .B1(new_n818), .B2(new_n822), .C1(new_n643), .C2(new_n645), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n818), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n824), .A2(new_n826), .A3(new_n673), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n703), .B1(new_n817), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n560), .A2(new_n813), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n830), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n705), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n706), .A2(new_n674), .A3(new_n744), .A4(new_n560), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n678), .A2(new_n470), .A3(new_n504), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n673), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n646), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n706), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n703), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G134gat), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT118), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n844), .A2(G134gat), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(KEYINPUT119), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(KEYINPUT119), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n846), .B(new_n851), .C1(new_n847), .C2(new_n849), .ZN(G1343gat));
  AOI21_X1  g651(.A(new_n696), .B1(new_n833), .B2(new_n834), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n673), .A2(new_n827), .ZN(new_n855));
  OAI22_X1  g654(.A1(new_n823), .A2(new_n855), .B1(new_n744), .B2(new_n813), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n560), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n831), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n834), .B1(new_n858), .B2(new_n706), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n451), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n853), .A2(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n678), .A2(new_n470), .A3(new_n497), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G141gat), .B1(new_n864), .B2(new_n674), .ZN(new_n865));
  XOR2_X1   g664(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n866));
  NAND3_X1  g665(.A1(new_n853), .A2(new_n677), .A3(new_n691), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT122), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(KEYINPUT122), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n501), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n674), .A2(G141gat), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n865), .B(new_n866), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n853), .A2(new_n863), .A3(new_n871), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT121), .B1(new_n862), .B2(new_n863), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n673), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(G1344gat));
  INV_X1    g680(.A(new_n870), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n208), .A3(new_n646), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G148gat), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n864), .B(new_n875), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n646), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n835), .A2(new_n451), .A3(new_n854), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n860), .A2(new_n861), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n744), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n863), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n884), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n883), .B1(new_n887), .B2(new_n894), .ZN(G1345gat));
  AOI21_X1  g694(.A(G155gat), .B1(new_n882), .B2(new_n706), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n705), .A2(new_n213), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n886), .B2(new_n897), .ZN(G1346gat));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n214), .A3(new_n703), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n886), .A2(new_n703), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n214), .ZN(G1347gat));
  NOR3_X1   g700(.A1(new_n677), .A2(new_n501), .A3(new_n504), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n835), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT124), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n674), .ZN(new_n906));
  INV_X1    g705(.A(new_n903), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n314), .A3(new_n673), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n907), .B2(new_n646), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n744), .A2(new_n315), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n904), .B2(new_n911), .ZN(G1349gat));
  OAI211_X1 g711(.A(new_n907), .B(new_n706), .C1(new_n342), .C2(new_n341), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n905), .A2(new_n705), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n334), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT60), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n917), .B(new_n913), .C1(new_n914), .C2(new_n334), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n907), .A2(new_n340), .A3(new_n703), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT125), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n703), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(G190gat), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT61), .B(new_n340), .C1(new_n904), .C2(new_n703), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  NOR3_X1   g725(.A1(new_n677), .A2(new_n501), .A3(new_n497), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n853), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(G197gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n673), .ZN(new_n930));
  INV_X1    g729(.A(new_n927), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n891), .A2(new_n674), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(new_n929), .ZN(G1352gat));
  INV_X1    g732(.A(G204gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n934), .A3(new_n646), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT62), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n892), .B2(new_n927), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n936), .A2(new_n937), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n928), .A2(new_n298), .A3(new_n706), .ZN(new_n939));
  INV_X1    g738(.A(new_n854), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n696), .B(new_n940), .C1(new_n833), .C2(new_n834), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT57), .B1(new_n859), .B2(new_n451), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n706), .B(new_n927), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n890), .A2(new_n945), .A3(new_n706), .A4(new_n927), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(G211gat), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(KEYINPUT127), .A3(new_n948), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n944), .A2(new_n946), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT127), .B1(new_n947), .B2(new_n948), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n939), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  AOI21_X1  g752(.A(G218gat), .B1(new_n928), .B2(new_n703), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n891), .A2(new_n931), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n560), .A2(new_n297), .A3(new_n296), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(G1355gat));
endmodule


