

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598;

  XNOR2_X1 U325 ( .A(G190GAT), .B(n293), .ZN(G1351GAT) );
  XOR2_X1 U326 ( .A(n581), .B(n580), .Z(n293) );
  XNOR2_X1 U327 ( .A(n316), .B(KEYINPUT74), .ZN(n456) );
  INV_X1 U328 ( .A(n509), .ZN(n466) );
  AND2_X1 U329 ( .A1(n536), .A2(n513), .ZN(n355) );
  XNOR2_X1 U330 ( .A(G176GAT), .B(G64GAT), .ZN(n316) );
  XNOR2_X1 U331 ( .A(n389), .B(n388), .ZN(n477) );
  INV_X1 U332 ( .A(KEYINPUT104), .ZN(n388) );
  NOR2_X1 U333 ( .A1(n387), .A2(n386), .ZN(n389) );
  XNOR2_X1 U334 ( .A(n534), .B(n533), .ZN(n563) );
  XNOR2_X1 U335 ( .A(n328), .B(n327), .ZN(n330) );
  INV_X1 U336 ( .A(n479), .ZN(n465) );
  XOR2_X1 U337 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n294) );
  XNOR2_X1 U338 ( .A(n356), .B(KEYINPUT103), .ZN(n357) );
  XNOR2_X1 U339 ( .A(n340), .B(KEYINPUT88), .ZN(n341) );
  XNOR2_X1 U340 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U341 ( .A(n375), .B(n341), .ZN(n342) );
  XNOR2_X1 U342 ( .A(n462), .B(n348), .ZN(n349) );
  NOR2_X1 U343 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U344 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U345 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U346 ( .A(KEYINPUT26), .B(KEYINPUT102), .ZN(n353) );
  NAND2_X1 U347 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U348 ( .A(n354), .B(n353), .ZN(n582) );
  XNOR2_X1 U349 ( .A(n467), .B(KEYINPUT110), .ZN(n468) );
  NOR2_X1 U350 ( .A1(n570), .A2(n569), .ZN(n579) );
  XOR2_X1 U351 ( .A(n332), .B(n331), .Z(n513) );
  XNOR2_X1 U352 ( .A(n469), .B(G43GAT), .ZN(n470) );
  XNOR2_X1 U353 ( .A(n471), .B(n470), .ZN(G1330GAT) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G127GAT), .Z(n396) );
  XOR2_X1 U355 ( .A(G120GAT), .B(G71GAT), .Z(n455) );
  XNOR2_X1 U356 ( .A(n396), .B(n455), .ZN(n297) );
  XOR2_X1 U357 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n296) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT84), .ZN(n295) );
  XNOR2_X1 U359 ( .A(n296), .B(n295), .ZN(n379) );
  XNOR2_X1 U360 ( .A(n297), .B(n379), .ZN(n303) );
  XOR2_X1 U361 ( .A(G183GAT), .B(KEYINPUT18), .Z(n299) );
  XNOR2_X1 U362 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n324) );
  XOR2_X1 U364 ( .A(G113GAT), .B(n324), .Z(n301) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U366 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U367 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U368 ( .A(KEYINPUT86), .B(G99GAT), .Z(n305) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U371 ( .A(G176GAT), .B(KEYINPUT87), .Z(n307) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n306) );
  XNOR2_X1 U373 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U374 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n570) );
  XOR2_X1 U376 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n313) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U378 ( .A(n313), .B(n312), .ZN(n315) );
  XOR2_X1 U379 ( .A(G218GAT), .B(KEYINPUT90), .Z(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n351) );
  INV_X1 U381 ( .A(n351), .ZN(n332) );
  XOR2_X1 U382 ( .A(G36GAT), .B(G190GAT), .Z(n413) );
  INV_X1 U383 ( .A(n413), .ZN(n317) );
  NAND2_X1 U384 ( .A1(n456), .A2(n317), .ZN(n320) );
  INV_X1 U385 ( .A(n456), .ZN(n318) );
  NAND2_X1 U386 ( .A1(n318), .A2(n413), .ZN(n319) );
  NAND2_X1 U387 ( .A1(n320), .A2(n319), .ZN(n322) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U389 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n323), .B(KEYINPUT100), .ZN(n328) );
  XOR2_X1 U391 ( .A(n324), .B(KEYINPUT79), .Z(n326) );
  INV_X1 U392 ( .A(G92GAT), .ZN(n325) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n433) );
  XNOR2_X1 U394 ( .A(n433), .B(G204GAT), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n331) );
  INV_X1 U396 ( .A(n513), .ZN(n562) );
  XOR2_X1 U397 ( .A(KEYINPUT27), .B(KEYINPUT101), .Z(n333) );
  XNOR2_X1 U398 ( .A(n562), .B(n333), .ZN(n385) );
  XOR2_X1 U399 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n336) );
  XOR2_X1 U400 ( .A(G141GAT), .B(G22GAT), .Z(n445) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(KEYINPUT77), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n334), .B(G162GAT), .ZN(n416) );
  XNOR2_X1 U403 ( .A(n445), .B(n416), .ZN(n335) );
  XOR2_X1 U404 ( .A(n336), .B(n335), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT91), .B(G155GAT), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n294), .B(n337), .ZN(n339) );
  INV_X1 U407 ( .A(KEYINPUT92), .ZN(n338) );
  XNOR2_X1 U408 ( .A(n339), .B(n338), .ZN(n375) );
  XOR2_X1 U409 ( .A(KEYINPUT93), .B(KEYINPUT22), .Z(n340) );
  XNOR2_X1 U410 ( .A(n343), .B(n342), .ZN(n350) );
  XNOR2_X1 U411 ( .A(G148GAT), .B(KEYINPUT70), .ZN(n344) );
  XNOR2_X1 U412 ( .A(n344), .B(KEYINPUT71), .ZN(n345) );
  XOR2_X1 U413 ( .A(n345), .B(G204GAT), .Z(n347) );
  XNOR2_X1 U414 ( .A(G78GAT), .B(G106GAT), .ZN(n346) );
  XNOR2_X1 U415 ( .A(n347), .B(n346), .ZN(n462) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n567) );
  NAND2_X1 U418 ( .A1(n567), .A2(n570), .ZN(n354) );
  NOR2_X1 U419 ( .A1(n385), .A2(n582), .ZN(n360) );
  INV_X1 U420 ( .A(n570), .ZN(n536) );
  OR2_X1 U421 ( .A1(n567), .A2(n355), .ZN(n358) );
  INV_X1 U422 ( .A(KEYINPUT25), .ZN(n356) );
  NOR2_X1 U423 ( .A1(n360), .A2(n359), .ZN(n384) );
  XOR2_X1 U424 ( .A(G113GAT), .B(G1GAT), .Z(n435) );
  XOR2_X1 U425 ( .A(G85GAT), .B(G162GAT), .Z(n362) );
  XNOR2_X1 U426 ( .A(G29GAT), .B(G141GAT), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U428 ( .A(n435), .B(n363), .Z(n365) );
  NAND2_X1 U429 ( .A1(G225GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n383) );
  XOR2_X1 U431 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n367) );
  XNOR2_X1 U432 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U434 ( .A(G57GAT), .B(G148GAT), .Z(n369) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G120GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U438 ( .A(KEYINPUT4), .B(KEYINPUT96), .Z(n373) );
  XNOR2_X1 U439 ( .A(KEYINPUT98), .B(KEYINPUT97), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U443 ( .A(n378), .B(KEYINPUT99), .Z(n381) );
  XNOR2_X1 U444 ( .A(n379), .B(KEYINPUT94), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U446 ( .A(n383), .B(n382), .Z(n565) );
  INV_X1 U447 ( .A(n565), .ZN(n510) );
  NOR2_X1 U448 ( .A1(n384), .A2(n510), .ZN(n387) );
  NOR2_X1 U449 ( .A1(n565), .A2(n385), .ZN(n549) );
  XOR2_X1 U450 ( .A(KEYINPUT28), .B(n567), .Z(n493) );
  NAND2_X1 U451 ( .A1(n549), .A2(n493), .ZN(n535) );
  NOR2_X1 U452 ( .A1(n535), .A2(n536), .ZN(n386) );
  XOR2_X1 U453 ( .A(G155GAT), .B(G211GAT), .Z(n391) );
  XNOR2_X1 U454 ( .A(G22GAT), .B(G78GAT), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U456 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n393) );
  XNOR2_X1 U457 ( .A(G183GAT), .B(G71GAT), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U459 ( .A(n395), .B(n394), .Z(n401) );
  XOR2_X1 U460 ( .A(G57GAT), .B(KEYINPUT13), .Z(n452) );
  XOR2_X1 U461 ( .A(n396), .B(n452), .Z(n398) );
  NAND2_X1 U462 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U464 ( .A(G8GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U466 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n403) );
  XNOR2_X1 U467 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U469 ( .A(KEYINPUT80), .B(KEYINPUT83), .Z(n405) );
  XNOR2_X1 U470 ( .A(G1GAT), .B(KEYINPUT14), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U472 ( .A(n407), .B(n406), .Z(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n556) );
  INV_X1 U474 ( .A(n556), .ZN(n592) );
  XOR2_X1 U475 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n411) );
  XNOR2_X1 U476 ( .A(G218GAT), .B(KEYINPUT78), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U478 ( .A(n412), .B(KEYINPUT10), .Z(n415) );
  XNOR2_X1 U479 ( .A(G106GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U481 ( .A(n416), .B(G134GAT), .Z(n418) );
  NAND2_X1 U482 ( .A1(G232GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U484 ( .A(n420), .B(n419), .Z(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT67), .B(KEYINPUT8), .Z(n422) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G29GAT), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U488 ( .A(KEYINPUT7), .B(n423), .Z(n436) );
  XOR2_X1 U489 ( .A(KEYINPUT72), .B(G92GAT), .Z(n425) );
  XNOR2_X1 U490 ( .A(G99GAT), .B(KEYINPUT73), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U492 ( .A(G85GAT), .B(n426), .Z(n461) );
  XNOR2_X1 U493 ( .A(n436), .B(n461), .ZN(n427) );
  XNOR2_X1 U494 ( .A(n428), .B(n427), .ZN(n578) );
  XOR2_X1 U495 ( .A(n578), .B(KEYINPUT36), .Z(n596) );
  NOR2_X1 U496 ( .A1(n592), .A2(n596), .ZN(n429) );
  NAND2_X1 U497 ( .A1(n477), .A2(n429), .ZN(n430) );
  XOR2_X1 U498 ( .A(n430), .B(KEYINPUT37), .Z(n509) );
  XOR2_X1 U499 ( .A(G15GAT), .B(G197GAT), .Z(n432) );
  XNOR2_X1 U500 ( .A(G36GAT), .B(G50GAT), .ZN(n431) );
  XNOR2_X1 U501 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U502 ( .A(n434), .B(n433), .Z(n438) );
  XNOR2_X1 U503 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U504 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U505 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n440) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U507 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U508 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U509 ( .A(KEYINPUT29), .B(KEYINPUT64), .Z(n444) );
  XNOR2_X1 U510 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n443) );
  XNOR2_X1 U511 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n550) );
  INV_X1 U514 ( .A(n550), .ZN(n584) );
  XOR2_X1 U515 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n450) );
  XNOR2_X1 U516 ( .A(KEYINPUT69), .B(KEYINPUT75), .ZN(n449) );
  XNOR2_X1 U517 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U518 ( .A(n451), .B(KEYINPUT33), .Z(n454) );
  XNOR2_X1 U519 ( .A(n452), .B(KEYINPUT32), .ZN(n453) );
  XNOR2_X1 U520 ( .A(n454), .B(n453), .ZN(n460) );
  XOR2_X1 U521 ( .A(n456), .B(n455), .Z(n458) );
  NAND2_X1 U522 ( .A1(G230GAT), .A2(G233GAT), .ZN(n457) );
  XNOR2_X1 U523 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U524 ( .A(n460), .B(n459), .Z(n464) );
  XNOR2_X1 U525 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(n588) );
  NAND2_X1 U527 ( .A1(n584), .A2(n588), .ZN(n479) );
  XNOR2_X1 U528 ( .A(KEYINPUT38), .B(n468), .ZN(n492) );
  NOR2_X1 U529 ( .A1(n570), .A2(n492), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n565), .A2(n492), .ZN(n475) );
  XNOR2_X1 U532 ( .A(KEYINPUT109), .B(KEYINPUT39), .ZN(n473) );
  INV_X1 U533 ( .A(G29GAT), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(G1328GAT) );
  NOR2_X1 U536 ( .A1(n578), .A2(n556), .ZN(n476) );
  XNOR2_X1 U537 ( .A(KEYINPUT16), .B(n476), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n478), .A2(n477), .ZN(n498) );
  NOR2_X1 U539 ( .A1(n479), .A2(n498), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n510), .A2(n488), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT106), .Z(n481) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(KEYINPUT105), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n488), .A2(n513), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT107), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U548 ( .A1(n488), .A2(n536), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U550 ( .A(G15GAT), .B(n487), .Z(G1326GAT) );
  INV_X1 U551 ( .A(n493), .ZN(n517) );
  NAND2_X1 U552 ( .A1(n488), .A2(n517), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n489), .B(KEYINPUT108), .ZN(n490) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(n490), .ZN(G1327GAT) );
  NOR2_X1 U555 ( .A1(n562), .A2(n492), .ZN(n491) );
  XOR2_X1 U556 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  NOR2_X1 U557 ( .A1(n493), .A2(n492), .ZN(n495) );
  INV_X1 U558 ( .A(KEYINPUT112), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n496), .ZN(G1331GAT) );
  XOR2_X2 U561 ( .A(KEYINPUT41), .B(n588), .Z(n572) );
  NOR2_X1 U562 ( .A1(n584), .A2(n572), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n497), .B(KEYINPUT113), .ZN(n508) );
  NOR2_X1 U564 ( .A1(n498), .A2(n508), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n499), .B(KEYINPUT114), .ZN(n504) );
  NAND2_X1 U566 ( .A1(n504), .A2(n510), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n513), .A2(n504), .ZN(n502) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n504), .A2(n536), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT43), .B(KEYINPUT115), .Z(n506) );
  NAND2_X1 U574 ( .A1(n517), .A2(n504), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NOR2_X1 U577 ( .A1(n509), .A2(n508), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n518), .A2(n510), .ZN(n511) );
  XNOR2_X1 U579 ( .A(KEYINPUT116), .B(n511), .ZN(n512) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n518), .A2(n513), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n514), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT117), .Z(n516) );
  NAND2_X1 U584 ( .A1(n518), .A2(n536), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n516), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT118), .Z(n520) );
  NAND2_X1 U587 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n521), .Z(G1339GAT) );
  XNOR2_X1 U590 ( .A(KEYINPUT121), .B(KEYINPUT48), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n550), .A2(n588), .ZN(n524) );
  NOR2_X1 U592 ( .A1(n596), .A2(n556), .ZN(n522) );
  XOR2_X1 U593 ( .A(KEYINPUT45), .B(n522), .Z(n523) );
  NOR2_X1 U594 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U595 ( .A(KEYINPUT120), .B(n525), .Z(n532) );
  NOR2_X1 U596 ( .A1(n550), .A2(n572), .ZN(n526) );
  XNOR2_X1 U597 ( .A(n526), .B(KEYINPUT46), .ZN(n527) );
  NOR2_X1 U598 ( .A1(n592), .A2(n527), .ZN(n528) );
  XNOR2_X1 U599 ( .A(n528), .B(KEYINPUT119), .ZN(n529) );
  NOR2_X1 U600 ( .A1(n578), .A2(n529), .ZN(n530) );
  XNOR2_X1 U601 ( .A(KEYINPUT47), .B(n530), .ZN(n531) );
  NAND2_X1 U602 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U603 ( .A1(n563), .A2(n535), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n550), .A2(n545), .ZN(n538) );
  XOR2_X1 U606 ( .A(G113GAT), .B(n538), .Z(G1340GAT) );
  NOR2_X1 U607 ( .A1(n572), .A2(n545), .ZN(n540) );
  XNOR2_X1 U608 ( .A(KEYINPUT122), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NOR2_X1 U611 ( .A1(n556), .A2(n545), .ZN(n543) );
  XNOR2_X1 U612 ( .A(KEYINPUT123), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  INV_X1 U615 ( .A(n578), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n559), .A2(n545), .ZN(n547) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U618 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n563), .A2(n582), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n549), .A2(n548), .ZN(n558) );
  NOR2_X1 U621 ( .A1(n550), .A2(n558), .ZN(n551) );
  XOR2_X1 U622 ( .A(KEYINPUT124), .B(n551), .Z(n552) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U624 ( .A1(n572), .A2(n558), .ZN(n554) );
  XNOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U626 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U628 ( .A1(n556), .A2(n558), .ZN(n557) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U630 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(KEYINPUT125), .ZN(n560) );
  XNOR2_X1 U632 ( .A(n561), .B(n560), .ZN(G1347GAT) );
  XNOR2_X1 U633 ( .A(KEYINPUT54), .B(n564), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n583) );
  NOR2_X1 U635 ( .A1(n567), .A2(n583), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT55), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n579), .A2(n584), .ZN(n571) );
  XNOR2_X1 U638 ( .A(G169GAT), .B(n571), .ZN(G1348GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n575) );
  INV_X1 U640 ( .A(n572), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n579), .A2(n573), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(G176GAT), .B(n576), .ZN(G1349GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n592), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n581) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n586) );
  NOR2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n593) );
  NAND2_X1 U650 ( .A1(n593), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(n587), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n590) );
  INV_X1 U654 ( .A(n593), .ZN(n595) );
  OR2_X1 U655 ( .A1(n595), .A2(n588), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U657 ( .A(G204GAT), .B(n591), .Z(G1353GAT) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n594), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(KEYINPUT62), .B(n597), .Z(n598) );
  XNOR2_X1 U662 ( .A(G218GAT), .B(n598), .ZN(G1355GAT) );
endmodule

