//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G125), .ZN(new_n460));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT67), .Z(new_n483));
  AOI211_X1 g058(.A(new_n476), .B(new_n483), .C1(G136), .C2(new_n467), .ZN(G162));
  NAND2_X1  g059(.A1(G126), .A2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n461), .B2(new_n462), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n480), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n477), .C2(new_n478), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n480), .C1(new_n477), .C2(new_n478), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n500), .A3(G138), .A4(new_n480), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n490), .A2(new_n496), .B1(new_n498), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT69), .A3(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(G88), .B1(G50), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n506), .A2(KEYINPUT69), .A3(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n506), .B2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT70), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n513), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n510), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(new_n511), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n529), .B(new_n530), .C1(new_n533), .C2(KEYINPUT71), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n516), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n508), .A2(new_n509), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n511), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n516), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT72), .B(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n539), .A2(new_n546), .B1(new_n547), .B2(new_n511), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n522), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n508), .A2(G65), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n560), .A2(KEYINPUT73), .A3(new_n555), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(G651), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n511), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n509), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  AOI22_X1  g141(.A1(G91), .A2(new_n510), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  XNOR2_X1  g144(.A(G171), .B(new_n569), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n526), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n513), .A2(new_n517), .A3(KEYINPUT75), .A4(new_n525), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(G303));
  NAND2_X1  g150(.A1(new_n510), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n512), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  OAI211_X1 g154(.A(G61), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n508), .A2(KEYINPUT76), .A3(G61), .ZN(new_n583));
  AND2_X1   g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n539), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n510), .A2(G85), .B1(G47), .B2(new_n512), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT78), .Z(new_n594));
  AOI22_X1  g169(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n516), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(new_n510), .A2(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  MUX2_X1   g181(.A(new_n606), .B(G301), .S(G868), .Z(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT79), .Z(G284));
  XNOR2_X1  g183(.A(new_n607), .B(KEYINPUT80), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(G868), .B2(new_n611), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(G868), .B2(new_n611), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n619), .B(new_n620), .C1(G868), .C2(new_n549), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n499), .A2(new_n470), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n481), .A2(G123), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT82), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G2105), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(G135), .B2(new_n467), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n625), .A2(new_n626), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(G2096), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n627), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n642), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT83), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  XOR2_X1   g236(.A(new_n659), .B(KEYINPUT17), .Z(new_n662));
  INV_X1    g237(.A(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n664), .B1(new_n666), .B2(KEYINPUT84), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(KEYINPUT84), .B2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n657), .A2(new_n662), .A3(new_n663), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n661), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n626), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT85), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT86), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n690), .B2(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G29), .A2(G35), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G162), .B2(G29), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT29), .ZN(new_n699));
  INV_X1    g274(.A(G2090), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G20), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT23), .Z(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G299), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1956), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G26), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n481), .A2(G128), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  NOR2_X1   g286(.A1(G104), .A2(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT91), .ZN(new_n713));
  INV_X1    g288(.A(G116), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n469), .B1(new_n714), .B2(G2105), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n713), .A2(new_n715), .B1(G140), .B2(new_n467), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT92), .B(G2067), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n702), .A2(G19), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n549), .B2(new_n702), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT89), .B(G1341), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G4), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n614), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1348), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n701), .A2(new_n706), .A3(new_n725), .A4(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT97), .B1(G16), .B2(G21), .ZN(new_n731));
  NAND2_X1  g306(.A1(G168), .A2(G16), .ZN(new_n732));
  MUX2_X1   g307(.A(KEYINPUT97), .B(new_n731), .S(new_n732), .Z(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT98), .Z(new_n736));
  OR2_X1    g311(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  INV_X1    g312(.A(G11), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT31), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G28), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n707), .B1(new_n741), .B2(G28), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n739), .B(new_n740), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n634), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT24), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n707), .B1(new_n747), .B2(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n747), .B2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G160), .B2(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2084), .ZN(new_n751));
  INV_X1    g326(.A(G2072), .ZN(new_n752));
  OR2_X1    g327(.A1(G29), .A2(G33), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT25), .ZN(new_n756));
  NAND2_X1  g331(.A1(G115), .A2(G2104), .ZN(new_n757));
  INV_X1    g332(.A(G127), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n479), .B2(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n759), .A2(G2105), .B1(G139), .B2(new_n467), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(new_n707), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n746), .B(new_n751), .C1(new_n752), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G5), .A2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT99), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G171), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1961), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n707), .A2(G27), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT101), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n490), .A2(new_n496), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n498), .A2(new_n501), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n769), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n763), .A2(new_n767), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G32), .ZN(new_n777));
  AOI21_X1  g352(.A(KEYINPUT96), .B1(new_n707), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n470), .A2(G105), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT95), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n467), .A2(G141), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n481), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT26), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(KEYINPUT26), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  MUX2_X1   g365(.A(KEYINPUT96), .B(new_n778), .S(new_n790), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT27), .B(G1996), .Z(new_n792));
  OR2_X1    g367(.A1(new_n750), .A2(G2084), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n792), .B1(KEYINPUT100), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(KEYINPUT100), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n794), .B(new_n795), .C1(new_n792), .C2(new_n791), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n762), .A2(new_n752), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n736), .A2(new_n737), .A3(new_n776), .A4(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT102), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT102), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n730), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n481), .A2(G119), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT87), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(G107), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G2105), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G131), .B2(new_n467), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT88), .ZN(new_n812));
  MUX2_X1   g387(.A(G25), .B(new_n812), .S(G29), .Z(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NOR2_X1   g390(.A1(G6), .A2(G16), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n590), .B1(new_n586), .B2(G651), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(G166), .A2(G16), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G16), .B2(G22), .ZN(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n702), .A2(G23), .ZN(new_n826));
  INV_X1    g401(.A(G288), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n702), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT33), .B(G1976), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n818), .A2(new_n819), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OR3_X1    g407(.A1(new_n825), .A2(KEYINPUT34), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(KEYINPUT34), .B1(new_n825), .B2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n702), .A2(G24), .ZN(new_n835));
  INV_X1    g410(.A(G290), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(new_n702), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n686), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n815), .A2(new_n833), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT36), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n803), .A2(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  NOR2_X1   g417(.A1(new_n606), .A2(new_n615), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n516), .ZN(new_n847));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n539), .A2(new_n848), .B1(new_n849), .B2(new_n511), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n549), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n549), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n845), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT104), .ZN(new_n860));
  OAI21_X1  g435(.A(G860), .B1(new_n847), .B2(new_n850), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n634), .B(G160), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G162), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n811), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n624), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n481), .A2(G130), .ZN(new_n871));
  OR2_X1    g446(.A1(G106), .A2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n872), .B(G2104), .C1(G118), .C2(new_n480), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(G142), .B2(new_n467), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n870), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n761), .A2(KEYINPUT105), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n717), .Z(new_n878));
  NOR2_X1   g453(.A1(new_n486), .A2(new_n489), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n771), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n789), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n789), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n876), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT107), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n883), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n876), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n884), .A2(new_n885), .ZN(new_n893));
  INV_X1    g468(.A(new_n876), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n867), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n866), .B1(new_n893), .B2(new_n894), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n897), .B2(new_n886), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n864), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n887), .A2(new_n891), .B1(new_n894), .B2(new_n893), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n898), .B(KEYINPUT40), .C1(new_n901), .C2(new_n867), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(G395));
  XNOR2_X1  g478(.A(new_n617), .B(new_n854), .ZN(new_n904));
  OR2_X1    g479(.A1(G299), .A2(KEYINPUT108), .ZN(new_n905));
  NAND2_X1  g480(.A1(G299), .A2(KEYINPUT108), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n614), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n606), .A2(KEYINPUT108), .A3(G299), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(KEYINPUT41), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n904), .A2(new_n909), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n915), .A2(KEYINPUT42), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G288), .B(KEYINPUT110), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n526), .B(new_n817), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n919), .B(new_n920), .Z(new_n921));
  OAI21_X1  g496(.A(KEYINPUT42), .B1(new_n915), .B2(new_n916), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n917), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(G868), .B2(new_n851), .ZN(G295));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n851), .ZN(G331));
  XNOR2_X1  g502(.A(G171), .B(KEYINPUT74), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(G168), .ZN(new_n929));
  NOR2_X1   g504(.A1(G168), .A2(G171), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n929), .B2(new_n931), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n854), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  NOR2_X1   g512(.A1(G301), .A2(G286), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT111), .B1(new_n938), .B2(new_n930), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n933), .A3(new_n855), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n939), .A2(new_n933), .A3(KEYINPUT112), .A4(new_n855), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n913), .A3(new_n914), .A4(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n936), .A2(new_n908), .A3(new_n907), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n945), .B2(new_n921), .ZN(new_n946));
  INV_X1    g521(.A(new_n921), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT43), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n909), .B1(new_n941), .B2(new_n942), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n936), .A2(new_n940), .B1(new_n910), .B2(new_n912), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n921), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  AND4_X1   g528(.A1(KEYINPUT43), .A2(new_n952), .A3(new_n953), .A4(new_n948), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT44), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n946), .B2(new_n948), .ZN(new_n958));
  AND4_X1   g533(.A1(new_n957), .A2(new_n952), .A3(new_n953), .A4(new_n948), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n960), .ZN(G397));
  AOI21_X1  g536(.A(G1384), .B1(new_n771), .B2(new_n879), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n465), .A2(G40), .A3(new_n471), .A4(new_n468), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G2067), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n717), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n789), .B(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n811), .B(new_n814), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n836), .A2(new_n686), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n836), .A2(new_n686), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT113), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n968), .B1(new_n976), .B2(KEYINPUT113), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n966), .A2(new_n962), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G8), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1976), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n827), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(G305), .A2(G1981), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n817), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n584), .B1(new_n580), .B2(new_n581), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n516), .B1(new_n991), .B2(new_n583), .ZN(new_n992));
  NOR4_X1   g567(.A1(new_n992), .A2(KEYINPUT117), .A3(new_n590), .A4(G1981), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n983), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT49), .B(new_n987), .C1(new_n990), .C2(new_n993), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n986), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n990), .A2(new_n993), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n984), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n982), .B(G8), .C1(new_n985), .C2(G288), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT52), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n827), .B2(G1976), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1002), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n996), .B2(new_n997), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n770), .B2(new_n771), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT114), .B(new_n964), .C1(G164), .C2(G1384), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n965), .B1(new_n962), .B2(KEYINPUT45), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1007), .B1(new_n1013), .B2(new_n823), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1007), .A3(new_n823), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n965), .B1(new_n962), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(new_n1021), .B2(G2090), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1019), .A2(KEYINPUT116), .A3(new_n1020), .A4(new_n700), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1015), .A2(new_n1016), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n573), .A2(G8), .A3(new_n574), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n573), .A2(KEYINPUT55), .A3(G8), .A4(new_n574), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1006), .A2(new_n1024), .A3(G8), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1000), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1000), .B2(new_n1030), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n772), .A2(KEYINPUT45), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n491), .A2(new_n494), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n498), .B2(new_n501), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n964), .B1(new_n1038), .B2(G1384), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1039), .A3(new_n966), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n734), .ZN(new_n1041));
  INV_X1    g616(.A(G2084), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1019), .A2(new_n1042), .A3(new_n1020), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(G8), .A3(G286), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(G168), .A3(new_n1043), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(KEYINPUT122), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1046), .A2(KEYINPUT51), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1045), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT62), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1010), .A2(new_n774), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  INV_X1    g629(.A(G1961), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1053), .A2(new_n1054), .B1(new_n1055), .B2(new_n1021), .ZN(new_n1056));
  OR3_X1    g631(.A1(new_n1040), .A2(new_n1054), .A3(G2078), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1045), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1052), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n561), .A2(G651), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT73), .B1(new_n560), .B2(new_n555), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n567), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1062), .B1(new_n562), .B2(new_n567), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1009), .A2(new_n1018), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT50), .B1(new_n1038), .B2(G1384), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n966), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1956), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n982), .A2(G2067), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1348), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n614), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1068), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1076), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n614), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1085), .B2(new_n614), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1078), .A2(new_n1084), .A3(new_n1077), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1089), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n880), .A2(new_n1018), .A3(new_n1035), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n966), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1018), .B1(new_n772), .B2(new_n1035), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n728), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n982), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n969), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT60), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT121), .B1(new_n1098), .B2(new_n606), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1085), .A2(new_n1086), .A3(new_n614), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1091), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1090), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1067), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1073), .A2(new_n1075), .B1(new_n1103), .B2(new_n1065), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT61), .B1(new_n1076), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1082), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT58), .B(G1341), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1013), .A2(G1996), .B1(new_n1096), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n549), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1110), .B(new_n549), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1105), .A2(new_n1108), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1083), .B1(new_n1102), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1054), .B(G2078), .C1(new_n965), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n966), .A2(KEYINPUT123), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1039), .A4(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1056), .A2(G301), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1119), .B1(new_n1125), .B2(new_n1058), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1056), .A2(G301), .A3(new_n1057), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1021), .A2(new_n1055), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1124), .ZN(new_n1130));
  INV_X1    g705(.A(G171), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1127), .B(KEYINPUT54), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1126), .A2(new_n1132), .A3(new_n1051), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1061), .B1(new_n1118), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1016), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1135));
  OAI211_X1 g710(.A(G8), .B(new_n1029), .C1(new_n1135), .C2(new_n1014), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1071), .A2(G2090), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n823), .B2(new_n1013), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1027), .B(new_n1028), .C1(new_n1138), .C2(new_n1047), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1136), .A2(new_n1139), .A3(new_n1006), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1034), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1024), .A2(G8), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1047), .B(G286), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1144), .A2(KEYINPUT63), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1143), .A2(new_n1006), .A3(new_n1136), .A4(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1136), .A2(new_n1139), .A3(new_n1006), .A4(new_n1144), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n981), .B1(new_n1141), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n717), .A2(G2067), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n972), .A2(new_n968), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n812), .A2(new_n814), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n967), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1159), .B2(new_n1158), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT46), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n970), .B(new_n789), .C1(new_n1162), .C2(G1996), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n968), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n967), .B2(G1996), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT125), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT47), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT48), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n977), .A2(new_n1169), .A3(new_n967), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1169), .B1(new_n977), .B2(new_n967), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n974), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1161), .B(new_n1168), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT126), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT127), .B1(new_n1154), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1099), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1089), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1083), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1133), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1061), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1140), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1034), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n1153), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n981), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1173), .B(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1175), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g768(.A(G319), .B1(new_n652), .B2(new_n653), .ZN(new_n1195));
  NOR2_X1   g769(.A1(G227), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g770(.A1(new_n694), .A2(new_n695), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1197), .B1(new_n896), .B2(new_n899), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n959), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1199), .ZN(G308));
  OAI221_X1 g774(.A(new_n1197), .B1(new_n896), .B2(new_n899), .C1(new_n958), .C2(new_n959), .ZN(G225));
endmodule


