//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT1), .A3(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(new_n198), .C1(G128), .C2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n194), .A2(new_n196), .A3(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n199), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G224), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G953), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n209), .B(KEYINPUT76), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n207), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G110), .B(G122), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n214), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G101), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n215), .A2(new_n218), .A3(new_n222), .A4(new_n219), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT4), .B(new_n221), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G116), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT65), .B1(new_n230), .B2(G119), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(G119), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT2), .A2(G113), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n233), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n215), .A2(new_n218), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n222), .A4(new_n219), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n217), .A2(G104), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n219), .A2(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n243), .A2(new_n244), .B1(G101), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n236), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n233), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT5), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n232), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(G113), .B(new_n251), .C1(new_n233), .C2(new_n250), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  AOI211_X1 g067(.A(KEYINPUT6), .B(new_n213), .C1(new_n240), .C2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n240), .A2(new_n253), .A3(new_n213), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT75), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n240), .A2(new_n253), .A3(new_n257), .A4(new_n213), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n213), .B1(new_n240), .B2(new_n253), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n212), .B(new_n254), .C1(new_n259), .C2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  INV_X1    g078(.A(new_n259), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n213), .B(KEYINPUT8), .Z(new_n267));
  NAND2_X1  g081(.A1(new_n246), .A2(G101), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(new_n224), .B2(new_n225), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n249), .A2(new_n252), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(new_n253), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n206), .B(new_n274), .C1(G125), .C2(new_n200), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT7), .B1(new_n208), .B2(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n201), .A2(new_n206), .A3(new_n278), .A4(new_n274), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n266), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n267), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n269), .A2(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n243), .A2(new_n244), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n284), .A2(new_n268), .B1(new_n249), .B2(new_n252), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT78), .A3(new_n277), .A4(new_n279), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n264), .B1(new_n265), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n190), .B1(new_n263), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n281), .A2(new_n287), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n291), .B2(new_n259), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n259), .A2(new_n262), .ZN(new_n293));
  INV_X1    g107(.A(new_n254), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n211), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n295), .A3(new_n189), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n188), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT9), .B(G234), .Z(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G221), .B1(new_n299), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  XNOR2_X1  g115(.A(G110), .B(G140), .ZN(new_n302));
  INV_X1    g116(.A(G953), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(G227), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n302), .B(new_n304), .Z(new_n305));
  INV_X1    g119(.A(KEYINPUT11), .ZN(new_n306));
  INV_X1    g120(.A(G134), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(G137), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(G137), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT11), .A3(G134), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  INV_X1    g127(.A(G131), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n308), .A2(new_n311), .A3(new_n314), .A4(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n205), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n226), .A2(new_n239), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n268), .B(new_n200), .C1(new_n224), .C2(new_n225), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT73), .B1(new_n319), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n319), .B2(new_n320), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n247), .A2(KEYINPUT74), .A3(KEYINPUT10), .A4(new_n200), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n316), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n320), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n316), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n318), .A3(new_n335), .A4(new_n327), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n305), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n319), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n200), .B1(new_n284), .B2(new_n268), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n316), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(KEYINPUT12), .B(new_n316), .C1(new_n338), .C2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n336), .A2(new_n344), .A3(new_n305), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n301), .B(new_n264), .C1(new_n337), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(G469), .A2(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(new_n305), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n329), .A2(new_n336), .A3(new_n305), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(G469), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n297), .A2(new_n300), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G125), .B(G140), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n193), .ZN(new_n356));
  AND2_X1   g170(.A1(KEYINPUT66), .A2(G237), .ZN(new_n357));
  NOR2_X1   g171(.A1(KEYINPUT66), .A2(G237), .ZN(new_n358));
  OAI211_X1 g172(.A(G214), .B(new_n303), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n195), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT66), .B(G237), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(G143), .A3(G214), .A4(new_n303), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n314), .B1(new_n360), .B2(new_n362), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n365), .A2(KEYINPUT79), .A3(KEYINPUT18), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT79), .B1(new_n365), .B2(KEYINPUT18), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n356), .B(new_n364), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G125), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n369), .A2(KEYINPUT16), .A3(G140), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(G146), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(G146), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n365), .A2(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n360), .A2(new_n362), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n360), .A2(new_n362), .A3(new_n314), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n374), .B(new_n375), .C1(new_n379), .C2(KEYINPUT17), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n368), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n368), .A2(new_n380), .A3(new_n383), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G475), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G478), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(KEYINPUT15), .ZN(new_n391));
  INV_X1    g205(.A(G122), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT83), .B1(new_n392), .B2(G116), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n230), .A3(G122), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(G116), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n217), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT85), .ZN(new_n399));
  XNOR2_X1  g213(.A(G128), .B(G143), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n307), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n396), .A2(KEYINPUT14), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n397), .B1(new_n396), .B2(KEYINPUT14), .ZN(new_n403));
  OAI21_X1  g217(.A(G107), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n396), .A2(new_n397), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G107), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n398), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT13), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n191), .B2(G143), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n195), .A2(KEYINPUT13), .A3(G128), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n410), .B(new_n411), .C1(G128), .C2(new_n195), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT84), .A3(G134), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n400), .A2(new_n307), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(G134), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n408), .A2(new_n413), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G217), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n299), .A2(new_n419), .A3(G953), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n405), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n405), .B2(new_n418), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n391), .B1(new_n424), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n423), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  INV_X1    g241(.A(new_n391), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n264), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(G234), .A2(G237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(G952), .A3(new_n303), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT21), .B(G898), .Z(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(G902), .A3(G953), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n386), .ZN(new_n436));
  INV_X1    g250(.A(new_n372), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n355), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n355), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n355), .B2(new_n438), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(new_n440), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n379), .B(new_n437), .C1(new_n445), .C2(G146), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n368), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n383), .B1(new_n447), .B2(KEYINPUT82), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n368), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n436), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT20), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n368), .A2(new_n449), .A3(new_n446), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n449), .B1(new_n368), .B2(new_n446), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n456), .A2(new_n457), .A3(new_n383), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n455), .B(new_n452), .C1(new_n458), .C2(new_n436), .ZN(new_n459));
  AOI211_X1 g273(.A(new_n389), .B(new_n435), .C1(new_n454), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT86), .B1(new_n354), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n300), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n352), .A2(new_n347), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n346), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n297), .A4(new_n460), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n316), .A2(new_n317), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n307), .A2(G137), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT64), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n309), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(G131), .C1(new_n472), .C2(new_n469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n200), .A2(new_n315), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n237), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(G210), .B(new_n303), .C1(new_n357), .C2(new_n358), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT27), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n361), .A2(new_n478), .A3(G210), .A4(new_n303), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT26), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n477), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n222), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n479), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT26), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(G101), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n468), .A2(new_n474), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n238), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT67), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n475), .A2(new_n483), .A3(new_n487), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n489), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT31), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n468), .A2(new_n237), .A3(new_n474), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n237), .B1(new_n468), .B2(new_n474), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT28), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT28), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n475), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n483), .A2(new_n487), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT31), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n489), .A2(new_n507), .A3(new_n494), .A4(new_n496), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n498), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G472), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n264), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT32), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n505), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n501), .A2(new_n514), .A3(KEYINPUT29), .A4(new_n503), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n501), .A2(new_n503), .A3(new_n514), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n514), .B1(new_n494), .B2(new_n475), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n264), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G472), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT68), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n509), .A2(KEYINPUT32), .A3(new_n510), .A4(new_n264), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT68), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n524), .A3(G472), .ZN(new_n525));
  AND4_X1   g339(.A1(new_n513), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n419), .B1(G234), .B2(new_n264), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n372), .B1(new_n193), .B2(new_n355), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT23), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n228), .B2(G128), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n228), .A2(G128), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n534));
  OR3_X1    g348(.A1(new_n533), .A2(new_n534), .A3(G110), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n533), .B2(G110), .ZN(new_n536));
  XNOR2_X1  g350(.A(G119), .B(G128), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT24), .B(G110), .Z(new_n538));
  OAI211_X1 g352(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n528), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n537), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n541), .A2(KEYINPUT69), .B1(G110), .B2(new_n533), .ZN(new_n542));
  OAI221_X1 g356(.A(new_n542), .B1(KEYINPUT69), .B2(new_n541), .C1(new_n372), .C2(new_n373), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n303), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT22), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(G137), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n540), .A2(new_n543), .A3(new_n547), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n264), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT25), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n551), .A2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n527), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n527), .A2(G902), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n549), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n526), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n462), .A2(new_n467), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G101), .ZN(G3));
  NAND2_X1  g376(.A1(new_n454), .A2(new_n459), .ZN(new_n563));
  INV_X1    g377(.A(new_n389), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT88), .B(KEYINPUT33), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n427), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n426), .A2(new_n421), .B1(new_n568), .B2(KEYINPUT33), .ZN(new_n569));
  OAI21_X1  g383(.A(G478), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n390), .A2(new_n264), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n427), .A2(new_n390), .A3(new_n264), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n297), .A2(new_n565), .A3(new_n434), .A4(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT87), .ZN(new_n578));
  INV_X1    g392(.A(new_n559), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n509), .A2(new_n264), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n511), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n353), .A2(new_n300), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n511), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(new_n559), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n465), .A2(new_n586), .A3(KEYINPUT87), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n577), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT34), .B(G104), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT89), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n588), .B(new_n590), .ZN(G6));
  NAND2_X1  g405(.A1(new_n297), .A2(new_n434), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT90), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n454), .A2(new_n459), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n425), .A2(new_n429), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n389), .ZN(new_n597));
  OAI211_X1 g411(.A(KEYINPUT90), .B(KEYINPUT20), .C1(new_n451), .C2(new_n453), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n584), .A3(new_n587), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  INV_X1    g417(.A(KEYINPUT91), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n540), .A2(new_n604), .A3(new_n543), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n540), .B2(new_n543), .ZN(new_n609));
  OR3_X1    g423(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n606), .B2(new_n609), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n557), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n556), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n614), .A2(new_n511), .A3(new_n581), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n462), .A2(new_n467), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT37), .B(G110), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G12));
  NAND2_X1  g432(.A1(new_n290), .A2(new_n296), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n187), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n583), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n513), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n614), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n433), .A2(G900), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n431), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n594), .A2(new_n597), .A3(new_n598), .A4(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n621), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G128), .ZN(G30));
  XNOR2_X1  g443(.A(new_n625), .B(KEYINPUT93), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT39), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n465), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT40), .Z(new_n633));
  XOR2_X1   g447(.A(new_n619), .B(KEYINPUT38), .Z(new_n634));
  AOI21_X1  g448(.A(new_n389), .B1(new_n454), .B2(new_n459), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(new_n188), .A3(new_n596), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n634), .A2(new_n614), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n505), .B1(new_n499), .B2(new_n500), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n497), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(G472), .B1(new_n640), .B2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n513), .A2(new_n523), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT92), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n633), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT94), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G143), .ZN(G45));
  INV_X1    g461(.A(new_n625), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n635), .A2(new_n574), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n621), .A2(new_n623), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G146), .ZN(G48));
  OAI21_X1  g465(.A(new_n264), .B1(new_n337), .B2(new_n345), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G469), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n300), .A3(new_n346), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n526), .A2(new_n559), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT95), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n577), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n653), .A2(new_n300), .A3(new_n346), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n579), .A3(new_n622), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT95), .B1(new_n659), .B2(new_n576), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT41), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G113), .ZN(G15));
  NAND2_X1  g477(.A1(new_n655), .A2(new_n600), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  AND3_X1   g479(.A1(new_n622), .A2(new_n460), .A3(new_n614), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n620), .A2(new_n654), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT96), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G119), .ZN(G21));
  NOR2_X1   g484(.A1(new_n592), .A2(new_n654), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n565), .A3(new_n595), .A4(new_n586), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G122), .ZN(G24));
  AND2_X1   g487(.A1(new_n649), .A2(new_n615), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n667), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G125), .ZN(G27));
  NAND3_X1  g490(.A1(new_n290), .A2(new_n296), .A3(new_n187), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n290), .A2(new_n296), .A3(KEYINPUT97), .A4(new_n187), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n679), .A2(new_n465), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n560), .A3(new_n649), .ZN(new_n682));
  NOR2_X1   g496(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n683), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G131), .ZN(G33));
  AND2_X1   g502(.A1(new_n626), .A2(KEYINPUT99), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n626), .A2(KEYINPUT99), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n681), .B(new_n560), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G134), .ZN(G36));
  XNOR2_X1  g506(.A(new_n635), .B(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n575), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n565), .A2(new_n574), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n694), .B(KEYINPUT43), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n696), .B2(KEYINPUT101), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n697), .A2(new_n585), .A3(new_n614), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT44), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n679), .A2(new_n680), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n350), .A2(new_n351), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  OAI21_X1  g519(.A(G469), .B1(new_n705), .B2(G902), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n346), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n707), .A2(new_n711), .A3(new_n346), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(new_n300), .A3(new_n631), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n703), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G137), .ZN(G39));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n300), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT47), .ZN(new_n718));
  INV_X1    g532(.A(new_n702), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n559), .A3(new_n649), .ZN(new_n720));
  OR3_X1    g534(.A1(new_n718), .A2(new_n622), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G140), .ZN(G42));
  INV_X1    g536(.A(new_n431), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n697), .A2(new_n723), .A3(new_n699), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n697), .A2(KEYINPUT112), .A3(new_n723), .A4(new_n699), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n654), .B(new_n702), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n560), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT48), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n582), .B1(new_n726), .B2(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n667), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n643), .A2(new_n579), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n723), .A3(new_n658), .A4(new_n719), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n565), .A2(new_n575), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(G952), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(G953), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n730), .A2(new_n732), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n634), .A2(new_n188), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n731), .A2(new_n658), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n743));
  AOI211_X1 g557(.A(KEYINPUT114), .B(KEYINPUT50), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n742), .B2(KEYINPUT114), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n743), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n744), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n728), .A2(new_n615), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n735), .A2(new_n565), .A3(new_n575), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n653), .A2(new_n346), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n463), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n702), .B1(new_n718), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n753), .B1(new_n756), .B2(new_n731), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n749), .A2(new_n746), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n747), .A2(new_n748), .A3(new_n745), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n757), .A3(new_n752), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT51), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n740), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n621), .B(new_n623), .C1(new_n627), .C2(new_n649), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n675), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n642), .A2(new_n556), .A3(new_n613), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n583), .A2(new_n648), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n619), .A4(new_n636), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n675), .A3(new_n770), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n771), .A2(new_n773), .B1(KEYINPUT106), .B2(new_n772), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n772), .A2(KEYINPUT106), .A3(new_n767), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n389), .A2(new_n595), .A3(new_n648), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n594), .A2(new_n778), .A3(new_n598), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n681), .A2(new_n623), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT105), .B1(new_n681), .B2(new_n674), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n679), .A2(new_n465), .A3(new_n680), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n649), .A2(new_n615), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n691), .B(new_n780), .C1(new_n781), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n597), .A2(new_n563), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT104), .B1(new_n592), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n787), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT104), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n790), .A3(new_n297), .A4(new_n434), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n788), .A2(new_n584), .A3(new_n587), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n561), .A2(new_n616), .A3(new_n792), .A4(new_n588), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n687), .A2(new_n794), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n655), .A2(new_n600), .B1(new_n666), .B2(new_n667), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n656), .B1(new_n655), .B2(new_n577), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n659), .A2(KEYINPUT95), .A3(new_n576), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n796), .B(new_n672), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT103), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT103), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n661), .A2(new_n801), .A3(new_n672), .A4(new_n796), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n776), .A2(new_n777), .A3(new_n795), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n772), .B(new_n767), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n687), .A3(new_n805), .A4(new_n794), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n804), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT107), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n799), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n684), .B2(new_n686), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n777), .B1(new_n812), .B2(KEYINPUT109), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n687), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n776), .A2(new_n813), .A3(new_n794), .A4(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT108), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n806), .A2(new_n819), .A3(new_n777), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n806), .B2(new_n777), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n816), .B(new_n818), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n809), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n810), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n810), .A2(KEYINPUT111), .A3(new_n822), .A4(new_n823), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n763), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n763), .A2(KEYINPUT115), .A3(new_n826), .A4(new_n827), .ZN(new_n831));
  NOR2_X1   g645(.A1(G952), .A2(G953), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT116), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n694), .A2(new_n188), .A3(new_n463), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n754), .B(KEYINPUT49), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n734), .A3(new_n634), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n834), .A2(new_n837), .ZN(G75));
  OAI21_X1  g652(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n264), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n841), .A2(G210), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n293), .A2(new_n294), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n211), .ZN(new_n845));
  XOR2_X1   g659(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n846));
  XNOR2_X1  g660(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n843), .A2(new_n847), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n303), .A2(G952), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G51));
  AND3_X1   g665(.A1(new_n841), .A2(G469), .A3(new_n705), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n839), .A2(new_n817), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n822), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n347), .B(KEYINPUT57), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g672(.A(KEYINPUT118), .B(new_n856), .C1(new_n854), .C2(new_n822), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n337), .A2(new_n345), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n852), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT119), .B1(new_n863), .B2(new_n850), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n865));
  INV_X1    g679(.A(new_n850), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n852), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n864), .A2(new_n868), .ZN(G54));
  NAND3_X1  g683(.A1(new_n841), .A2(KEYINPUT58), .A3(G475), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(new_n451), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n451), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n871), .A2(KEYINPUT120), .A3(new_n866), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(G60));
  NOR2_X1   g691(.A1(new_n567), .A2(new_n569), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n571), .B(KEYINPUT59), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n855), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n826), .B2(new_n827), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n866), .B(new_n881), .C1(new_n882), .C2(new_n878), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(G63));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT60), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n840), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n612), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n549), .A2(new_n550), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n888), .B(new_n866), .C1(new_n889), .C2(new_n887), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g705(.A(new_n303), .B1(new_n432), .B2(G224), .ZN(new_n892));
  INV_X1    g706(.A(new_n803), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(new_n793), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n894), .B2(new_n303), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n844), .B1(G898), .B2(new_n303), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n895), .B(new_n896), .Z(G69));
  AND3_X1   g711(.A1(new_n721), .A2(new_n691), .A3(new_n766), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n560), .A2(new_n619), .A3(new_n636), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n714), .B1(new_n703), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n900), .A3(new_n687), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(G953), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n492), .A2(new_n493), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n445), .ZN(new_n904));
  NAND2_X1  g718(.A1(G900), .A2(G953), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n646), .A2(new_n766), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT62), .Z(new_n908));
  AOI211_X1 g722(.A(new_n559), .B(new_n526), .C1(new_n736), .C2(new_n787), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n465), .A3(new_n631), .A4(new_n719), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n715), .A2(KEYINPUT121), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT121), .B1(new_n715), .B2(new_n910), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n908), .B(new_n721), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n904), .B1(new_n913), .B2(new_n303), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n906), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n303), .B1(G227), .B2(G900), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n916), .B(new_n919), .ZN(G72));
  XNOR2_X1  g734(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n510), .A2(new_n264), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n494), .A2(new_n475), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n497), .B1(new_n926), .B2(new_n514), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n804), .A2(new_n807), .A3(new_n924), .A4(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT126), .Z(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n901), .B2(new_n894), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n505), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n866), .B(new_n929), .C1(new_n931), .C2(new_n925), .ZN(new_n932));
  OAI211_X1 g746(.A(KEYINPUT125), .B(new_n924), .C1(new_n913), .C2(new_n894), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(new_n925), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n924), .B1(new_n913), .B2(new_n894), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n505), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n934), .B2(new_n937), .ZN(G57));
endmodule


