//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  XNOR2_X1  g034(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n462), .B1(new_n479), .B2(new_n480), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n477), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT69), .A2(G114), .ZN(new_n489));
  OAI211_X1 g064(.A(G2104), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n463), .B2(new_n464), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n479), .A2(new_n480), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(new_n494), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n492), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT71), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n507), .B1(new_n504), .B2(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n501), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n506), .A2(new_n510), .A3(new_n514), .A4(new_n511), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(G88), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n506), .A2(new_n510), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(G50), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n518), .A2(new_n519), .B1(G651), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT73), .B1(new_n516), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n516), .A2(new_n526), .A3(KEYINPUT73), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n517), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n506), .A2(new_n510), .A3(KEYINPUT75), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n532), .A2(G51), .A3(G543), .A4(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n523), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n511), .A2(KEYINPUT74), .A3(G63), .A4(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n537), .A2(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n513), .A2(new_n515), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n534), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  AOI22_X1  g121(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n501), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT76), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT77), .B(G52), .Z(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n513), .A2(G90), .A3(new_n515), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND4_X1  g130(.A1(new_n532), .A2(G43), .A3(G543), .A4(new_n533), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n501), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n556), .B(new_n558), .C1(new_n543), .C2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND4_X1  g141(.A1(new_n532), .A2(G53), .A3(G543), .A4(new_n533), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n513), .A2(G91), .A3(new_n515), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n511), .A2(G65), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT78), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n568), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(new_n529), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n527), .ZN(G303));
  NAND3_X1  g152(.A1(new_n513), .A2(G87), .A3(new_n515), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n579));
  AND2_X1   g154(.A1(G49), .A2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n532), .A2(new_n533), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n513), .A2(G86), .A3(new_n515), .ZN(new_n583));
  AND2_X1   g158(.A1(G48), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n523), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n518), .A2(new_n584), .B1(new_n587), .B2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n550), .A2(G47), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n513), .A2(G85), .A3(new_n515), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n501), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n513), .A2(G92), .A3(new_n515), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n523), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n550), .A2(G54), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n497), .A2(new_n470), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT79), .B(G2100), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n483), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n462), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT80), .Z(new_n647));
  NOR2_X1   g222(.A1(G2072), .A2(G2078), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n444), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(KEYINPUT17), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n645), .B(new_n646), .C1(new_n444), .C2(new_n648), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n647), .A3(new_n645), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n665), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n666), .A2(KEYINPUT20), .A3(new_n665), .ZN(new_n671));
  OAI221_X1 g246(.A(new_n667), .B1(new_n665), .B2(new_n663), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NOR2_X1   g256(.A1(G166), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(G22), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(G1971), .ZN(new_n685));
  INV_X1    g260(.A(G305), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G16), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G6), .B2(G16), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT32), .B(G1981), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n684), .A2(G1971), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(G16), .A2(G23), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT84), .ZN(new_n694));
  NAND2_X1  g269(.A1(G288), .A2(KEYINPUT85), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n578), .A2(new_n581), .A3(new_n696), .A4(new_n579), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n694), .B1(new_n698), .B2(new_n681), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT33), .B(G1976), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n685), .A2(new_n692), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n481), .A2(G131), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n462), .A2(G107), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n483), .A2(KEYINPUT82), .A3(G119), .ZN(new_n709));
  AOI21_X1  g284(.A(KEYINPUT82), .B1(new_n483), .B2(G119), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n706), .B1(new_n707), .B2(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT83), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n705), .B1(new_n712), .B2(G29), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT35), .B(G1991), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n713), .B(new_n714), .Z(new_n715));
  MUX2_X1   g290(.A(G24), .B(G290), .S(G16), .Z(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G1986), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(G1986), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n685), .A2(new_n692), .A3(new_n720), .A4(new_n701), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n703), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n723), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n703), .A2(new_n719), .A3(new_n725), .A4(new_n721), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n724), .A2(new_n726), .B1(KEYINPUT86), .B2(KEYINPUT36), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT97), .ZN(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  NAND2_X1  g305(.A1(G162), .A2(G29), .ZN(new_n731));
  OR2_X1    g306(.A1(G29), .A2(G35), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n731), .A2(new_n730), .A3(new_n732), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n481), .A2(G140), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n483), .A2(G128), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n462), .A2(G116), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n704), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n704), .A2(G32), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT26), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G129), .B2(new_n483), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n754), .A2(new_n755), .B1(new_n481), .B2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n749), .B1(new_n757), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT24), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G34), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G160), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n737), .A2(new_n748), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n758), .A2(new_n759), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT91), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n704), .A2(G27), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G164), .B2(new_n704), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(new_n443), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n704), .B1(new_n778), .B2(G28), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(KEYINPUT93), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(G28), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n779), .B2(KEYINPUT93), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n777), .B1(new_n780), .B2(new_n782), .C1(new_n627), .C2(new_n704), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n768), .B2(new_n767), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n773), .A2(new_n776), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n735), .B1(new_n734), .B2(new_n736), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n771), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n681), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n604), .B2(new_n681), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n497), .A2(G127), .ZN(new_n792));
  INV_X1    g367(.A(G115), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n469), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(G2105), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT25), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n481), .A2(G139), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n795), .A2(KEYINPUT88), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT88), .B1(new_n795), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT89), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(KEYINPUT89), .B1(new_n800), .B2(new_n801), .ZN(new_n805));
  OR3_X1    g380(.A1(new_n804), .A2(new_n704), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G33), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n442), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n804), .A2(new_n805), .A3(new_n704), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n810), .A2(G2072), .A3(new_n807), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n787), .B(new_n791), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n681), .A2(G20), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT96), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT23), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G299), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1956), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n561), .A2(G16), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G16), .B2(G19), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT87), .B(G1341), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n681), .A2(G5), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G171), .B2(new_n681), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(G1961), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n819), .A2(new_n821), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n817), .A2(new_n822), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n812), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(G16), .A2(G21), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G286), .B2(new_n681), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G1966), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(G1966), .A3(new_n832), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n824), .A2(KEYINPUT94), .A3(G1961), .ZN(new_n837));
  AOI21_X1  g412(.A(KEYINPUT94), .B1(new_n824), .B2(G1961), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n729), .B1(new_n828), .B2(new_n840), .ZN(new_n841));
  NOR4_X1   g416(.A1(new_n812), .A2(new_n827), .A3(KEYINPUT97), .A4(new_n839), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n728), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n842), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n845), .A2(new_n727), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(G311));
  NAND2_X1  g423(.A1(new_n728), .A2(new_n843), .ZN(G150));
  NAND2_X1  g424(.A1(new_n604), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n513), .A2(G93), .A3(new_n515), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n532), .A2(G55), .A3(G543), .A4(new_n533), .ZN(new_n853));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n523), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(KEYINPUT99), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(KEYINPUT99), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G651), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n852), .B(new_n853), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(new_n560), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n560), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n851), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n860), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT100), .Z(G145));
  XOR2_X1   g446(.A(new_n742), .B(KEYINPUT101), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n496), .A2(new_n499), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT69), .ZN(new_n874));
  INV_X1    g449(.A(G114), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(KEYINPUT69), .A2(G114), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(G2105), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(G126), .A2(new_n483), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n872), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n757), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n872), .B(G164), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n757), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n802), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n483), .A2(G130), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n462), .A2(G118), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(G142), .B2(new_n481), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n618), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n712), .B(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n885), .B(new_n887), .C1(new_n804), .C2(new_n805), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n890), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n890), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n627), .B(G160), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G162), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g482(.A(G868), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n698), .A2(G303), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  NAND2_X1  g485(.A1(G290), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n590), .A2(KEYINPUT102), .A3(new_n591), .A4(new_n593), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n686), .ZN(new_n914));
  NAND3_X1  g489(.A1(G166), .A2(new_n695), .A3(new_n697), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(G305), .A3(new_n912), .ZN(new_n916));
  AND4_X1   g491(.A1(new_n909), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n914), .A2(new_n916), .B1(new_n915), .B2(new_n909), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n917), .A2(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n613), .B(new_n863), .Z(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n603), .A2(G299), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n603), .A2(G299), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n929), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n927), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n925), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n613), .B(new_n863), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n928), .B2(new_n929), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n924), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n937), .B(new_n935), .C1(new_n920), .C2(new_n923), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n908), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n860), .A2(new_n908), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OR3_X1    g518(.A1(new_n941), .A2(KEYINPUT103), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT103), .B1(new_n941), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(G295));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n940), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(G868), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n949), .B2(new_n942), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n941), .A2(KEYINPUT104), .A3(new_n943), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(G331));
  NOR2_X1   g527(.A1(new_n928), .A2(new_n929), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n861), .A2(G286), .A3(new_n862), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G286), .B1(new_n861), .B2(new_n862), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n955), .A2(G301), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n863), .A2(G168), .ZN(new_n958));
  AOI21_X1  g533(.A(G171), .B1(new_n958), .B2(new_n954), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n953), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(G301), .B1(new_n955), .B2(new_n956), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(G171), .A3(new_n954), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n933), .A3(new_n930), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n919), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  INV_X1    g541(.A(G37), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n921), .A2(new_n960), .A3(new_n963), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT105), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n964), .B2(new_n919), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n966), .A4(new_n968), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(KEYINPUT44), .A3(new_n969), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(G397));
  INV_X1    g555(.A(KEYINPUT125), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n528), .A2(G8), .A3(new_n529), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n468), .A2(new_n471), .ZN(new_n987));
  INV_X1    g562(.A(G125), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n479), .B2(new_n480), .ZN(new_n989));
  INV_X1    g564(.A(new_n466), .ZN(new_n990));
  OAI21_X1  g565(.A(G2105), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n991), .A3(G40), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(G160), .A2(KEYINPUT106), .A3(G40), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G164), .B2(G1384), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n873), .B2(new_n881), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT45), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n996), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G164), .B2(G1384), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n882), .A2(KEYINPUT112), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n996), .ZN(new_n1011));
  INV_X1    g586(.A(new_n999), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1004), .A2(G1971), .B1(new_n1014), .B2(G2090), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n986), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1007), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n882), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(new_n994), .A3(new_n995), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1018), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT112), .B1(new_n882), .B2(new_n1008), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1005), .B(G1384), .C1(new_n873), .C2(new_n881), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT50), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1020), .A2(new_n994), .A3(new_n995), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(KEYINPUT115), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1027), .A3(new_n730), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1001), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1029));
  NOR3_X1   g604(.A1(G164), .A2(new_n997), .A3(G1384), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1003), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1011), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1971), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1017), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1016), .B1(new_n1036), .B2(new_n986), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n695), .A2(G1976), .A3(new_n697), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1006), .A2(new_n994), .A3(new_n1009), .A4(new_n995), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1038), .A2(G8), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n583), .A2(new_n588), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n583), .B2(new_n588), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n583), .A2(new_n588), .A3(new_n1044), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1047), .A2(new_n1050), .A3(G8), .A4(new_n1039), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1042), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1017), .B1(new_n1053), .B2(new_n1011), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1038), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT113), .B1(new_n1055), .B2(KEYINPUT52), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1057), .B(new_n1058), .C1(new_n1054), .C2(new_n1038), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1052), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1037), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n996), .B1(KEYINPUT50), .B2(new_n1012), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1961), .B1(new_n1063), .B2(new_n1010), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1004), .A2(new_n443), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n996), .A2(new_n1030), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n997), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n443), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT123), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1068), .A2(new_n1069), .A3(new_n1072), .A4(new_n443), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G301), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1066), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1004), .B2(new_n443), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n992), .B(new_n1078), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1079));
  NOR4_X1   g654(.A1(new_n1077), .A2(new_n1079), .A3(new_n1064), .A4(G171), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1062), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n1083));
  AND3_X1   g658(.A1(G286), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(G286), .B2(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1086), .B2(KEYINPUT121), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT45), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1000), .A2(new_n994), .A3(new_n995), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n834), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1010), .A2(new_n1011), .A3(new_n768), .A4(new_n1013), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1085), .ZN(new_n1093));
  NAND3_X1  g668(.A1(G286), .A2(new_n1083), .A3(G8), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1017), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1087), .B(new_n1096), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1092), .A2(G8), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n1086), .C1(KEYINPUT121), .C2(new_n1082), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1067), .A2(new_n1074), .A3(G301), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1077), .A2(new_n1064), .A3(new_n1079), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1102), .B(KEYINPUT54), .C1(G301), .C2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1061), .A2(new_n1081), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1004), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n568), .A2(new_n1109), .A3(new_n574), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1108), .A2(new_n1113), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT61), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1108), .A2(new_n1113), .A3(new_n1106), .A4(new_n1110), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1053), .A2(new_n1011), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1039), .A2(KEYINPUT117), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(G1341), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1996), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1004), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n561), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1134), .A3(new_n561), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1116), .A2(new_n1122), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(G2067), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1348), .B1(new_n1063), .B2(new_n1010), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n604), .B1(new_n1140), .B2(KEYINPUT119), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n747), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1139), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(KEYINPUT60), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(new_n603), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1141), .A2(new_n1147), .B1(KEYINPUT119), .B2(new_n1140), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1136), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n603), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1121), .B1(new_n1152), .B2(new_n1115), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1105), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G288), .A2(G1976), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1051), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1054), .B1(new_n1156), .B2(new_n1045), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1060), .B2(new_n1016), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT114), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT114), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1157), .B(new_n1160), .C1(new_n1060), .C2(new_n1016), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n986), .B1(G8), .B2(new_n1015), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT116), .B1(new_n1060), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1057), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1055), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1015), .A2(G8), .ZN(new_n1169));
  INV_X1    g744(.A(new_n986), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT116), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .A4(new_n1052), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1099), .A2(G286), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1174), .A2(KEYINPUT63), .A3(new_n1016), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1164), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n1061), .B2(new_n1174), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1162), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n981), .B1(new_n1154), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1042), .A2(new_n1051), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1181));
  AOI21_X1  g756(.A(G2090), .B1(new_n1111), .B2(new_n1018), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1182), .A2(new_n1027), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1170), .B1(new_n1183), .B2(new_n1017), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1181), .A2(new_n1184), .A3(new_n1016), .A4(new_n1174), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1164), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1187), .A2(new_n1188), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1153), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1140), .A2(KEYINPUT119), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1140), .A2(KEYINPUT119), .A3(new_n604), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n603), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1150), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1190), .B1(new_n1196), .B2(new_n1136), .ZN(new_n1197));
  OAI211_X1 g772(.A(KEYINPUT125), .B(new_n1189), .C1(new_n1197), .C2(new_n1105), .ZN(new_n1198));
  OR2_X1    g773(.A1(new_n1101), .A2(KEYINPUT62), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1101), .A2(KEYINPUT62), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1199), .A2(new_n1061), .A3(new_n1075), .A4(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1179), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n996), .A2(new_n998), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1203), .A2(G1996), .A3(new_n757), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT109), .Z(new_n1205));
  XNOR2_X1  g780(.A(new_n742), .B(new_n747), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1206), .B1(G1996), .B2(new_n757), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1203), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT110), .Z(new_n1210));
  AND2_X1   g785(.A1(new_n712), .A2(new_n714), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n712), .A2(new_n714), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1203), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(G290), .A2(G1986), .ZN(new_n1215));
  XOR2_X1   g790(.A(new_n1215), .B(KEYINPUT107), .Z(new_n1216));
  NAND2_X1  g791(.A1(G290), .A2(G1986), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT108), .ZN(new_n1218));
  OR2_X1    g793(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1214), .B1(new_n1203), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1202), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1203), .ZN(new_n1222));
  OR3_X1    g797(.A1(new_n1222), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1223));
  OAI21_X1  g798(.A(KEYINPUT46), .B1(new_n1222), .B2(G1996), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1206), .A2(new_n884), .ZN(new_n1225));
  AOI22_X1  g800(.A1(new_n1223), .A2(new_n1224), .B1(new_n1203), .B2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(KEYINPUT47), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1228));
  OR2_X1    g803(.A1(new_n742), .A2(G2067), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1216), .A2(new_n1203), .ZN(new_n1231));
  XOR2_X1   g806(.A(new_n1231), .B(KEYINPUT126), .Z(new_n1232));
  NAND2_X1  g807(.A1(new_n1232), .A2(KEYINPUT48), .ZN(new_n1233));
  NOR2_X1   g808(.A1(new_n1232), .A2(KEYINPUT48), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1234), .A2(new_n1214), .ZN(new_n1235));
  AOI211_X1 g810(.A(new_n1227), .B(new_n1230), .C1(new_n1233), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1221), .A2(new_n1236), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g812(.A(G319), .ZN(new_n1239));
  NOR3_X1   g813(.A1(G401), .A2(new_n1239), .A3(G227), .ZN(new_n1240));
  OAI21_X1  g814(.A(new_n1240), .B1(new_n678), .B2(new_n679), .ZN(new_n1241));
  AOI21_X1  g815(.A(new_n1241), .B1(new_n904), .B2(new_n905), .ZN(new_n1242));
  AND3_X1   g816(.A1(new_n976), .A2(KEYINPUT127), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g817(.A(KEYINPUT127), .B1(new_n976), .B2(new_n1242), .ZN(new_n1244));
  NOR2_X1   g818(.A1(new_n1243), .A2(new_n1244), .ZN(G308));
  NAND2_X1  g819(.A1(new_n976), .A2(new_n1242), .ZN(G225));
endmodule


