//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G107), .C2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G77), .B2(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n209), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n229), .A2(new_n232), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT65), .B(G250), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G257), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n222), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  XOR2_X1   g0049(.A(G97), .B(G107), .Z(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G274), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT66), .B(G45), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n235), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n257), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n261), .A2(new_n215), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n226), .B2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n223), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n265), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n259), .B1(new_n211), .B2(new_n264), .C1(new_n272), .C2(new_n262), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT13), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT14), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(G179), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(new_n279), .A3(G169), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n235), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT67), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(KEYINPUT67), .A3(new_n235), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n210), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n234), .A2(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n202), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT11), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n295), .A2(new_n210), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n254), .A2(G20), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n285), .A2(new_n299), .A3(new_n286), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n293), .B(new_n298), .C1(new_n210), .C2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n296), .B1(new_n295), .B2(new_n210), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n281), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n275), .B2(G190), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n275), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT74), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n234), .B1(new_n201), .B2(new_n203), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(G150), .B2(new_n288), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n225), .A2(KEYINPUT8), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT8), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G58), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT68), .B1(new_n225), .B2(KEYINPUT8), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT69), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n317), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT69), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n319), .B(new_n320), .C1(new_n321), .C2(new_n312), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n311), .B1(new_n323), .B2(new_n290), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n287), .B1(new_n222), .B2(new_n295), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n222), .B2(new_n300), .ZN(new_n326));
  XOR2_X1   g0126(.A(new_n326), .B(KEYINPUT9), .Z(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n261), .ZN(new_n329));
  NAND2_X1  g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n270), .A2(G222), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G223), .A2(G1698), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n335), .C1(G77), .C2(new_n331), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(new_n259), .C1(new_n223), .C2(new_n264), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT71), .B(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n344));
  OR2_X1    g0144(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n340), .A2(KEYINPUT72), .A3(KEYINPUT10), .A4(new_n342), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n337), .A2(new_n276), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n326), .B(new_n348), .C1(G179), .C2(new_n337), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n300), .A2(new_n202), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n290), .ZN(new_n353));
  XOR2_X1   g0153(.A(new_n353), .B(KEYINPUT70), .Z(new_n354));
  INV_X1    g0154(.A(new_n288), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n354), .B1(new_n234), .B2(new_n202), .C1(new_n355), .C2(new_n321), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n351), .B1(new_n356), .B2(new_n287), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n295), .A2(new_n202), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G238), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n331), .B(new_n359), .C1(new_n226), .C2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n335), .C1(G107), .C2(new_n331), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n262), .A2(G244), .A3(new_n263), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n259), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n341), .ZN(new_n364));
  INV_X1    g0164(.A(new_n363), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G190), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n357), .A2(new_n358), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n350), .A2(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n318), .A2(new_n300), .A3(new_n322), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n295), .B1(new_n318), .B2(new_n322), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT76), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n314), .A2(G58), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n225), .A2(KEYINPUT8), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT68), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n320), .B1(new_n375), .B2(new_n319), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n316), .A2(KEYINPUT69), .A3(new_n317), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n294), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT76), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n318), .A2(new_n300), .A3(new_n322), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT75), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n268), .B2(new_n234), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n234), .A4(new_n330), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n225), .A2(new_n210), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n203), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n288), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n383), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n329), .A2(new_n234), .A3(new_n330), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n210), .B1(new_n398), .B2(new_n385), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n383), .B(new_n394), .C1(new_n399), .C2(new_n391), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n287), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n399), .A2(new_n391), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n382), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n223), .A2(G1698), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n407), .B1(G223), .B2(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n262), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n262), .A2(G232), .A3(new_n263), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n410), .A2(new_n411), .A3(new_n258), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n412), .A2(new_n306), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(G190), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n406), .A2(KEYINPUT17), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n372), .A2(new_n381), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n394), .B1(new_n399), .B2(new_n391), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT75), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n405), .A2(new_n418), .A3(new_n400), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n416), .A2(new_n419), .A3(new_n413), .A4(new_n414), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n412), .A2(new_n276), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n412), .A2(G179), .ZN(new_n425));
  AOI221_X4 g0225(.A(new_n423), .B1(new_n424), .B2(new_n425), .C1(new_n416), .C2(new_n419), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n416), .A2(new_n419), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n425), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT18), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n415), .B(new_n422), .C1(new_n426), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n357), .A2(new_n358), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n363), .A2(new_n276), .ZN(new_n432));
  INV_X1    g0232(.A(G179), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n365), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n309), .A2(new_n369), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(G238), .B(new_n270), .C1(new_n266), .C2(new_n267), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT81), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n331), .A2(new_n442), .A3(G238), .A4(new_n270), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G116), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT82), .ZN(new_n446));
  OAI21_X1  g0246(.A(G244), .B1(new_n266), .B2(new_n267), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(new_n270), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n331), .A2(KEYINPUT82), .A3(G244), .A4(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n335), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n214), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n255), .A2(new_n452), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n262), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n433), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT19), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n290), .B2(new_n215), .ZN(new_n459));
  AOI21_X1  g0259(.A(G20), .B1(new_n329), .B2(new_n330), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G68), .ZN(new_n461));
  XOR2_X1   g0261(.A(KEYINPUT83), .B(G87), .Z(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n207), .ZN(new_n463));
  AOI21_X1  g0263(.A(G20), .B1(new_n265), .B2(KEYINPUT19), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n459), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n287), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n352), .A2(new_n295), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n352), .B(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n254), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n285), .A2(new_n294), .A3(new_n469), .A4(new_n286), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n451), .A2(new_n456), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n457), .B(new_n471), .C1(new_n472), .C2(G169), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n214), .B1(new_n329), .B2(new_n330), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT4), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(KEYINPUT78), .ZN(new_n476));
  OAI21_X1  g0276(.A(G1698), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G283), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n261), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n447), .B2(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n331), .A2(G244), .A3(new_n270), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n475), .B1(new_n482), .B2(KEYINPUT78), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n335), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT79), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT5), .B(G41), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n453), .ZN(new_n487));
  INV_X1    g0287(.A(G274), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(KEYINPUT79), .A3(G274), .A4(new_n453), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(G257), .A3(new_n262), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT80), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n335), .B1(new_n453), .B2(new_n486), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(KEYINPUT80), .A3(G257), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n484), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n276), .ZN(new_n499));
  OAI21_X1  g0299(.A(G107), .B1(new_n384), .B2(new_n386), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n215), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n503), .B2(new_n206), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(KEYINPUT6), .A3(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n288), .A2(G77), .ZN(new_n508));
  XOR2_X1   g0308(.A(new_n508), .B(KEYINPUT77), .Z(new_n509));
  NAND3_X1  g0309(.A1(new_n500), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n287), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n294), .A2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n470), .A2(new_n215), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n484), .A2(new_n433), .A3(new_n497), .A4(new_n491), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n499), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n498), .A2(G200), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n512), .B(new_n514), .C1(new_n510), .C2(new_n287), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n484), .A2(G190), .A3(new_n497), .A4(new_n491), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n451), .A2(new_n456), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n341), .ZN(new_n524));
  INV_X1    g0324(.A(new_n470), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G87), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n466), .A2(new_n467), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n451), .A2(G190), .A3(new_n456), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n473), .A2(new_n518), .A3(new_n522), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n295), .A2(new_n502), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT25), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n470), .A2(new_n502), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n216), .A2(G1698), .ZN(new_n535));
  OAI221_X1 g0335(.A(new_n535), .B1(G250), .B2(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n536));
  INV_X1    g0336(.A(G294), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n261), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n335), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n487), .A2(G264), .A3(new_n262), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT90), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n495), .A2(KEYINPUT90), .A3(G264), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n539), .A2(new_n491), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n306), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n539), .A2(new_n491), .A3(new_n338), .A4(new_n540), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n234), .A2(G33), .A3(G116), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n502), .A2(KEYINPUT23), .A3(G20), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT23), .B1(new_n502), .B2(G20), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n213), .A2(KEYINPUT87), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n234), .C1(new_n267), .C2(new_n266), .ZN(new_n554));
  XNOR2_X1  g0354(.A(KEYINPUT88), .B(KEYINPUT22), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n460), .B2(new_n553), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT24), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n554), .A2(new_n556), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n331), .A2(new_n555), .A3(new_n234), .A4(new_n553), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n552), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT89), .B1(new_n566), .B2(new_n287), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n563), .B2(new_n552), .ZN(new_n568));
  AOI211_X1 g0368(.A(KEYINPUT24), .B(new_n551), .C1(new_n561), .C2(new_n562), .ZN(new_n569));
  OAI211_X1 g0369(.A(KEYINPUT89), .B(new_n287), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n534), .B(new_n547), .C1(new_n567), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT91), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n534), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n287), .B1(new_n568), .B2(new_n569), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT89), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n575), .B1(new_n578), .B2(new_n570), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(KEYINPUT91), .A3(new_n547), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n534), .B1(new_n567), .B2(new_n571), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n539), .A2(new_n491), .A3(new_n540), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G169), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n433), .B2(new_n544), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G116), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n295), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n525), .A2(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(G20), .ZN(new_n590));
  AOI21_X1  g0390(.A(G20), .B1(G33), .B2(G283), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n261), .A2(G97), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n591), .B2(new_n592), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n283), .B(new_n590), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n588), .B(new_n589), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G264), .A2(G1698), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n331), .B(new_n601), .C1(new_n216), .C2(G1698), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(new_n335), .C1(G303), .C2(new_n331), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n495), .A2(G270), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n491), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n600), .A2(G169), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n605), .A2(new_n433), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n600), .ZN(new_n611));
  INV_X1    g0411(.A(new_n608), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n600), .A2(G169), .A3(new_n605), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n605), .A2(new_n338), .ZN(new_n615));
  AOI211_X1 g0415(.A(new_n600), .B(new_n615), .C1(G200), .C2(new_n605), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n530), .A2(new_n581), .A3(new_n586), .A4(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n439), .A2(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n304), .A2(new_n435), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n420), .B(KEYINPUT17), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n307), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n427), .A2(new_n428), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n423), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n428), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n346), .A3(new_n347), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n349), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n473), .A2(new_n529), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(new_n518), .ZN(new_n632));
  XOR2_X1   g0432(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n634), .B(KEYINPUT94), .C1(KEYINPUT26), .C2(new_n632), .ZN(new_n635));
  INV_X1    g0435(.A(new_n473), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT94), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n518), .A2(new_n522), .A3(new_n473), .A4(new_n529), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n574), .B2(new_n580), .ZN(new_n641));
  INV_X1    g0441(.A(new_n614), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n586), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n641), .A2(KEYINPUT92), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT92), .B1(new_n641), .B2(new_n643), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n635), .B(new_n639), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n630), .B1(new_n438), .B2(new_n647), .ZN(G369));
  XOR2_X1   g0448(.A(new_n617), .B(KEYINPUT96), .Z(new_n649));
  INV_X1    g0449(.A(G13), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G20), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n235), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT95), .ZN(new_n654));
  INV_X1    g0454(.A(G213), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n652), .B2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(KEYINPUT95), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n600), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n649), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n614), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n660), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n586), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT97), .ZN(new_n669));
  INV_X1    g0469(.A(new_n585), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n579), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n574), .B2(new_n580), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n579), .B2(new_n667), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n614), .A2(new_n667), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n674), .A2(new_n677), .B1(new_n586), .B2(new_n660), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(G399));
  NAND2_X1  g0480(.A1(new_n463), .A2(new_n587), .ZN(new_n681));
  INV_X1    g0481(.A(new_n230), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(new_n254), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT98), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  INV_X1    g0487(.A(new_n683), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n686), .B(new_n687), .C1(new_n233), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n484), .A2(new_n491), .A3(new_n497), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n472), .A3(new_n610), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT30), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n523), .A2(new_n605), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n433), .A3(new_n498), .A4(new_n544), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n660), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT100), .ZN(new_n699));
  XNOR2_X1  g0499(.A(KEYINPUT99), .B(KEYINPUT31), .ZN(new_n700));
  OR3_X1    g0500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT31), .B1(new_n697), .B2(new_n660), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n702), .A2(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n672), .A2(new_n530), .A3(new_n617), .A4(new_n667), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT101), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n701), .B(new_n703), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n646), .A2(new_n710), .A3(new_n667), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n641), .A2(new_n643), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n631), .A2(new_n518), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT26), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n633), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n712), .A2(new_n714), .A3(new_n473), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n667), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n709), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n690), .B1(new_n720), .B2(G1), .ZN(G364));
  AOI21_X1  g0521(.A(KEYINPUT102), .B1(new_n665), .B2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n664), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n254), .B1(new_n651), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n683), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n665), .A2(KEYINPUT102), .A3(G330), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n724), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n433), .A2(new_n306), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n234), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(KEYINPUT33), .A2(G317), .ZN(new_n733));
  NAND2_X1  g0533(.A1(KEYINPUT33), .A2(G317), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n331), .B1(new_n738), .B2(G329), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n234), .B1(new_n736), .B2(G190), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n537), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n234), .A2(new_n338), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n433), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n735), .B(new_n741), .C1(G322), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n730), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT105), .B(G326), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n731), .A2(new_n743), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(new_n749), .B1(new_n751), .B2(G311), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n341), .A2(new_n433), .A3(new_n731), .ZN(new_n754));
  INV_X1    g0554(.A(G303), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n341), .A2(new_n433), .A3(new_n742), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT104), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n753), .B1(new_n478), .B2(new_n754), .C1(new_n755), .C2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n331), .B1(new_n747), .B2(new_n222), .ZN(new_n762));
  INV_X1    g0562(.A(new_n754), .ZN(new_n763));
  INV_X1    g0563(.A(new_n732), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n763), .A2(G107), .B1(G68), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n202), .B2(new_n750), .ZN(new_n766));
  INV_X1    g0566(.A(new_n740), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n762), .B(new_n766), .C1(G97), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n760), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n462), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n738), .A2(G159), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT32), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n771), .A2(KEYINPUT32), .B1(G58), .B2(new_n745), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n768), .A2(new_n770), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n761), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT106), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n235), .B1(G20), .B2(new_n276), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n682), .A2(new_n331), .ZN(new_n779));
  INV_X1    g0579(.A(new_n256), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n779), .B1(new_n233), .B2(new_n780), .C1(new_n249), .C2(new_n452), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n331), .A2(new_n230), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(G116), .B2(new_n230), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n650), .A2(new_n261), .A3(KEYINPUT103), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT103), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G13), .B2(G33), .ZN(new_n787));
  AOI21_X1  g0587(.A(G20), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n777), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n778), .A2(new_n727), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n664), .B2(new_n788), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n729), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  OAI21_X1  g0594(.A(new_n473), .B1(new_n634), .B2(KEYINPUT94), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT92), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n578), .A2(new_n570), .ZN(new_n797));
  AND4_X1   g0597(.A1(KEYINPUT91), .A2(new_n797), .A3(new_n534), .A4(new_n547), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT91), .B1(new_n579), .B2(new_n547), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n530), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n671), .A2(new_n614), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n641), .A2(KEYINPUT92), .A3(new_n643), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n795), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n660), .B1(new_n804), .B2(new_n635), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n436), .A2(new_n667), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n431), .A2(new_n660), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n367), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n435), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n805), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n709), .ZN(new_n815));
  INV_X1    g0615(.A(new_n727), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT109), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n709), .B2(new_n814), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n785), .A2(new_n787), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n777), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n202), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n769), .A2(G50), .B1(G58), .B2(new_n767), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n268), .B1(new_n738), .B2(G132), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(new_n210), .C2(new_n754), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT108), .B(G143), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n745), .A2(new_n828), .B1(new_n751), .B2(G159), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n748), .A2(G137), .ZN(new_n830));
  INV_X1    g0630(.A(G150), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n732), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  NOR2_X1   g0633(.A1(new_n744), .A2(new_n537), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n769), .A2(G107), .ZN(new_n835));
  XOR2_X1   g0635(.A(KEYINPUT107), .B(G283), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n764), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n763), .A2(G87), .B1(G97), .B2(new_n767), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n747), .A2(new_n755), .B1(new_n737), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n331), .B(new_n840), .C1(G116), .C2(new_n751), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n835), .A2(new_n837), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n827), .A2(new_n833), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n777), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n822), .A2(new_n727), .A3(new_n824), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n820), .A2(new_n845), .ZN(G384));
  AND3_X1   g0646(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n618), .A2(KEYINPUT101), .A3(new_n667), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n704), .A2(new_n705), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n698), .A2(new_n700), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n303), .A2(new_n660), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n304), .A2(new_n307), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n304), .A2(new_n667), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(KEYINPUT113), .A2(KEYINPUT40), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n852), .A2(new_n812), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n658), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n405), .A2(new_n417), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n370), .B2(new_n371), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n430), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n427), .B1(new_n428), .B2(new_n859), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n420), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n428), .B2(new_n859), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n866), .A2(new_n420), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n867), .B2(new_n864), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n812), .B1(new_n854), .B2(new_n855), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n850), .B2(new_n851), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n858), .B(new_n873), .C1(KEYINPUT113), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n427), .A2(new_n859), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n621), .B2(new_n626), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n863), .A2(new_n864), .A3(new_n420), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n864), .B1(new_n863), .B2(new_n420), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n870), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n872), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT40), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n886), .A2(new_n852), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(G330), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n723), .B1(new_n850), .B2(new_n851), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n439), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n887), .A2(new_n439), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n719), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n438), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n629), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n871), .B2(new_n872), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n882), .A2(new_n872), .A3(new_n895), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT112), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n281), .A2(new_n303), .A3(new_n667), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n862), .B2(new_n868), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT39), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT112), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n882), .A2(new_n872), .A3(new_n895), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n900), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n626), .A2(new_n859), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n646), .A2(new_n667), .A3(new_n812), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n806), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n856), .A3(new_n873), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n894), .B(new_n913), .Z(new_n914));
  XNOR2_X1  g0714(.A(new_n891), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n254), .B2(new_n651), .ZN(new_n916));
  OR3_X1    g0716(.A1(new_n388), .A2(new_n233), .A3(new_n202), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n201), .A2(G68), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n254), .B(G13), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT111), .ZN(new_n920));
  OAI211_X1 g0720(.A(G20), .B(new_n260), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n587), .B(new_n921), .C1(KEYINPUT35), .C2(new_n506), .ZN(new_n922));
  XNOR2_X1  g0722(.A(KEYINPUT110), .B(KEYINPUT36), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n916), .A2(new_n920), .A3(new_n924), .ZN(G367));
  INV_X1    g0725(.A(KEYINPUT114), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT42), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n674), .A2(new_n677), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n518), .A2(new_n667), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n518), .B(new_n522), .C1(new_n520), .C2(new_n667), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n927), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n930), .A2(new_n586), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n660), .B1(new_n933), .B2(new_n518), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n926), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n932), .A2(new_n926), .A3(new_n934), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT43), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n667), .A2(new_n527), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n631), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n636), .A2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n928), .A2(new_n927), .A3(new_n931), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n938), .A2(new_n939), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n937), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n945), .A3(new_n935), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n939), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n931), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n676), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n946), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n946), .B2(new_n951), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n683), .B(KEYINPUT41), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT115), .B1(new_n678), .B2(new_n952), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n678), .A2(KEYINPUT115), .A3(new_n952), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n678), .A2(new_n952), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT44), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n963), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n675), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n963), .A2(new_n965), .A3(new_n968), .A4(new_n676), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n674), .B(new_n677), .Z(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n666), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n970), .A2(new_n720), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n958), .B1(new_n974), .B2(new_n720), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n956), .B1(new_n975), .B2(new_n726), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n740), .A2(new_n210), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n769), .B2(G58), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n763), .A2(G77), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G159), .A2(new_n764), .B1(new_n738), .B2(G137), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n748), .A2(new_n828), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n745), .A2(G150), .ZN(new_n983));
  INV_X1    g0783(.A(new_n201), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n268), .B1(new_n751), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n760), .A2(new_n587), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n987), .A2(KEYINPUT46), .B1(new_n537), .B2(new_n732), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n987), .A2(KEYINPUT46), .ZN(new_n989));
  INV_X1    g0789(.A(new_n836), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n750), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n748), .A2(G311), .B1(new_n767), .B2(G107), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n755), .B2(new_n744), .ZN(new_n993));
  NOR4_X1   g0793(.A1(new_n988), .A2(new_n989), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n994), .B1(new_n215), .B2(new_n754), .C1(new_n995), .C2(new_n737), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n986), .B1(new_n996), .B2(new_n331), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n777), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n944), .A2(new_n788), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n779), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n789), .B1(new_n230), .B2(new_n352), .C1(new_n245), .C2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n999), .A2(new_n727), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n976), .A2(new_n1003), .ZN(G387));
  OR2_X1    g0804(.A1(new_n973), .A2(new_n720), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n973), .A2(new_n720), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n683), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n674), .A2(new_n788), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n779), .B1(new_n241), .B2(new_n256), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n681), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n783), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n210), .A2(new_n202), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n321), .A2(G50), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT116), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n681), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n452), .C1(KEYINPUT50), .C2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1011), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n682), .A2(new_n502), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n788), .B(new_n777), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G322), .A2(new_n748), .B1(new_n764), .B2(G311), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n755), .B2(new_n750), .C1(new_n995), .C2(new_n744), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT48), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n537), .B2(new_n760), .C1(new_n740), .C2(new_n990), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n738), .A2(new_n749), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n331), .B1(new_n763), .B2(G116), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n744), .A2(new_n222), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n468), .A2(new_n740), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n760), .A2(new_n202), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G150), .C2(new_n738), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n318), .A2(new_n322), .A3(new_n764), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n754), .A2(new_n215), .B1(new_n210), .B2(new_n750), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n268), .B(new_n1033), .C1(G159), .C2(new_n748), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1027), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n816), .B(new_n1019), .C1(new_n1036), .C2(new_n777), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n973), .A2(new_n726), .B1(new_n1008), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1007), .A2(new_n1038), .ZN(G393));
  AOI22_X1  g0839(.A1(new_n769), .A2(G68), .B1(new_n738), .B2(new_n828), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT117), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n763), .A2(G87), .B1(G77), .B2(new_n767), .ZN(new_n1042));
  INV_X1    g0842(.A(G159), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n747), .A2(new_n831), .B1(new_n744), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT51), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1044), .A2(new_n1045), .B1(new_n984), .B2(new_n764), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1041), .A2(new_n331), .A3(new_n1042), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n750), .A2(new_n321), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n747), .A2(new_n995), .B1(new_n744), .B2(new_n839), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT52), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n331), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .C1(new_n502), .C2(new_n754), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G322), .A2(new_n738), .B1(new_n767), .B2(G116), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n760), .B2(new_n990), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n732), .A2(new_n755), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n750), .A2(new_n537), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n777), .B1(new_n1050), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n952), .A2(new_n788), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n789), .B1(new_n215), .B2(new_n230), .C1(new_n252), .C2(new_n1001), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1060), .A2(new_n727), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n970), .A2(new_n971), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n725), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n688), .B1(new_n1064), .B2(new_n1006), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n974), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(G390));
  AND3_X1   g0868(.A1(new_n708), .A2(G330), .A3(new_n812), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n856), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n883), .A2(new_n899), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n806), .B1(new_n717), .B2(new_n811), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n856), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n900), .B1(new_n911), .B2(new_n856), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1070), .B(new_n1074), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n807), .B1(new_n805), .B2(new_n812), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n856), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n899), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n898), .A2(new_n906), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1073), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n852), .A2(G330), .A3(new_n812), .A4(new_n856), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1086), .A2(new_n725), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1083), .A2(new_n821), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n323), .A2(new_n823), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n331), .B1(new_n754), .B2(new_n201), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT119), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n760), .A2(new_n831), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT53), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n767), .A2(G159), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT54), .B(G143), .Z(new_n1096));
  AOI22_X1  g0896(.A1(new_n1090), .A2(KEYINPUT119), .B1(new_n751), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(G128), .ZN(new_n1098));
  INV_X1    g0898(.A(G132), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n747), .A2(new_n1098), .B1(new_n744), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G137), .B2(new_n764), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1092), .B(new_n1102), .C1(G125), .C2(new_n738), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n732), .A2(new_n502), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n769), .A2(G87), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n763), .A2(G68), .B1(G77), .B2(new_n767), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n331), .B1(new_n748), .B2(G283), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G116), .A2(new_n745), .B1(new_n738), .B2(G294), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1104), .B(new_n1109), .C1(G97), .C2(new_n751), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n777), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1088), .A2(new_n727), .A3(new_n1089), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n856), .B1(new_n889), .B2(new_n812), .ZN(new_n1113));
  AND4_X1   g0913(.A1(G330), .A2(new_n708), .A3(new_n856), .A4(new_n812), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1072), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1085), .B1(new_n1069), .B2(new_n856), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1115), .A2(new_n1116), .B1(new_n1117), .B2(new_n911), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n894), .A2(new_n890), .ZN(new_n1119));
  OR3_X1    g0919(.A1(new_n1086), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1117), .A2(new_n911), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n852), .A2(G330), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1081), .B1(new_n1122), .B2(new_n813), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n1116), .A3(new_n1070), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n438), .A2(new_n1122), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n893), .A2(new_n1126), .A3(new_n629), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT118), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n1086), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1120), .A2(new_n683), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n1128), .B2(new_n1086), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1087), .B(new_n1112), .C1(new_n1131), .C2(new_n1132), .ZN(G378));
  OAI21_X1  g0933(.A(new_n1127), .B1(new_n1086), .B2(new_n1118), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n723), .B1(new_n876), .B2(new_n885), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1136));
  NAND2_X1  g0936(.A1(new_n350), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n346), .A2(new_n347), .A3(new_n349), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n326), .A2(new_n859), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1137), .A2(new_n326), .A3(new_n859), .A4(new_n1139), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(new_n907), .A3(new_n909), .A4(new_n912), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n913), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1135), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1145), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n888), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1134), .A2(KEYINPUT57), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n683), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT121), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1150), .A2(new_n1148), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1134), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1151), .A2(KEYINPUT121), .A3(new_n683), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1155), .A2(new_n726), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1144), .A2(new_n821), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n222), .B1(new_n266), .B2(G41), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n769), .A2(new_n1096), .B1(G132), .B2(new_n764), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n748), .A2(G125), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n745), .A2(G128), .B1(new_n767), .B2(G150), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G137), .B2(new_n751), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT59), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n763), .A2(G159), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G33), .B1(new_n738), .B2(G124), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1170), .A2(new_n257), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1163), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1030), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n468), .A2(new_n750), .B1(new_n215), .B2(new_n732), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT120), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n763), .A2(G58), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(KEYINPUT120), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G116), .B2(new_n748), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n268), .B1(new_n737), .B2(new_n478), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n977), .B(new_n1183), .C1(G107), .C2(new_n745), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n257), .A3(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT58), .Z(new_n1186));
  OAI21_X1  g0986(.A(new_n777), .B1(new_n1175), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n823), .A2(new_n201), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1162), .A2(new_n727), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1161), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1160), .A2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1193), .A2(new_n1128), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n957), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT122), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1125), .A2(new_n726), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1081), .A2(new_n821), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n823), .A2(new_n210), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1179), .B(new_n331), .C1(new_n831), .C2(new_n750), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n769), .B2(G159), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n745), .A2(G137), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n748), .A2(G132), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1096), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1204), .A2(new_n732), .B1(new_n1098), .B2(new_n737), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G50), .B2(new_n767), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n760), .A2(new_n215), .B1(new_n755), .B2(new_n737), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT124), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n979), .A2(new_n268), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT123), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n747), .A2(new_n537), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1209), .A2(new_n1029), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n502), .B2(new_n750), .C1(new_n478), .C2(new_n744), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n732), .A2(new_n587), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1207), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n777), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1198), .A2(new_n727), .A3(new_n1199), .A4(new_n1217), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1197), .A2(KEYINPUT125), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT125), .B1(new_n1197), .B2(new_n1218), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1196), .A2(new_n1222), .ZN(G381));
  NOR2_X1   g1023(.A1(G375), .A2(G378), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n976), .A2(new_n1067), .A3(new_n1003), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G396), .A3(G393), .ZN(new_n1226));
  INV_X1    g1026(.A(G384), .ZN(new_n1227));
  INV_X1    g1027(.A(G381), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(G407));
  NAND2_X1  g1029(.A1(new_n659), .A2(G213), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT126), .Z(new_n1231));
  AOI21_X1  g1031(.A(new_n655), .B1(new_n1224), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(G407), .ZN(G409));
  XNOR2_X1  g1033(.A(G393), .B(new_n793), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1225), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1067), .B1(new_n976), .B2(new_n1003), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(G390), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1234), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1225), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1151), .A2(KEYINPUT121), .A3(new_n683), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT121), .B1(new_n1151), .B2(new_n683), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1134), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(G378), .B1(new_n1245), .B2(new_n1190), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1231), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n683), .B(new_n1249), .C1(new_n1194), .C2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1222), .A2(new_n1251), .A3(G384), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n1193), .B2(new_n1128), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1253), .A2(new_n688), .A3(new_n1248), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1227), .B1(new_n1254), .B2(new_n1221), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1161), .B(new_n1189), .C1(new_n1156), .C2(new_n958), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(G378), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1246), .A2(new_n1247), .A3(new_n1257), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1231), .B1(G375), .B2(G378), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1257), .A4(new_n1260), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1160), .B2(new_n1191), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1269), .A2(new_n1231), .A3(new_n1259), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1231), .A2(G2897), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1256), .B(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1267), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1241), .B1(new_n1266), .B2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1246), .A2(new_n1247), .A3(new_n1260), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT127), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1272), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1263), .A2(new_n1278), .A3(new_n1260), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1241), .B1(new_n1281), .B2(new_n1261), .ZN(new_n1282));
  NOR4_X1   g1082(.A1(new_n1269), .A2(new_n1231), .A3(new_n1256), .A4(new_n1259), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1283), .B2(KEYINPUT63), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1282), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1274), .A2(new_n1285), .ZN(G405));
  OR3_X1    g1086(.A1(new_n1224), .A2(new_n1257), .A3(new_n1269), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1241), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1257), .B1(new_n1224), .B2(new_n1269), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


