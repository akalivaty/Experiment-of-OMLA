//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1147, new_n1148, new_n1149,
    new_n1150;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT67), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(G137), .A3(new_n470), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n464), .A2(new_n465), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n466), .B1(new_n469), .B2(new_n468), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n470), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n484), .A2(G124), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n482), .A2(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n470), .A2(G138), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n466), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n466), .A2(G138), .A3(new_n470), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(new_n493), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n495), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n504), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(G88), .B1(G50), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n511), .A2(new_n512), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n516), .A2(G89), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT72), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n505), .A2(new_n525), .A3(new_n506), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n524), .A2(new_n526), .A3(G63), .A4(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n517), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n521), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND3_X1  g107(.A1(new_n524), .A2(new_n526), .A3(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n502), .B1(new_n533), .B2(new_n534), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n516), .A2(G90), .B1(G52), .B2(new_n517), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n524), .A2(new_n526), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n516), .A2(G81), .B1(G43), .B2(new_n517), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT74), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n515), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n517), .A2(KEYINPUT76), .A3(G53), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n559), .B(new_n565), .C1(new_n560), .C2(new_n561), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n516), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n522), .A2(new_n523), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n564), .A2(new_n566), .A3(new_n567), .A4(new_n572), .ZN(G299));
  OAI21_X1  g148(.A(new_n541), .B1(new_n539), .B2(KEYINPUT73), .ZN(new_n574));
  AOI211_X1 g149(.A(new_n537), .B(new_n502), .C1(new_n533), .C2(new_n534), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT77), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n538), .A2(new_n577), .A3(new_n540), .A4(new_n541), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G301));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n502), .B1(new_n545), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n517), .A2(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n515), .A2(new_n507), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n502), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n516), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n517), .A2(G48), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n517), .A2(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n585), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n545), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n596), .B1(new_n599), .B2(G651), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND3_X1  g179(.A1(new_n516), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n585), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n569), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n579), .B2(G868), .ZN(G284));
  XOR2_X1   g191(.A(G284), .B(KEYINPUT79), .Z(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(G168), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n618), .B2(G168), .ZN(G280));
  AND2_X1   g196(.A1(new_n609), .A2(new_n613), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n614), .A2(G559), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT80), .ZN(new_n626));
  MUX2_X1   g201(.A(new_n550), .B(new_n626), .S(G868), .Z(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n466), .A2(new_n475), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n484), .A2(G123), .B1(G135), .B2(new_n480), .ZN(new_n635));
  OAI221_X1 g210(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2096), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT82), .B(G2438), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n641), .B(new_n642), .Z(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n641), .B(new_n642), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n644), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  OAI21_X1  g234(.A(KEYINPUT83), .B1(new_n655), .B2(new_n657), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n651), .B(new_n654), .Z(new_n661));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n662), .A3(new_n656), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n659), .B1(new_n660), .B2(new_n663), .ZN(G401));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n632), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(new_n638), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(KEYINPUT84), .ZN(new_n680));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(KEYINPUT84), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n677), .A2(new_n678), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(new_n679), .ZN(new_n687));
  MUX2_X1   g262(.A(new_n687), .B(new_n686), .S(new_n682), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT85), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(G166), .A2(G16), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G16), .B2(G22), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n587), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n698), .A2(new_n699), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n700), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G6), .A2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G305), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT87), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  MUX2_X1   g293(.A(G24), .B(G290), .S(G16), .Z(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G1986), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n484), .A2(G119), .B1(G131), .B2(new_n480), .ZN(new_n721));
  OAI221_X1 g296(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n719), .B2(G1986), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n717), .A2(new_n718), .A3(new_n720), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n729), .A2(KEYINPUT88), .A3(KEYINPUT36), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G33), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G139), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n736), .B(new_n739), .C1(new_n470), .C2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT93), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n734), .B1(new_n743), .B2(new_n733), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G2072), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n701), .A2(G20), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT23), .Z(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G299), .B2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1956), .ZN(new_n749));
  NAND2_X1  g324(.A1(G286), .A2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n701), .A2(G21), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G4), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n622), .B2(G16), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n753), .A2(G1966), .B1(new_n755), .B2(G1348), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G1966), .B2(new_n753), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n745), .A2(new_n749), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n733), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n733), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G2090), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT99), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n551), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT89), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1341), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n758), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n761), .A2(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n733), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OAI22_X1  g349(.A1(G160), .A2(new_n733), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2084), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G1348), .B2(new_n755), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT30), .B(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  NAND2_X1  g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n778), .A2(new_n733), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n637), .B2(new_n733), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT97), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  NOR2_X1   g359(.A1(G27), .A2(G29), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G164), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n783), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n733), .A2(G26), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT28), .Z(new_n790));
  AOI22_X1  g365(.A1(new_n484), .A2(G128), .B1(G140), .B2(new_n480), .ZN(new_n791));
  NOR2_X1   g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT90), .Z(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n790), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G2078), .B2(new_n786), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n770), .A2(new_n777), .A3(new_n788), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G29), .A2(G32), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n480), .A2(G141), .ZN(new_n802));
  INV_X1    g377(.A(G105), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n476), .ZN(new_n804));
  NAND3_X1  g379(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT26), .Z(new_n806));
  INV_X1    g381(.A(G129), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n483), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n809));
  OR3_X1    g384(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n804), .B2(new_n808), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n801), .B1(new_n813), .B2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT27), .B(G1996), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G171), .A2(new_n701), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G5), .B2(new_n701), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n814), .A2(new_n816), .B1(new_n819), .B2(G1961), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(KEYINPUT98), .B2(new_n769), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n814), .A2(new_n816), .B1(new_n819), .B2(G1961), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n800), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n730), .A2(new_n732), .A3(new_n768), .A4(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n516), .A2(G93), .B1(G55), .B2(new_n517), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n524), .A2(new_n526), .A3(G67), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n826), .B(new_n827), .C1(new_n830), .C2(new_n502), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n502), .B1(new_n828), .B2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n517), .A2(G55), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n585), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT100), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n550), .A3(new_n836), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n548), .B(new_n549), .C1(new_n832), .C2(new_n835), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n622), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n846), .A2(new_n847), .A3(G860), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n831), .A2(new_n836), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n848), .A2(new_n851), .ZN(G145));
  NAND2_X1  g427(.A1(new_n495), .A2(new_n500), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n795), .B(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n810), .A2(new_n811), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n742), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n813), .A2(new_n742), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n855), .B(KEYINPUT96), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n743), .ZN(new_n861));
  INV_X1    g436(.A(new_n854), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n856), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n723), .B(new_n630), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n480), .A2(G142), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT103), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n484), .A2(G130), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n470), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n867), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n865), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n859), .A2(new_n863), .A3(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n637), .ZN(new_n877));
  XOR2_X1   g452(.A(G160), .B(KEYINPUT102), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(KEYINPUT104), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n859), .A2(new_n863), .A3(new_n883), .A4(new_n872), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n882), .A2(new_n874), .A3(new_n884), .A4(new_n879), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g463(.A(new_n849), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT105), .B1(new_n889), .B2(G868), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n566), .A2(new_n567), .A3(new_n572), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n891), .A2(new_n564), .A3(new_n609), .A4(new_n613), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n891), .A2(new_n564), .B1(new_n609), .B2(new_n613), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT41), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(new_n614), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n893), .A2(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n837), .A2(new_n838), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT101), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n837), .A2(new_n839), .A3(new_n838), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n626), .ZN(new_n905));
  MUX2_X1   g480(.A(new_n899), .B(new_n900), .S(new_n905), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT42), .ZN(new_n907));
  NAND2_X1  g482(.A1(G290), .A2(new_n710), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n602), .A2(G305), .A3(new_n603), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(G303), .B(G288), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n910), .B(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n618), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n910), .B(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n890), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n914), .A2(new_n918), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G295));
  AOI21_X1  g497(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G331));
  NAND3_X1  g498(.A1(new_n576), .A2(new_n578), .A3(G168), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n542), .B2(G168), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n576), .A2(new_n578), .A3(new_n925), .A4(G168), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n842), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n927), .B(new_n928), .C1(new_n841), .C2(new_n840), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n900), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n904), .B1(new_n928), .B2(new_n927), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n929), .A2(new_n842), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n899), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n930), .A2(KEYINPUT107), .A3(new_n931), .A4(new_n900), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n934), .A2(new_n937), .A3(new_n913), .A4(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n939), .A2(new_n886), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n898), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n896), .A2(new_n892), .A3(KEYINPUT108), .A4(new_n897), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n944), .A2(new_n895), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n935), .B2(new_n936), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n932), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n949), .B2(new_n916), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n930), .A2(new_n900), .A3(new_n931), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n946), .B1(new_n930), .B2(new_n931), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n916), .B(new_n942), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n941), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n934), .A2(new_n938), .A3(new_n937), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n916), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n940), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n956), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n940), .B2(new_n958), .ZN(new_n962));
  NOR2_X1   g537(.A1(KEYINPUT43), .A2(G37), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n939), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT110), .B1(new_n955), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n939), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n916), .B1(new_n951), .B2(new_n952), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n953), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n962), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n966), .A2(new_n969), .A3(new_n970), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n970), .B1(new_n966), .B2(new_n969), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT111), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n960), .B1(new_n974), .B2(new_n980), .ZN(G397));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n853), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G160), .A2(G40), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n984), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n813), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n795), .A2(G2067), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n791), .A2(new_n797), .A3(new_n794), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n987), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n986), .A2(G1996), .A3(new_n812), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT112), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT113), .Z(new_n997));
  XNOR2_X1  g572(.A(new_n723), .B(new_n725), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n987), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(G290), .B(G1986), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n986), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G168), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1003), .A2(KEYINPUT51), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n985), .B1(new_n983), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1966), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n983), .A2(KEYINPUT50), .ZN(new_n1011));
  AND2_X1   g586(.A1(G160), .A2(G40), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n853), .A2(new_n1013), .A3(new_n982), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G2084), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G8), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1004), .B1(new_n1019), .B2(KEYINPUT122), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1002), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT51), .B1(new_n1021), .B2(new_n1003), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1020), .A2(new_n1023), .B1(new_n1024), .B2(KEYINPUT121), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1024), .A2(KEYINPUT121), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1025), .A2(new_n1026), .B1(new_n1018), .B2(new_n1003), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1028));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n1008), .B2(G2078), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1006), .A2(new_n1007), .A3(KEYINPUT53), .A4(new_n784), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1030), .B(new_n1031), .C1(G1961), .C2(new_n1015), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1032), .A2(new_n579), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n579), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1028), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n984), .A2(new_n1012), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n587), .A2(G1976), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n587), .B2(G1976), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1002), .B1(new_n984), .B2(new_n1012), .ZN(new_n1042));
  INV_X1    g617(.A(G1981), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n590), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(G305), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI221_X1 g624(.A(new_n1039), .B1(new_n1038), .B2(new_n1041), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G2090), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1971), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G303), .A2(G8), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT55), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1057), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(G8), .C1(new_n1054), .C2(new_n1053), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1051), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1032), .A2(G171), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(KEYINPUT54), .C1(new_n579), .C2(new_n1032), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1035), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  OR3_X1    g639(.A1(new_n1027), .A2(new_n1064), .A3(KEYINPUT124), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT124), .B1(new_n1027), .B2(new_n1064), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1015), .A2(G1348), .B1(G2067), .B2(new_n1036), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1067), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n622), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1069), .B2(KEYINPUT60), .ZN(new_n1070));
  XOR2_X1   g645(.A(G299), .B(KEYINPUT57), .Z(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1015), .A2(G1956), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1006), .A2(new_n1007), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1075), .B(new_n1071), .C1(G1956), .C2(new_n1015), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1077), .A2(KEYINPUT61), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT61), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT58), .B(G1341), .Z(new_n1083));
  NAND3_X1  g658(.A1(new_n1036), .A2(KEYINPUT118), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n985), .B2(new_n983), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1084), .B(new_n1087), .C1(new_n1008), .C2(G1996), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n551), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1089), .B(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1081), .A2(new_n1082), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1082), .B1(new_n1081), .B2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1070), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1078), .A2(new_n1067), .A3(new_n622), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(new_n1077), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1065), .A2(new_n1066), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1019), .A2(G286), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(new_n1051), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT63), .B1(new_n1100), .B2(KEYINPUT116), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(KEYINPUT116), .A3(KEYINPUT63), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G305), .A2(G1981), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT115), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1107));
  OR2_X1    g682(.A1(G288), .A2(G1976), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1104), .B1(new_n1042), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1102), .A2(KEYINPUT117), .A3(new_n1103), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1101), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1061), .B(new_n1033), .C1(new_n1027), .C2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1027), .A2(new_n1115), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1111), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1001), .B1(new_n1098), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n997), .A2(new_n725), .A3(new_n722), .A4(new_n721), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n987), .B1(new_n1120), .B2(new_n991), .ZN(new_n1121));
  INV_X1    g696(.A(new_n992), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n986), .B1(new_n1122), .B2(new_n812), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n987), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT46), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n986), .B2(new_n988), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1123), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT47), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n987), .A2(G1986), .A3(G290), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT125), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT48), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1128), .B1(new_n999), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1119), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n1136));
  NOR2_X1   g710(.A1(G227), .A2(new_n462), .ZN(new_n1137));
  AND2_X1   g711(.A1(new_n663), .A2(new_n660), .ZN(new_n1138));
  OAI211_X1 g712(.A(new_n1136), .B(new_n1137), .C1(new_n1138), .C2(new_n659), .ZN(new_n1139));
  INV_X1    g713(.A(new_n1137), .ZN(new_n1140));
  OAI21_X1  g714(.A(KEYINPUT126), .B1(G401), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g715(.A(G229), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AND2_X1   g716(.A1(new_n887), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g717(.A1(new_n978), .A2(new_n1143), .A3(KEYINPUT127), .ZN(new_n1144));
  AOI21_X1  g718(.A(KEYINPUT127), .B1(new_n978), .B2(new_n1143), .ZN(new_n1145));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n1145), .ZN(G308));
  NAND2_X1  g720(.A1(new_n978), .A2(new_n1143), .ZN(new_n1147));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n1148));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g723(.A1(new_n978), .A2(new_n1143), .A3(KEYINPUT127), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1150), .ZN(G225));
endmodule


