

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595;

  NOR2_X1 U322 ( .A1(n550), .A2(n365), .ZN(n366) );
  XNOR2_X1 U323 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U324 ( .A(n493), .B(KEYINPUT100), .ZN(n494) );
  XNOR2_X1 U325 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U326 ( .A(n391), .B(n390), .Z(n525) );
  NOR2_X1 U327 ( .A1(n536), .A2(n392), .ZN(n395) );
  INV_X1 U328 ( .A(n406), .ZN(n407) );
  XNOR2_X1 U329 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U330 ( .A(G71GAT), .B(G57GAT), .ZN(n327) );
  XNOR2_X1 U331 ( .A(n353), .B(n330), .ZN(n332) );
  XNOR2_X1 U332 ( .A(n410), .B(n409), .ZN(n416) );
  INV_X1 U333 ( .A(G78GAT), .ZN(n356) );
  INV_X1 U334 ( .A(KEYINPUT37), .ZN(n493) );
  INV_X1 U335 ( .A(KEYINPUT110), .ZN(n362) );
  XNOR2_X1 U336 ( .A(n357), .B(n356), .ZN(n358) );
  INV_X1 U337 ( .A(KEYINPUT118), .ZN(n454) );
  NAND2_X1 U338 ( .A1(n453), .A2(n537), .ZN(n455) );
  XNOR2_X1 U339 ( .A(n495), .B(n494), .ZN(n522) );
  XNOR2_X1 U340 ( .A(n464), .B(KEYINPUT28), .ZN(n540) );
  XNOR2_X1 U341 ( .A(n341), .B(n390), .ZN(n584) );
  XNOR2_X1 U342 ( .A(n455), .B(n454), .ZN(n571) );
  INV_X1 U343 ( .A(n540), .ZN(n530) );
  XNOR2_X1 U344 ( .A(n456), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U345 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n291) );
  XNOR2_X1 U347 ( .A(G218GAT), .B(G92GAT), .ZN(n290) );
  XNOR2_X1 U348 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U349 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n293) );
  XNOR2_X1 U350 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n292) );
  XNOR2_X1 U351 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U352 ( .A(n295), .B(n294), .Z(n306) );
  XOR2_X1 U353 ( .A(G29GAT), .B(KEYINPUT67), .Z(n297) );
  XNOR2_X1 U354 ( .A(KEYINPUT7), .B(G43GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n299) );
  XOR2_X1 U356 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n298) );
  XOR2_X1 U357 ( .A(n299), .B(n298), .Z(n323) );
  INV_X1 U358 ( .A(n323), .ZN(n304) );
  XOR2_X1 U359 ( .A(G36GAT), .B(G190GAT), .Z(n377) );
  XNOR2_X1 U360 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n300), .B(G162GAT), .ZN(n405) );
  XOR2_X1 U362 ( .A(n377), .B(n405), .Z(n302) );
  NAND2_X1 U363 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U364 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U365 ( .A(n304), .B(n303), .Z(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U367 ( .A(n307), .B(KEYINPUT10), .Z(n310) );
  XNOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n308), .B(KEYINPUT71), .ZN(n331) );
  XNOR2_X1 U370 ( .A(G134GAT), .B(n331), .ZN(n309) );
  XOR2_X1 U371 ( .A(n310), .B(n309), .Z(n566) );
  INV_X1 U372 ( .A(n566), .ZN(n550) );
  XOR2_X1 U373 ( .A(G141GAT), .B(G22GAT), .Z(n312) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(G197GAT), .ZN(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n314) );
  XNOR2_X1 U377 ( .A(G15GAT), .B(G8GAT), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G36GAT), .Z(n316) );
  XOR2_X1 U380 ( .A(G113GAT), .B(G1GAT), .Z(n419) );
  XNOR2_X1 U381 ( .A(n419), .B(KEYINPUT29), .ZN(n315) );
  XNOR2_X1 U382 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U383 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U384 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U387 ( .A(n324), .B(n323), .Z(n581) );
  INV_X1 U388 ( .A(n581), .ZN(n555) );
  XOR2_X1 U389 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n326) );
  XNOR2_X1 U390 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n327), .B(KEYINPUT13), .ZN(n353) );
  AND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  INV_X1 U394 ( .A(KEYINPUT72), .ZN(n328) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n335) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n333), .B(G148GAT), .ZN(n406) );
  XNOR2_X1 U398 ( .A(G120GAT), .B(n406), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U401 ( .A(G92GAT), .B(KEYINPUT73), .Z(n339) );
  XNOR2_X1 U402 ( .A(G204GAT), .B(G64GAT), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U404 ( .A(G176GAT), .B(n340), .ZN(n390) );
  XNOR2_X1 U405 ( .A(KEYINPUT41), .B(n584), .ZN(n560) );
  NOR2_X1 U406 ( .A1(n555), .A2(n560), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n342), .B(KEYINPUT46), .ZN(n363) );
  XOR2_X1 U408 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n344) );
  XNOR2_X1 U409 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n343) );
  XNOR2_X1 U410 ( .A(n344), .B(n343), .ZN(n361) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(G183GAT), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n345), .B(G211GAT), .ZN(n381) );
  XOR2_X1 U413 ( .A(G22GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U414 ( .A(n381), .B(n401), .ZN(n349) );
  INV_X1 U415 ( .A(n349), .ZN(n347) );
  AND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  INV_X1 U417 ( .A(n348), .ZN(n346) );
  NAND2_X1 U418 ( .A1(n347), .A2(n346), .ZN(n351) );
  NAND2_X1 U419 ( .A1(n349), .A2(n348), .ZN(n350) );
  NAND2_X1 U420 ( .A1(n351), .A2(n350), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n352), .B(KEYINPUT12), .ZN(n355) );
  XOR2_X1 U422 ( .A(n353), .B(KEYINPUT78), .Z(n354) );
  XNOR2_X1 U423 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U424 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XNOR2_X1 U425 ( .A(G1GAT), .B(n439), .ZN(n357) );
  XOR2_X1 U426 ( .A(n361), .B(n360), .Z(n563) );
  XNOR2_X1 U427 ( .A(n563), .B(n362), .ZN(n546) );
  NOR2_X1 U428 ( .A1(n363), .A2(n546), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n364), .B(KEYINPUT111), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(KEYINPUT47), .ZN(n371) );
  XNOR2_X1 U431 ( .A(KEYINPUT36), .B(n566), .ZN(n592) );
  NOR2_X1 U432 ( .A1(n592), .A2(n563), .ZN(n367) );
  XOR2_X1 U433 ( .A(KEYINPUT45), .B(n367), .Z(n368) );
  NOR2_X1 U434 ( .A1(n584), .A2(n368), .ZN(n369) );
  NAND2_X1 U435 ( .A1(n369), .A2(n555), .ZN(n370) );
  NAND2_X1 U436 ( .A1(n371), .A2(n370), .ZN(n373) );
  XOR2_X1 U437 ( .A(KEYINPUT64), .B(KEYINPUT48), .Z(n372) );
  XNOR2_X1 U438 ( .A(n373), .B(n372), .ZN(n536) );
  XOR2_X1 U439 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n375) );
  XNOR2_X1 U440 ( .A(KEYINPUT92), .B(KEYINPUT90), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U442 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U443 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U445 ( .A(n381), .B(n380), .Z(n389) );
  XNOR2_X1 U446 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n382), .B(KEYINPUT19), .ZN(n383) );
  XOR2_X1 U448 ( .A(n383), .B(KEYINPUT82), .Z(n385) );
  XNOR2_X1 U449 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n450) );
  XOR2_X1 U451 ( .A(KEYINPUT21), .B(KEYINPUT84), .Z(n387) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(G218GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n414) );
  XNOR2_X1 U454 ( .A(n450), .B(n414), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n391) );
  INV_X1 U456 ( .A(n525), .ZN(n392) );
  INV_X1 U457 ( .A(n395), .ZN(n394) );
  INV_X1 U458 ( .A(KEYINPUT54), .ZN(n393) );
  NAND2_X1 U459 ( .A1(n394), .A2(n393), .ZN(n397) );
  NAND2_X1 U460 ( .A1(KEYINPUT54), .A2(n395), .ZN(n396) );
  NAND2_X1 U461 ( .A1(n397), .A2(n396), .ZN(n577) );
  XOR2_X1 U462 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n399) );
  XNOR2_X1 U463 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n403) );
  AND2_X1 U466 ( .A1(G228GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U468 ( .A(n404), .B(G211GAT), .Z(n410) );
  XNOR2_X1 U469 ( .A(n405), .B(KEYINPUT24), .ZN(n408) );
  XOR2_X1 U470 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n412) );
  XNOR2_X1 U471 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U473 ( .A(G141GAT), .B(n413), .Z(n423) );
  XNOR2_X1 U474 ( .A(n423), .B(n414), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n468) );
  XOR2_X1 U476 ( .A(G85GAT), .B(G162GAT), .Z(n421) );
  XOR2_X1 U477 ( .A(G120GAT), .B(KEYINPUT81), .Z(n418) );
  XNOR2_X1 U478 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n440) );
  XNOR2_X1 U480 ( .A(n419), .B(n440), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n436) );
  XOR2_X1 U483 ( .A(G155GAT), .B(G148GAT), .Z(n425) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G127GAT), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U486 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n427) );
  XNOR2_X1 U487 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U489 ( .A(n429), .B(n428), .Z(n434) );
  XOR2_X1 U490 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n431) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(KEYINPUT1), .B(n432), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U495 ( .A(n436), .B(n435), .Z(n576) );
  AND2_X1 U496 ( .A1(n468), .A2(n576), .ZN(n437) );
  NAND2_X1 U497 ( .A1(n577), .A2(n437), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n438), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT20), .Z(n444) );
  XNOR2_X1 U503 ( .A(G113GAT), .B(G183GAT), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U505 ( .A(n446), .B(n445), .Z(n452) );
  XOR2_X1 U506 ( .A(G71GAT), .B(G99GAT), .Z(n448) );
  XNOR2_X1 U507 ( .A(G43GAT), .B(G190GAT), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(n537) );
  NAND2_X1 U511 ( .A1(n550), .A2(n571), .ZN(n458) );
  XOR2_X1 U512 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n456) );
  INV_X1 U513 ( .A(n560), .ZN(n508) );
  NAND2_X1 U514 ( .A1(n571), .A2(n508), .ZN(n462) );
  XOR2_X1 U515 ( .A(G176GAT), .B(KEYINPUT120), .Z(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  NOR2_X1 U519 ( .A1(n584), .A2(n555), .ZN(n463) );
  XOR2_X1 U520 ( .A(n463), .B(KEYINPUT74), .Z(n496) );
  INV_X1 U521 ( .A(n576), .ZN(n523) );
  XNOR2_X1 U522 ( .A(n525), .B(KEYINPUT27), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n523), .A2(n470), .ZN(n535) );
  NOR2_X1 U524 ( .A1(n537), .A2(n535), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n468), .B(KEYINPUT66), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n465), .A2(n540), .ZN(n475) );
  NAND2_X1 U527 ( .A1(n537), .A2(n525), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n468), .A2(n466), .ZN(n467) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n467), .Z(n472) );
  NOR2_X1 U530 ( .A1(n468), .A2(n537), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(KEYINPUT26), .ZN(n578) );
  NAND2_X1 U532 ( .A1(n470), .A2(n578), .ZN(n471) );
  NAND2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n473), .A2(n576), .ZN(n474) );
  NAND2_X1 U535 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT94), .B(n476), .ZN(n492) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n478) );
  INV_X1 U538 ( .A(n563), .ZN(n587) );
  NAND2_X1 U539 ( .A1(n587), .A2(n566), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U541 ( .A1(n492), .A2(n479), .ZN(n509) );
  NOR2_X1 U542 ( .A1(n496), .A2(n509), .ZN(n489) );
  NAND2_X1 U543 ( .A1(n489), .A2(n523), .ZN(n483) );
  XOR2_X1 U544 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n481) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  XOR2_X1 U548 ( .A(G8GAT), .B(KEYINPUT97), .Z(n485) );
  NAND2_X1 U549 ( .A1(n489), .A2(n525), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U552 ( .A1(n489), .A2(n537), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n530), .A2(n489), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U557 ( .A1(n587), .A2(n592), .ZN(n491) );
  NAND2_X1 U558 ( .A1(n492), .A2(n491), .ZN(n495) );
  OR2_X1 U559 ( .A1(n496), .A2(n522), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT38), .ZN(n498) );
  XNOR2_X1 U561 ( .A(KEYINPUT101), .B(n498), .ZN(n506) );
  NAND2_X1 U562 ( .A1(n506), .A2(n523), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n499), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U566 ( .A1(n506), .A2(n525), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n506), .A2(n537), .ZN(n504) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U571 ( .A(G43GAT), .B(n505), .Z(G1330GAT) );
  NAND2_X1 U572 ( .A1(n530), .A2(n506), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n512) );
  NAND2_X1 U575 ( .A1(n555), .A2(n508), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n521), .A2(n509), .ZN(n510) );
  XOR2_X1 U577 ( .A(KEYINPUT103), .B(n510), .Z(n516) );
  NAND2_X1 U578 ( .A1(n516), .A2(n523), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U580 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NAND2_X1 U581 ( .A1(n525), .A2(n516), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n516), .A2(n537), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U586 ( .A1(n516), .A2(n530), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT105), .Z(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n523), .A2(n531), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  XOR2_X1 U593 ( .A(G92GAT), .B(KEYINPUT107), .Z(n527) );
  NAND2_X1 U594 ( .A1(n531), .A2(n525), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n531), .A2(n537), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n528), .B(KEYINPUT108), .ZN(n529) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n533) );
  NAND2_X1 U600 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n554) );
  NAND2_X1 U604 ( .A1(n537), .A2(n554), .ZN(n538) );
  XOR2_X1 U605 ( .A(KEYINPUT112), .B(n538), .Z(n539) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n545) );
  NOR2_X1 U607 ( .A1(n555), .A2(n545), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1340GAT) );
  NOR2_X1 U610 ( .A1(n560), .A2(n545), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n548) );
  INV_X1 U614 ( .A(n545), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n551), .A2(n546), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n578), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n555), .A2(n565), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n560), .A2(n565), .ZN(n561) );
  XOR2_X1 U629 ( .A(n562), .B(n561), .Z(G1345GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n565), .ZN(n564) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1347GAT) );
  XOR2_X1 U635 ( .A(G169GAT), .B(KEYINPUT119), .Z(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n581), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n571), .A2(n546), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n574) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(n575), .Z(n583) );
  AND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(KEYINPUT122), .B(n580), .ZN(n591) );
  INV_X1 U647 ( .A(n591), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n588), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U651 ( .A1(n588), .A2(n584), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  XOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT125), .Z(n590) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1354GAT) );
  XNOR2_X1 U656 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n594) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(G218GAT), .B(n595), .Z(G1355GAT) );
endmodule

