//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT70), .B(G50), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT71), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G45), .ZN(new_n251));
  AOI21_X1  g0051(.A(G1), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n254), .A3(G274), .ZN(new_n255));
  INV_X1    g0055(.A(G226), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n263), .A2(new_n264), .B1(new_n265), .B2(new_n261), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT72), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n254), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n260), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G169), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n274), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT73), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n278), .A2(new_n279), .A3(new_n216), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n279), .B1(new_n278), .B2(new_n216), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n204), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT76), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT8), .A2(G58), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT74), .B(G58), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(KEYINPUT8), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n217), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n290), .B1(G150), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n204), .A2(KEYINPUT76), .A3(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n285), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n282), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n217), .A3(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n278), .A2(new_n216), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n278), .A2(new_n279), .A3(new_n216), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n202), .B1(new_n257), .B2(G20), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n303), .A2(new_n304), .B1(new_n202), .B2(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n277), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT9), .B1(new_n297), .B2(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(new_n260), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n268), .B(KEYINPUT72), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n266), .B1(new_n311), .B2(G223), .ZN(new_n312));
  OAI211_X1 g0112(.A(G190), .B(new_n310), .C1(new_n312), .C2(new_n254), .ZN(new_n313));
  XOR2_X1   g0113(.A(KEYINPUT77), .B(G200), .Z(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n274), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n305), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n318), .A2(new_n293), .A3(new_n294), .A4(new_n285), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n319), .B2(new_n282), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n320), .A2(KEYINPUT78), .A3(KEYINPUT9), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT78), .B1(new_n320), .B2(KEYINPUT9), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT78), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n306), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n320), .A2(KEYINPUT78), .A3(KEYINPUT9), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(new_n316), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n308), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G33), .ZN(new_n334));
  INV_X1    g0134(.A(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(KEYINPUT81), .A3(KEYINPUT7), .A4(new_n217), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n261), .B2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(G20), .B1(new_n334), .B2(new_n336), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT81), .B1(new_n342), .B2(KEYINPUT7), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n201), .B1(new_n287), .B2(G68), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT82), .ZN(new_n347));
  INV_X1    g0147(.A(new_n291), .ZN(new_n348));
  INV_X1    g0148(.A(G159), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n291), .A2(KEYINPUT82), .A3(G159), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n346), .A2(G20), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n344), .A2(new_n352), .A3(KEYINPUT16), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n351), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n345), .B2(new_n217), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT83), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n335), .B2(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n333), .A2(KEYINPUT83), .A3(G33), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n336), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n339), .A2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n357), .B1(new_n363), .B2(new_n340), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n354), .B1(new_n356), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n353), .A2(new_n365), .A3(new_n282), .ZN(new_n366));
  INV_X1    g0166(.A(G232), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n255), .B1(new_n367), .B2(new_n259), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n256), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n261), .B(new_n369), .C1(G223), .C2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n372), .B2(new_n273), .ZN(new_n373));
  INV_X1    g0173(.A(G190), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G200), .B2(new_n373), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n257), .A2(G20), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n288), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n288), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n378), .A2(new_n303), .B1(new_n299), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n381));
  NAND4_X1  g0181(.A1(new_n366), .A2(new_n376), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(KEYINPUT86), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n382), .A2(KEYINPUT86), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n366), .A2(new_n376), .A3(new_n380), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT17), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n366), .A2(new_n380), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT84), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT84), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n366), .A2(new_n390), .A3(new_n380), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n373), .A2(G179), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n373), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT18), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n389), .A2(new_n397), .A3(new_n391), .A4(new_n394), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G244), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n255), .B1(new_n400), .B2(new_n259), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G107), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n263), .A2(new_n367), .B1(new_n403), .B2(new_n261), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n311), .B2(G238), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n402), .B1(new_n405), .B2(new_n254), .ZN(new_n406));
  INV_X1    g0206(.A(new_n314), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n303), .A2(G77), .A3(new_n377), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT8), .B(G58), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n410), .A2(new_n348), .B1(new_n217), .B2(new_n265), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n289), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n282), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n299), .A2(new_n265), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n409), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n408), .B(new_n416), .C1(new_n374), .C2(new_n406), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n406), .B2(new_n393), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n276), .B(new_n402), .C1(new_n405), .C2(new_n254), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT14), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n256), .A2(new_n262), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n367), .A2(G1698), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n334), .A2(new_n424), .A3(new_n336), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n273), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n254), .A2(G238), .A3(new_n258), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n255), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n423), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n254), .B1(new_n426), .B2(new_n427), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n434), .A2(new_n431), .A3(KEYINPUT13), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n422), .B(G169), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(new_n432), .A3(new_n423), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT13), .B1(new_n434), .B2(new_n431), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G179), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n422), .B1(new_n441), .B2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT80), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(G169), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n439), .A4(new_n436), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n357), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n265), .B2(new_n289), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n282), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT11), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT79), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n298), .A2(G1), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G20), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT12), .B1(new_n455), .B2(G68), .ZN(new_n456));
  OR3_X1    g0256(.A1(new_n455), .A2(KEYINPUT12), .A3(G68), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n357), .B1(new_n257), .B2(G20), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n456), .A2(new_n457), .B1(new_n303), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n452), .A2(KEYINPUT79), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n448), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n441), .A2(G200), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n462), .B(new_n465), .C1(new_n374), .C2(new_n441), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n421), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n332), .A2(new_n387), .A3(new_n399), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n333), .A2(G33), .ZN(new_n471));
  OAI21_X1  g0271(.A(G303), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n334), .A2(new_n336), .A3(G264), .A4(G1698), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n334), .A2(new_n336), .A3(G257), .A4(new_n262), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(new_n273), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT90), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(new_n250), .A3(KEYINPUT5), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT5), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(KEYINPUT90), .B2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n251), .A2(G1), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G270), .A3(new_n254), .ZN(new_n483));
  INV_X1    g0283(.A(G274), .ZN(new_n484));
  AND2_X1   g0284(.A1(G1), .A2(G13), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n253), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G200), .B1(new_n476), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT95), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n257), .A2(G33), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n455), .B(new_n491), .C1(new_n280), .C2(new_n281), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n303), .A2(KEYINPUT95), .A3(G116), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR4_X1   g0296(.A1(new_n298), .A2(new_n217), .A3(G1), .A4(G116), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n217), .ZN(new_n500));
  OR2_X1    g0300(.A1(KEYINPUT88), .A2(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(KEYINPUT88), .A2(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n503), .B2(new_n335), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n278), .A2(new_n216), .B1(G20), .B2(new_n493), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n498), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(KEYINPUT88), .A2(G97), .ZN(new_n508));
  NOR2_X1   g0308(.A1(KEYINPUT88), .A2(G97), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G33), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT20), .B(new_n505), .C1(new_n511), .C2(new_n500), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n497), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n483), .A2(new_n487), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n475), .A2(new_n273), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(G190), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n489), .A2(new_n496), .A3(new_n513), .A4(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT96), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n496), .A2(new_n513), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n393), .B1(new_n514), .B2(new_n515), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n514), .A2(G179), .A3(new_n515), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n519), .A2(KEYINPUT21), .A3(new_n520), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n454), .A2(G20), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT89), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n530), .B(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n529), .B2(new_n492), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  AND2_X1   g0334(.A1(G97), .A2(G107), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n206), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n403), .A2(KEYINPUT6), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n510), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT87), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n348), .B2(new_n265), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n291), .A2(KEYINPUT87), .A3(G77), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n538), .A2(G20), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n337), .A2(new_n217), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(new_n339), .B1(new_n361), .B2(new_n362), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n403), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n533), .B1(new_n545), .B2(new_n282), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n482), .A2(G257), .A3(new_n254), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n487), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n334), .A2(new_n336), .A3(G244), .A4(new_n262), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n499), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n548), .B1(new_n554), .B2(new_n273), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G169), .ZN(new_n556));
  AOI211_X1 g0356(.A(G179), .B(new_n548), .C1(new_n273), .C2(new_n554), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n546), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI211_X1 g0358(.A(G190), .B(new_n548), .C1(new_n273), .C2(new_n554), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n273), .ZN(new_n560));
  INV_X1    g0360(.A(new_n548), .ZN(new_n561));
  AOI21_X1  g0361(.A(G200), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n546), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT91), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n546), .B(new_n565), .C1(new_n559), .C2(new_n562), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n558), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n334), .A2(new_n336), .A3(new_n217), .A4(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT22), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT22), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n261), .A2(new_n570), .A3(new_n217), .A4(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G116), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(G20), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n217), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n403), .A2(KEYINPUT23), .A3(G20), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n572), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n573), .B1(new_n572), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n282), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n299), .A2(new_n403), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n583), .B(KEYINPUT25), .ZN(new_n584));
  INV_X1    g0384(.A(new_n492), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(G107), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n482), .A2(G264), .A3(new_n254), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n334), .A2(new_n336), .A3(G257), .A4(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n334), .A2(new_n336), .A3(G250), .A4(new_n262), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n254), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT97), .A4(new_n592), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n589), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n276), .A3(new_n487), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n594), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n273), .A3(new_n596), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(new_n487), .A3(new_n588), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n393), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n587), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(G200), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n597), .A2(G190), .A3(new_n487), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n582), .A4(new_n586), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n334), .A2(new_n336), .A3(G244), .A4(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n334), .A2(new_n336), .A3(G238), .A4(new_n262), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n574), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n273), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT92), .B1(new_n251), .B2(G1), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT92), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n257), .A3(G45), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n254), .A2(new_n611), .A3(new_n613), .A4(G250), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n254), .A2(G274), .A3(new_n481), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n276), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n273), .B2(new_n609), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(G169), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n334), .A2(new_n336), .A3(new_n217), .A4(G68), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n289), .B1(new_n501), .B2(new_n502), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n622), .B1(new_n623), .B2(KEYINPUT19), .ZN(new_n624));
  NOR2_X1   g0424(.A1(G87), .A2(G107), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n501), .A2(new_n502), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT19), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n217), .B1(new_n427), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n282), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n412), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(new_n455), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n303), .A2(new_n631), .A3(new_n491), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT93), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n627), .B1(new_n510), .B2(new_n289), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n626), .A2(new_n628), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(new_n622), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n632), .B1(new_n640), .B2(new_n282), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT93), .B1(new_n641), .B2(new_n634), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n621), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n610), .A2(new_n616), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n407), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n303), .A2(G87), .A3(new_n491), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(KEYINPUT94), .A3(new_n641), .A4(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT94), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n630), .A2(new_n633), .A3(new_n646), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n314), .B1(new_n610), .B2(new_n616), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n610), .A2(G190), .A3(new_n616), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n603), .A2(new_n606), .A3(new_n643), .A4(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n469), .A2(new_n528), .A3(new_n567), .A4(new_n654), .ZN(G372));
  NAND2_X1  g0455(.A1(new_n388), .A2(new_n394), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(new_n397), .ZN(new_n657));
  INV_X1    g0457(.A(new_n420), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n466), .A2(new_n658), .B1(new_n448), .B2(new_n463), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n386), .A2(KEYINPUT86), .A3(new_n382), .ZN(new_n660));
  INV_X1    g0460(.A(new_n383), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n657), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT102), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n324), .A2(new_n331), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT102), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n666), .B(new_n657), .C1(new_n659), .C2(new_n662), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n307), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n635), .A2(new_n636), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n641), .A2(KEYINPUT93), .A3(new_n634), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n620), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n652), .B1(new_n314), .B2(new_n619), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT98), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n641), .A2(new_n677), .A3(new_n646), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n671), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n650), .B1(G190), .B2(new_n619), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n641), .A2(new_n677), .A3(new_n646), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n641), .B2(new_n646), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n643), .A2(new_n684), .A3(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(new_n567), .A3(new_n606), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT100), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n603), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n603), .A2(new_n688), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n527), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n643), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT26), .B1(new_n686), .B2(new_n558), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n558), .A2(new_n643), .A3(new_n653), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n693), .A2(KEYINPUT101), .B1(KEYINPUT26), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT101), .ZN(new_n696));
  OR3_X1    g0496(.A1(new_n546), .A2(new_n556), .A3(new_n557), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n680), .B2(new_n685), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n698), .B2(KEYINPUT26), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n692), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n670), .B1(new_n468), .B2(new_n700), .ZN(G369));
  NAND2_X1  g0501(.A1(new_n454), .A2(new_n217), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G343), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n519), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n528), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n527), .A2(new_n519), .A3(new_n707), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n603), .A2(new_n606), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n587), .A2(new_n707), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n603), .A2(new_n706), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n689), .A2(new_n690), .A3(new_n706), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n713), .A2(new_n527), .A3(new_n706), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n720), .A2(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n210), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n626), .A2(G116), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n214), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n603), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n686), .A2(new_n567), .A3(new_n606), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT104), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n566), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n560), .A2(new_n374), .A3(new_n561), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G200), .B2(new_n555), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n565), .B1(new_n739), .B2(new_n546), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n697), .B(new_n606), .C1(new_n737), .C2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT104), .A3(new_n686), .A4(new_n733), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT103), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n643), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n674), .A2(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT26), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n558), .A2(new_n653), .A3(new_n643), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n674), .A2(new_n679), .A3(new_n671), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT99), .B1(new_n643), .B2(new_n684), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n558), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n750), .B1(new_n753), .B2(KEYINPUT26), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n736), .A2(new_n743), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n706), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT29), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n753), .A2(KEYINPUT101), .A3(new_n748), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n694), .A2(KEYINPUT26), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n699), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n751), .A2(new_n752), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n741), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n603), .B(new_n688), .ZN(new_n763));
  INV_X1    g0563(.A(new_n527), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n674), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT29), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n767), .A2(new_n768), .A3(new_n706), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G330), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n524), .A2(new_n555), .A3(new_n597), .A4(new_n619), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT30), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n514), .A2(new_n515), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n775), .A2(new_n644), .A3(new_n276), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n776), .A2(KEYINPUT30), .A3(new_n555), .A4(new_n597), .ZN(new_n777));
  INV_X1    g0577(.A(new_n555), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n619), .A2(G179), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n601), .A2(new_n778), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n774), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g0581(.A1(new_n781), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n782));
  AOI21_X1  g0582(.A(KEYINPUT31), .B1(new_n781), .B2(new_n707), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n528), .A2(new_n654), .A3(new_n567), .A4(new_n706), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n771), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n770), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n732), .B1(new_n787), .B2(G1), .ZN(G364));
  NOR2_X1   g0588(.A1(new_n298), .A2(G20), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n257), .B1(new_n789), .B2(G45), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n727), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G355), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n261), .A2(new_n210), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n794), .B1(G116), .B2(new_n210), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n244), .A2(new_n251), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n337), .A2(new_n210), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n251), .B2(new_n215), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n216), .B1(G20), .B2(new_n393), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n792), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n803), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n217), .A2(G179), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n407), .A2(G190), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n407), .A2(new_n374), .A3(new_n808), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G87), .A2(new_n810), .B1(new_n812), .B2(G107), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n217), .A2(new_n276), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G190), .A2(G200), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n261), .B1(new_n816), .B2(new_n265), .ZN(new_n817));
  INV_X1    g0617(.A(G200), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(G190), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n817), .B1(new_n287), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n808), .A2(new_n815), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n349), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n374), .A2(G179), .A3(G200), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n217), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n824), .A2(KEYINPUT32), .B1(new_n827), .B2(G97), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n813), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n814), .A2(G200), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n374), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(G190), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G50), .A2(new_n831), .B1(new_n832), .B2(G68), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n829), .B(new_n833), .C1(KEYINPUT32), .C2(new_n824), .ZN(new_n834));
  INV_X1    g0634(.A(new_n831), .ZN(new_n835));
  INV_X1    g0635(.A(G326), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n832), .ZN(new_n838));
  OR2_X1    g0638(.A1(KEYINPUT33), .A2(G317), .ZN(new_n839));
  NAND2_X1  g0639(.A1(KEYINPUT33), .A2(G317), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n837), .B(new_n841), .C1(G294), .C2(new_n827), .ZN(new_n842));
  INV_X1    g0642(.A(G322), .ZN(new_n843));
  INV_X1    g0643(.A(G311), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n819), .A2(new_n843), .B1(new_n816), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n822), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n261), .B(new_n845), .C1(G329), .C2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n809), .B(KEYINPUT105), .Z(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G303), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n812), .A2(G283), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n842), .A2(new_n847), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n807), .B1(new_n834), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n806), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n802), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n711), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT106), .Z(new_n856));
  INV_X1    g0656(.A(new_n712), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n792), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(G330), .B2(new_n711), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(G396));
  NOR2_X1   g0660(.A1(new_n700), .A2(new_n707), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n420), .A2(new_n707), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n417), .B1(new_n416), .B2(new_n706), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n420), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n421), .A2(new_n706), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n861), .A2(new_n864), .B1(new_n700), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n786), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n792), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  INV_X1    g0669(.A(G132), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n261), .B1(new_n822), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n811), .A2(new_n357), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(new_n287), .C2(new_n827), .ZN(new_n873));
  INV_X1    g0673(.A(new_n848), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n202), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT110), .ZN(new_n876));
  XNOR2_X1  g0676(.A(KEYINPUT109), .B(G143), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n816), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n820), .A2(new_n878), .B1(new_n879), .B2(G159), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  INV_X1    g0681(.A(G137), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n880), .B1(new_n838), .B2(new_n881), .C1(new_n882), .C2(new_n835), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT34), .Z(new_n884));
  NOR2_X1   g0684(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n261), .B1(new_n848), .B2(G107), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT108), .Z(new_n887));
  AOI22_X1  g0687(.A1(G97), .A2(new_n827), .B1(new_n831), .B2(G303), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT107), .B(G283), .Z(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n838), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n812), .A2(G87), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(G116), .A2(new_n879), .B1(new_n846), .B2(G311), .ZN(new_n893));
  INV_X1    g0693(.A(G294), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n819), .ZN(new_n895));
  NOR4_X1   g0695(.A1(new_n887), .A2(new_n890), .A3(new_n892), .A4(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n803), .B1(new_n885), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n792), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n803), .A2(new_n800), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n265), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n897), .B(new_n900), .C1(new_n801), .C2(new_n864), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n869), .A2(new_n901), .ZN(G384));
  OR2_X1    g0702(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n903), .A2(G116), .A3(new_n218), .A4(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT36), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n287), .A2(G68), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G77), .A3(new_n215), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n202), .A2(G68), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT111), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n257), .B(G13), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n656), .B(KEYINPUT18), .ZN(new_n913));
  INV_X1    g0713(.A(new_n705), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  INV_X1    g0716(.A(new_n380), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n353), .A2(new_n282), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n344), .A2(new_n352), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n354), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n394), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n385), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n921), .A2(new_n914), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT37), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n389), .A2(new_n391), .A3(new_n705), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT37), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n385), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n395), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n396), .A2(new_n660), .A3(new_n661), .A4(new_n398), .ZN(new_n930));
  AOI221_X4 g0730(.A(new_n916), .B1(new_n925), .B2(new_n929), .C1(new_n930), .C2(new_n924), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n924), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n925), .A2(new_n929), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT38), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n463), .A2(new_n707), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n464), .A2(new_n466), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n448), .A2(new_n463), .A3(new_n707), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n865), .B1(new_n760), .B2(new_n766), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n862), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n932), .A2(new_n933), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n916), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n932), .A2(KEYINPUT38), .A3(new_n933), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(KEYINPUT39), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n926), .A2(new_n385), .A3(new_n656), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT37), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n929), .ZN(new_n949));
  INV_X1    g0749(.A(new_n926), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n662), .B2(new_n913), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT38), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n946), .B1(new_n931), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n464), .A2(new_n707), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n915), .B1(new_n935), .B2(new_n941), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n669), .B1(new_n770), .B2(new_n469), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n784), .A2(new_n785), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n960), .A2(new_n939), .A3(KEYINPUT40), .A4(new_n864), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n395), .A2(new_n928), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n962), .A2(new_n926), .B1(new_n947), .B2(KEYINPUT37), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n926), .B1(new_n387), .B2(new_n657), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n916), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n961), .B1(new_n965), .B2(new_n944), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n960), .A2(new_n939), .A3(new_n864), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n931), .B2(new_n934), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT40), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n469), .A2(new_n960), .ZN(new_n972));
  OAI21_X1  g0772(.A(G330), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n972), .B2(new_n971), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n959), .A2(new_n974), .B1(new_n257), .B2(new_n789), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n959), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n912), .B1(new_n975), .B2(new_n976), .ZN(G367));
  INV_X1    g0777(.A(new_n239), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n804), .B1(new_n210), .B2(new_n412), .C1(new_n978), .C2(new_n797), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n261), .B1(new_n820), .B2(G303), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n822), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n838), .A2(new_n894), .B1(new_n835), .B2(new_n844), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n503), .C2(new_n812), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n809), .A2(new_n493), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(KEYINPUT46), .B2(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n826), .A2(new_n403), .B1(new_n889), .B2(new_n816), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT114), .ZN(new_n988));
  NAND2_X1  g0788(.A1(KEYINPUT46), .A2(G116), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n874), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n826), .A2(new_n357), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n831), .B2(new_n878), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n349), .B2(new_n838), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n819), .A2(new_n881), .B1(new_n816), .B2(new_n202), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n337), .B(new_n994), .C1(G137), .C2(new_n846), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n812), .A2(G77), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n810), .A2(new_n287), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n986), .A2(new_n990), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  OAI211_X1 g0800(.A(new_n792), .B(new_n979), .C1(new_n1000), .C2(new_n807), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n676), .A2(new_n678), .A3(new_n707), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n686), .A2(KEYINPUT112), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n643), .B2(new_n1002), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT112), .B1(new_n686), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1001), .B1(new_n1006), .B2(new_n802), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n546), .A2(new_n706), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n697), .B(new_n1009), .C1(new_n737), .C2(new_n740), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT113), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT113), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n567), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n558), .A2(new_n707), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1016), .A2(KEYINPUT44), .A3(new_n723), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT44), .B1(new_n1016), .B2(new_n723), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n724), .A2(new_n1015), .A3(KEYINPUT45), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT45), .B1(new_n724), .B2(new_n1015), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1017), .A2(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n719), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n720), .B1(new_n1019), .B2(new_n1020), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n764), .A2(new_n707), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n722), .B1(new_n717), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n712), .B(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n787), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n727), .B(KEYINPUT41), .Z(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n791), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n697), .B1(new_n1032), .B2(new_n603), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1015), .A2(new_n713), .A3(new_n1025), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1033), .A2(new_n706), .B1(new_n1034), .B2(KEYINPUT42), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(KEYINPUT42), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1006), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT43), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT43), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1006), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1041), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1043), .A2(new_n1044), .B1(new_n720), .B2(new_n1016), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1044), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n720), .A2(new_n1016), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n1042), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1008), .B1(new_n1031), .B2(new_n1049), .ZN(G387));
  AND2_X1   g0850(.A1(new_n235), .A2(G45), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1051), .A2(new_n797), .B1(new_n729), .B2(new_n794), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n410), .A2(G50), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g0854(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n729), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1052), .A2(new_n1056), .B1(new_n403), .B2(new_n726), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n792), .B1(new_n1057), .B2(new_n805), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n820), .A2(G317), .B1(new_n879), .B2(G303), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n838), .B2(new_n844), .C1(new_n843), .C2(new_n835), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n809), .A2(new_n894), .B1(new_n826), .B2(new_n889), .ZN(new_n1064));
  OR3_X1    g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n337), .B1(new_n836), .B2(new_n822), .C1(new_n811), .C2(new_n493), .ZN(new_n1069));
  OR3_X1    g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n826), .A2(new_n412), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n337), .B1(new_n846), .B2(G150), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n202), .B2(new_n819), .C1(new_n357), .C2(new_n816), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G159), .C2(new_n831), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G77), .A2(new_n810), .B1(new_n812), .B2(G97), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n379), .C2(new_n838), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n807), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1058), .B(new_n1077), .C1(new_n718), .C2(new_n802), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1027), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n791), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n787), .A2(new_n1079), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1079), .A2(new_n867), .A3(new_n757), .A4(new_n769), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n727), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(G393));
  NAND2_X1  g0884(.A1(new_n1024), .A2(new_n1082), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n787), .A2(new_n1079), .A3(new_n1023), .A4(new_n1022), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n727), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1024), .A2(KEYINPUT115), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT115), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1022), .A2(new_n1023), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n791), .A3(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n248), .A2(new_n797), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n804), .B1(new_n210), .B2(new_n510), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n792), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n826), .A2(new_n493), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n337), .B1(new_n822), .B2(new_n843), .C1(new_n894), .C2(new_n816), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G303), .C2(new_n832), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n403), .B2(new_n811), .C1(new_n809), .C2(new_n889), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G317), .A2(new_n831), .B1(new_n820), .B2(G311), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G150), .A2(new_n831), .B1(new_n820), .B2(G159), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n810), .A2(G68), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n261), .B1(new_n816), .B2(new_n410), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n846), .B2(new_n878), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n826), .A2(new_n265), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G50), .B2(new_n832), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n891), .A2(new_n1104), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1098), .A2(new_n1101), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1094), .B1(new_n1110), .B2(new_n803), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1015), .B2(new_n854), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1087), .A2(new_n1091), .A3(new_n1112), .ZN(G390));
  NAND2_X1  g0913(.A1(new_n469), .A2(new_n786), .ZN(new_n1114));
  AND4_X1   g0914(.A1(G330), .A2(new_n960), .A3(new_n939), .A4(new_n864), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n939), .B1(new_n786), .B2(new_n864), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(new_n940), .B2(new_n862), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n960), .A2(G330), .A3(new_n864), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n939), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n863), .A2(new_n420), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n755), .A2(new_n706), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n862), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n786), .A2(new_n864), .A3(new_n939), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n958), .A2(new_n1114), .A3(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n953), .A2(new_n945), .B1(new_n941), .B2(new_n956), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n956), .B1(new_n931), .B2(new_n952), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n939), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1128), .A2(new_n1131), .A3(new_n1115), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n941), .A2(new_n956), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n954), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1130), .A2(new_n939), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n955), .B1(new_n965), .B2(new_n944), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1124), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1127), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1115), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1140));
  AOI211_X1 g0940(.A(KEYINPUT29), .B(new_n707), .C1(new_n760), .C2(new_n766), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n768), .B1(new_n755), .B2(new_n706), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n469), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n670), .A3(new_n1114), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n945), .A2(new_n953), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1123), .B1(new_n700), .B2(new_n865), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n955), .B1(new_n1148), .B2(new_n939), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1137), .B(new_n1124), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1140), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1139), .A2(new_n727), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1140), .A2(new_n1150), .A3(new_n791), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n898), .B1(new_n379), .B2(new_n899), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n261), .B1(new_n816), .B2(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n838), .A2(new_n882), .B1(new_n349), .B2(new_n826), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(G125), .C2(new_n846), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G128), .A2(new_n831), .B1(new_n820), .B2(G132), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT117), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n809), .A2(new_n881), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n812), .A2(G50), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1158), .A2(new_n1160), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n848), .A2(G87), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n838), .A2(new_n403), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1107), .B(new_n1167), .C1(G283), .C2(new_n831), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n872), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n819), .A2(new_n493), .B1(new_n816), .B2(new_n510), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n261), .B(new_n1170), .C1(G294), .C2(new_n846), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .A4(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1165), .A2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1154), .B1(new_n807), .B2(new_n1173), .C1(new_n1147), .C2(new_n801), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1153), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1152), .A2(KEYINPUT119), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT119), .B1(new_n1152), .B2(new_n1175), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(G378));
  NAND2_X1  g0979(.A1(new_n306), .A2(new_n705), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT120), .Z(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n330), .B1(new_n329), .B2(new_n316), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n307), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1186), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n332), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n332), .A2(new_n1188), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1181), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n968), .A2(new_n969), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n966), .ZN(new_n1196));
  AND4_X1   g0996(.A1(G330), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1194), .B1(new_n970), .B2(G330), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n957), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n915), .B1(new_n941), .B2(new_n935), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n955), .B2(new_n1147), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(G330), .A3(new_n1196), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1194), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n970), .A2(G330), .A3(new_n1194), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1201), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1199), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n791), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n337), .B2(new_n250), .ZN(new_n1210));
  INV_X1    g1010(.A(G283), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n250), .B(new_n337), .C1(new_n822), .C2(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n819), .A2(new_n403), .B1(new_n816), .B2(new_n412), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n810), .C2(G77), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n831), .A2(G116), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n991), .B1(G97), .B2(new_n832), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n812), .A2(new_n287), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1210), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(G128), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n819), .A2(new_n1221), .B1(new_n816), .B2(new_n882), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G132), .B2(new_n832), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G150), .A2(new_n827), .B1(new_n831), .B2(G125), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n809), .C2(new_n1155), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n812), .A2(G159), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n846), .C2(G124), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1220), .B1(new_n1219), .B2(new_n1218), .C1(new_n1226), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n803), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n898), .B1(new_n202), .B2(new_n899), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n1194), .C2(new_n801), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1208), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT121), .B1(new_n958), .B2(new_n1114), .ZN(new_n1236));
  AND4_X1   g1036(.A1(KEYINPUT121), .A2(new_n1143), .A3(new_n670), .A4(new_n1114), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1151), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1207), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n728), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1151), .B2(new_n1238), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n957), .B(KEYINPUT122), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1199), .A2(new_n1206), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1235), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1208), .A2(new_n1234), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1199), .A2(new_n1206), .B1(new_n1151), .B2(new_n1238), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n727), .B1(new_n1252), .B2(KEYINPUT57), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT123), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1250), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G375));
  NAND2_X1  g1058(.A1(new_n848), .A2(G97), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n838), .A2(new_n493), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1071), .B(new_n1260), .C1(G294), .C2(new_n831), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n819), .A2(new_n1211), .B1(new_n816), .B2(new_n403), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n261), .B(new_n1262), .C1(G303), .C2(new_n846), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1259), .A2(new_n1261), .A3(new_n996), .A4(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n831), .A2(G132), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1266), .B1(new_n882), .B2(new_n819), .C1(new_n838), .C2(new_n1155), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n874), .A2(new_n349), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1265), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n261), .B1(new_n822), .B2(new_n1221), .C1(new_n881), .C2(new_n816), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(G50), .B2(new_n827), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1217), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1264), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n803), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n898), .B1(new_n357), .B2(new_n899), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(new_n939), .C2(new_n801), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1126), .B1(new_n958), .B2(new_n1114), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1146), .A2(new_n1278), .A3(new_n1029), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1277), .B(new_n1279), .C1(new_n791), .C2(new_n1126), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(G381));
  NAND2_X1  g1081(.A1(new_n1152), .A2(new_n1175), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OR2_X1    g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  INV_X1    g1084(.A(G390), .ZN(new_n1285));
  INV_X1    g1085(.A(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(G381), .A2(G387), .A3(new_n1284), .A4(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1257), .A2(new_n1283), .A3(new_n1288), .ZN(G407));
  INV_X1    g1089(.A(G213), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(G343), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1257), .A2(new_n1283), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(new_n1292), .A3(G213), .ZN(G409));
  OAI211_X1 g1093(.A(G390), .B(new_n1008), .C1(new_n1031), .C2(new_n1049), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT126), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(G393), .B(G396), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(new_n1285), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1295), .A2(new_n1296), .B1(new_n1297), .B2(new_n1294), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  AND4_X1   g1099(.A1(new_n1299), .A2(new_n1297), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1246), .A2(new_n791), .A3(new_n1244), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1302), .B(new_n1234), .C1(new_n1029), .C2(new_n1240), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1283), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT119), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1282), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1176), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1304), .B1(new_n1255), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1291), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1277), .B1(new_n1126), .B2(new_n791), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1278), .B1(KEYINPUT60), .B2(new_n1127), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT60), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n727), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1310), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  OR2_X1    g1114(.A1(new_n1314), .A2(new_n1286), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1286), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1308), .A2(new_n1309), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(KEYINPUT125), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT125), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1308), .A2(new_n1321), .A3(new_n1309), .A4(new_n1318), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT62), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1291), .A2(G2897), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1315), .A2(new_n1316), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1248), .A2(G378), .B1(new_n1283), .B2(new_n1303), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1327), .B1(new_n1328), .B2(new_n1291), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(new_n727), .A3(new_n1247), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1332), .A2(new_n1306), .A3(new_n1176), .A4(new_n1251), .ZN(new_n1333));
  AOI211_X1 g1133(.A(new_n1291), .B(new_n1317), .C1(new_n1333), .C2(new_n1304), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT62), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1329), .B(new_n1330), .C1(new_n1334), .C2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1301), .B1(new_n1323), .B2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(KEYINPUT127), .B1(new_n1301), .B2(KEYINPUT61), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT127), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1339), .B(new_n1330), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1329), .A2(new_n1338), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT63), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1320), .A2(new_n1322), .A3(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1334), .A2(KEYINPUT63), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1337), .A2(new_n1345), .ZN(G405));
  NAND3_X1  g1146(.A1(new_n1250), .A2(new_n1256), .A3(new_n1283), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1333), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1301), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1301), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1347), .A2(new_n1350), .A3(new_n1333), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1349), .A2(new_n1318), .A3(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1318), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(G402));
endmodule


