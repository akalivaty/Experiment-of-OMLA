//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT65), .A2(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT65), .A2(G146), .ZN(new_n191));
  OAI21_X1  g005(.A(G143), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT65), .B(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G143), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G146), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n202), .B1(new_n197), .B2(G143), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT66), .B(G143), .C1(new_n190), .C2(new_n191), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n206), .A2(KEYINPUT70), .A3(new_n207), .A4(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT66), .B1(new_n195), .B2(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n192), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n210), .A2(new_n207), .A3(G128), .A4(new_n204), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n199), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n198), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n204), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G125), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G224), .ZN(new_n226));
  XOR2_X1   g040(.A(new_n226), .B(KEYINPUT91), .Z(new_n227));
  AND3_X1   g041(.A1(new_n216), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n216), .B2(new_n224), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G107), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(G104), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT82), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n232), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G101), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT3), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n234), .A2(new_n231), .A3(KEYINPUT82), .A4(G104), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n236), .A2(new_n237), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G104), .ZN(new_n242));
  OAI22_X1  g056(.A1(new_n238), .A2(KEYINPUT3), .B1(new_n242), .B2(G107), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(G107), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n240), .A3(new_n239), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n246), .A3(KEYINPUT4), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT2), .B(G113), .Z(new_n248));
  XNOR2_X1  g062(.A(G116), .B(G119), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n255), .A2(G119), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(G113), .C1(KEYINPUT5), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n232), .A2(KEYINPUT83), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n244), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n233), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G101), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n248), .A2(new_n249), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n262), .A3(new_n241), .A4(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n253), .A2(KEYINPUT88), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT88), .B1(new_n253), .B2(new_n264), .ZN(new_n266));
  XOR2_X1   g080(.A(G110), .B(G122), .Z(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n253), .A2(new_n264), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n253), .A2(KEYINPUT88), .A3(new_n264), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n275), .A2(new_n271), .A3(new_n267), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT90), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n267), .A3(new_n276), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n253), .A2(new_n268), .A3(new_n264), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(KEYINPUT6), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT89), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n279), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n280), .ZN(new_n284));
  AOI221_X4 g098(.A(new_n230), .B1(new_n272), .B2(new_n278), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n280), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n216), .A2(new_n224), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n227), .A2(KEYINPUT7), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n262), .A2(new_n241), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n293), .A2(KEYINPUT92), .A3(new_n263), .A4(new_n257), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n267), .B(KEYINPUT8), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n257), .A2(new_n263), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT92), .B1(new_n296), .B2(new_n292), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n297), .B2(new_n264), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n287), .A2(new_n289), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n189), .B1(new_n285), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n283), .A2(new_n284), .ZN(new_n303));
  INV_X1    g117(.A(new_n230), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n272), .A2(new_n278), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n188), .A3(new_n300), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(KEYINPUT93), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n201), .A2(G128), .ZN(new_n309));
  INV_X1    g123(.A(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G143), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(G134), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT99), .B(KEYINPUT13), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(G134), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G116), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n231), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n314), .A2(G134), .A3(new_n309), .A4(new_n311), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n231), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n321), .A2(KEYINPUT100), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n255), .A2(KEYINPUT14), .A3(G122), .ZN(new_n323));
  INV_X1    g137(.A(new_n317), .ZN(new_n324));
  OAI211_X1 g138(.A(G107), .B(new_n323), .C1(new_n324), .C2(KEYINPUT14), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(KEYINPUT100), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n322), .A2(new_n313), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT9), .B(G234), .Z(new_n329));
  AND3_X1   g143(.A1(new_n329), .A2(G217), .A3(new_n225), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G902), .ZN(new_n332));
  INV_X1    g146(.A(G478), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT15), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n332), .B(KEYINPUT101), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(new_n334), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT72), .B(G237), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(G214), .A3(new_n225), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT95), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G143), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(G143), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n340), .A2(G214), .A3(new_n225), .A4(new_n344), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT18), .ZN(new_n349));
  INV_X1    g163(.A(G131), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n197), .ZN(new_n353));
  OAI21_X1  g167(.A(G140), .B1(new_n215), .B2(KEYINPUT79), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n353), .B1(new_n359), .B2(new_n195), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n346), .A2(KEYINPUT18), .A3(G131), .A4(new_n347), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n351), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(G113), .B(G122), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(new_n242), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT97), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n348), .A2(new_n350), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT17), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n346), .A2(G131), .A3(new_n347), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT16), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n358), .A2(KEYINPUT80), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n356), .A3(G125), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT80), .B1(new_n358), .B2(new_n370), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n195), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n371), .A2(G146), .A3(new_n372), .A4(new_n373), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n346), .A2(KEYINPUT17), .A3(G131), .A4(new_n347), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT98), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n362), .B(new_n365), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT96), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT19), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n352), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(KEYINPUT19), .B2(new_n358), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n197), .ZN(new_n385));
  INV_X1    g199(.A(new_n368), .ZN(new_n386));
  AOI21_X1  g200(.A(G131), .B1(new_n346), .B2(new_n347), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n376), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n362), .ZN(new_n389));
  INV_X1    g203(.A(new_n364), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n381), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT96), .B(new_n364), .C1(new_n388), .C2(new_n362), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n380), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G475), .ZN(new_n394));
  INV_X1    g208(.A(G902), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n393), .A2(new_n399), .A3(new_n394), .A4(new_n395), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n377), .A2(new_n379), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n351), .A2(new_n360), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n361), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n380), .B1(new_n404), .B2(new_n364), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n395), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G475), .ZN(new_n407));
  INV_X1    g221(.A(G952), .ZN(new_n408));
  AOI211_X1 g222(.A(G953), .B(new_n408), .C1(G234), .C2(G237), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT21), .B(G898), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT102), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n395), .B(new_n225), .C1(G234), .C2(G237), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AND4_X1   g229(.A1(new_n339), .A2(new_n401), .A3(new_n407), .A4(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n189), .C1(new_n285), .C2(new_n301), .ZN(new_n418));
  AND4_X1   g232(.A1(new_n187), .A2(new_n308), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n223), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n420), .A2(new_n252), .A3(new_n247), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n207), .B1(G143), .B2(new_n195), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n222), .B1(new_n310), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n211), .A2(new_n212), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n211), .A2(new_n212), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n293), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n430));
  INV_X1    g244(.A(G134), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(G137), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT11), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(G137), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT11), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n430), .B(new_n435), .C1(new_n431), .C2(G137), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G131), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n433), .A2(new_n350), .A3(new_n434), .A4(new_n436), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n208), .A2(new_n213), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n194), .A2(new_n198), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n428), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(new_n293), .ZN(new_n445));
  NOR4_X1   g259(.A1(new_n214), .A2(KEYINPUT84), .A3(new_n428), .A4(new_n292), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n429), .B(new_n440), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G140), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n225), .A2(G227), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n438), .A2(new_n439), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n443), .B1(new_n424), .B2(new_n425), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n293), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n292), .B1(new_n442), .B2(new_n423), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT12), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n214), .A2(new_n292), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n427), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n451), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n447), .A2(new_n450), .A3(new_n456), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT86), .ZN(new_n462));
  INV_X1    g276(.A(new_n450), .ZN(new_n463));
  INV_X1    g277(.A(new_n447), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n452), .A2(KEYINPUT10), .A3(new_n293), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT84), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n452), .A2(new_n441), .A3(KEYINPUT10), .A4(new_n293), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n440), .B1(new_n468), .B2(new_n429), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n463), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n459), .B1(new_n458), .B2(new_n451), .ZN(new_n471));
  AOI211_X1 g285(.A(KEYINPUT12), .B(new_n440), .C1(new_n427), .C2(new_n457), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n447), .A4(new_n450), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n462), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT85), .B(G469), .Z(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n395), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n450), .B1(new_n464), .B2(new_n469), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n447), .A3(new_n463), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G469), .B1(new_n481), .B2(G902), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n329), .ZN(new_n484));
  OAI21_X1  g298(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n485), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n478), .B2(new_n482), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT87), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n419), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT103), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n375), .A2(new_n376), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n310), .A2(G119), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT23), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n310), .A2(KEYINPUT23), .A3(G119), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n498), .B(new_n499), .C1(G119), .C2(new_n310), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G110), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT78), .B1(new_n310), .B2(G119), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT24), .B(G110), .Z(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n495), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  OAI22_X1  g322(.A1(new_n505), .A2(new_n506), .B1(new_n500), .B2(G110), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n376), .A2(new_n509), .A3(new_n353), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n511), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n395), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT25), .Z(new_n517));
  INV_X1    g331(.A(G234), .ZN(new_n518));
  OAI21_X1  g332(.A(G217), .B1(new_n518), .B2(G902), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n519), .B(KEYINPUT77), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n395), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n521), .B(KEYINPUT81), .Z(new_n522));
  AOI22_X1  g336(.A1(new_n517), .A2(new_n520), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n431), .B2(G137), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n434), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n526), .A2(new_n431), .A3(G137), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n439), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT69), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(KEYINPUT71), .A3(new_n534), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n452), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n250), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n420), .A2(new_n451), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT28), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT75), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT75), .B1(new_n542), .B2(new_n543), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n440), .A2(new_n223), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n532), .A2(new_n534), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n452), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT73), .B1(new_n550), .B2(new_n540), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n541), .B1(new_n214), .B2(new_n535), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n250), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n542), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT28), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n555), .B2(KEYINPUT28), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n547), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n340), .A2(G210), .A3(new_n225), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n237), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n561), .B(new_n562), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT31), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n566));
  NAND2_X1  g380(.A1(new_n552), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n539), .A2(new_n541), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n250), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n542), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n565), .B1(new_n571), .B2(new_n564), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n570), .A2(KEYINPUT31), .A3(new_n542), .A4(new_n563), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n559), .A2(new_n564), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT76), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n573), .ZN(new_n579));
  INV_X1    g393(.A(new_n546), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n544), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n555), .A2(KEYINPUT28), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT74), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT28), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n579), .B1(new_n585), .B2(new_n563), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT76), .B1(new_n586), .B2(new_n576), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n525), .B1(new_n578), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n547), .B(new_n563), .C1(new_n557), .C2(new_n558), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n571), .A2(new_n564), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n568), .B(new_n540), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n543), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n581), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n564), .A2(new_n590), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n559), .A2(new_n564), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n577), .B1(new_n599), .B2(new_n579), .ZN(new_n600));
  AOI22_X1  g414(.A1(G472), .A2(new_n598), .B1(new_n600), .B2(KEYINPUT32), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n524), .B1(new_n588), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n419), .A2(new_n488), .A3(KEYINPUT103), .A4(new_n491), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n494), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n488), .A2(new_n491), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n575), .B1(new_n574), .B2(new_n577), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n586), .A2(KEYINPUT76), .A3(new_n576), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G472), .B1(new_n574), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n606), .A2(new_n611), .A3(new_n524), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n306), .A2(new_n188), .A3(new_n300), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n188), .B1(new_n306), .B2(new_n300), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT104), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n306), .A2(KEYINPUT104), .A3(new_n188), .A4(new_n300), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n187), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n613), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n331), .A2(KEYINPUT33), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n620), .A2(KEYINPUT106), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(KEYINPUT106), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n331), .A2(KEYINPUT33), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n623), .A2(KEYINPUT107), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(KEYINPUT107), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n621), .A2(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n333), .A2(G902), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n626), .A2(new_n627), .B1(new_n333), .B2(new_n338), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n394), .B1(new_n405), .B2(new_n395), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n398), .B2(new_n400), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n302), .A2(new_n632), .A3(new_n307), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n633), .A2(KEYINPUT105), .A3(new_n187), .A4(new_n617), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n415), .A2(new_n619), .A3(new_n631), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n612), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  OR2_X1    g452(.A1(new_n396), .A2(new_n397), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n629), .B1(new_n639), .B2(new_n398), .ZN(new_n640));
  INV_X1    g454(.A(new_n339), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n619), .A2(new_n415), .A3(new_n634), .A4(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n643), .A2(KEYINPUT108), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(KEYINPUT108), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n612), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  INV_X1    g462(.A(new_n611), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n517), .A2(new_n520), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT36), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n514), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT109), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n511), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n522), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n494), .A2(new_n603), .A3(new_n649), .A4(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AND3_X1   g473(.A1(new_n619), .A2(new_n634), .A3(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n588), .A2(new_n601), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n490), .B(new_n487), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n409), .B1(new_n413), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n642), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XNOR2_X1  g482(.A(new_n664), .B(KEYINPUT39), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n308), .A2(new_n418), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT38), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n630), .A2(new_n339), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n187), .ZN(new_n678));
  INV_X1    g492(.A(new_n656), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n586), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n571), .A2(new_n563), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n593), .A2(new_n564), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n395), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G472), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n588), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n679), .B(new_n685), .C1(new_n671), .C2(KEYINPUT40), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n677), .A2(new_n678), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n201), .ZN(G45));
  NOR3_X1   g502(.A1(new_n628), .A2(new_n630), .A3(new_n664), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  INV_X1    g505(.A(G469), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n476), .B2(new_n395), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n485), .A3(new_n478), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n524), .B(new_n695), .C1(new_n588), .C2(new_n601), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n635), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  OAI21_X1  g513(.A(new_n696), .B1(new_n644), .B2(new_n645), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(new_n478), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n702), .A2(new_n693), .A3(new_n489), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n660), .A2(new_n661), .A3(new_n416), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND4_X1  g519(.A1(new_n619), .A2(new_n415), .A3(new_n634), .A4(new_n676), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n579), .B1(new_n595), .B2(new_n563), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n576), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n703), .A2(new_n610), .A3(new_n523), .A4(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(G122), .Z(G24));
  NAND2_X1  g525(.A1(new_n610), .A2(new_n708), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n660), .A2(new_n689), .A3(new_n703), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  AND3_X1   g529(.A1(new_n673), .A2(new_n490), .A3(new_n187), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n631), .A2(new_n665), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n661), .A2(new_n523), .A3(new_n716), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n598), .A2(G472), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n525), .B1(new_n574), .B2(new_n577), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n680), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n523), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n689), .A2(new_n673), .A3(new_n490), .A4(new_n187), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT42), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n719), .A2(new_n725), .A3(KEYINPUT110), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT110), .B1(new_n719), .B2(new_n725), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n350), .ZN(G33));
  AND2_X1   g543(.A1(new_n602), .A2(new_n716), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(new_n666), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n431), .ZN(G36));
  NAND2_X1  g546(.A1(new_n673), .A2(new_n187), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n481), .B(KEYINPUT45), .Z(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G469), .ZN(new_n735));
  NAND2_X1  g549(.A1(G469), .A2(G902), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT46), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n702), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n489), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n401), .A2(new_n407), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n628), .A2(KEYINPUT43), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(KEYINPUT111), .ZN(new_n743));
  INV_X1    g557(.A(new_n628), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n742), .B1(new_n745), .B2(KEYINPUT43), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n746), .A2(new_n611), .A3(new_n656), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n740), .B(new_n670), .C1(KEYINPUT44), .C2(new_n747), .ZN(new_n748));
  AOI211_X1 g562(.A(new_n733), .B(new_n748), .C1(KEYINPUT44), .C2(new_n747), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT112), .B(G137), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G39));
  OR2_X1    g565(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n661), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n733), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n524), .A3(new_n689), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  INV_X1    g571(.A(new_n409), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n712), .A2(new_n524), .A3(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n746), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n703), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n678), .A3(new_n674), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT50), .Z(new_n763));
  INV_X1    g577(.A(new_n685), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n733), .A2(new_n758), .A3(new_n695), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n523), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT117), .Z(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n630), .A3(new_n628), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n694), .A2(new_n478), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n752), .B(new_n753), .C1(new_n485), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n755), .A3(new_n760), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n746), .A2(new_n765), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n656), .A3(new_n713), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n763), .A2(new_n768), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n773), .B2(KEYINPUT118), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n225), .A2(G952), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n761), .A2(new_n619), .A3(new_n634), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n779), .B(new_n780), .C1(new_n631), .C2(new_n767), .ZN(new_n781));
  INV_X1    g595(.A(new_n723), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n774), .A2(KEYINPUT119), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT48), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT119), .B1(new_n774), .B2(new_n782), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n784), .B(new_n785), .Z(new_n786));
  AND3_X1   g600(.A1(new_n781), .A2(KEYINPUT120), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT120), .B1(new_n781), .B2(new_n786), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n778), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n776), .A2(new_n777), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n630), .A2(new_n641), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n628), .B2(new_n630), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n793), .A2(new_n678), .A3(new_n673), .A4(new_n414), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n612), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n657), .A2(new_n604), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n657), .A2(new_n795), .A3(new_n604), .A4(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n710), .B1(new_n696), .B2(new_n635), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n700), .A2(new_n801), .A3(new_n704), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n728), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n661), .A2(new_n662), .A3(new_n339), .A4(new_n640), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n713), .A2(new_n490), .A3(new_n631), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n679), .B(new_n733), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n731), .B1(new_n806), .B2(new_n665), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n619), .A2(new_n634), .A3(new_n676), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n486), .A2(new_n664), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n685), .A2(new_n808), .A3(new_n679), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n667), .A3(new_n690), .A4(new_n714), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT32), .B1(new_n607), .B2(new_n608), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n720), .A2(new_n680), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n606), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n660), .C1(new_n666), .C2(new_n689), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT52), .A3(new_n714), .A4(new_n810), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n800), .A2(new_n803), .A3(new_n807), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n822), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(KEYINPUT115), .A3(new_n822), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n719), .A2(new_n725), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n830), .A2(new_n800), .A3(new_n807), .A4(new_n820), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n802), .A2(new_n822), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(KEYINPUT116), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n800), .A2(new_n820), .A3(new_n807), .A4(new_n830), .ZN(new_n835));
  INV_X1    g649(.A(new_n832), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n829), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n789), .A2(new_n790), .A3(new_n824), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(G952), .B2(G953), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n675), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n745), .A2(new_n524), .A3(new_n489), .A4(new_n678), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n844), .A2(new_n764), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n842), .A2(new_n847), .ZN(G75));
  AOI21_X1  g662(.A(new_n395), .B1(new_n829), .B2(new_n838), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n849), .B2(G210), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n303), .A2(new_n305), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(new_n304), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT55), .Z(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(KEYINPUT56), .B(new_n853), .C1(new_n849), .C2(G210), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n225), .A2(G952), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G51));
  AOI21_X1  g672(.A(KEYINPUT116), .B1(new_n831), .B2(new_n832), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n835), .A2(new_n834), .A3(new_n836), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n821), .A2(KEYINPUT115), .A3(new_n822), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT115), .B1(new_n821), .B2(new_n822), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n859), .A2(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n840), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n736), .B(KEYINPUT57), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n476), .B(KEYINPUT121), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n849), .A2(G469), .A3(new_n734), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n857), .B1(new_n869), .B2(new_n870), .ZN(G54));
  NAND4_X1  g685(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n873));
  INV_X1    g687(.A(new_n393), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n857), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(G60));
  NAND2_X1  g693(.A1(G478), .A2(G902), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT59), .Z(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n840), .B2(new_n824), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n876), .B1(new_n882), .B2(new_n626), .ZN(new_n883));
  INV_X1    g697(.A(new_n626), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n881), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT123), .B1(new_n865), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n887));
  INV_X1    g701(.A(new_n885), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n887), .B(new_n888), .C1(new_n864), .C2(new_n840), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n883), .A2(new_n886), .A3(new_n889), .ZN(G63));
  NAND2_X1  g704(.A1(G217), .A2(G902), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT60), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n863), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n515), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n857), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n863), .A2(new_n654), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT61), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n896), .B(new_n897), .C1(new_n899), .C2(KEYINPUT61), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G66));
  AOI21_X1  g717(.A(new_n802), .B1(new_n798), .B2(new_n799), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(G953), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT126), .Z(new_n906));
  AOI21_X1  g720(.A(new_n225), .B1(new_n411), .B2(G224), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n851), .B1(G898), .B2(new_n225), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n908), .B(new_n909), .Z(G69));
  NAND2_X1  g724(.A1(new_n818), .A2(new_n714), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n756), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n728), .ZN(new_n914));
  INV_X1    g728(.A(new_n731), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n740), .A2(new_n670), .A3(new_n808), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n723), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n749), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n913), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT127), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n913), .A2(new_n918), .A3(new_n921), .A4(new_n914), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n225), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(new_n384), .Z(new_n925));
  OAI21_X1  g739(.A(G953), .B1(new_n663), .B2(G227), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n925), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n671), .A2(new_n733), .A3(new_n793), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n749), .B1(new_n602), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n225), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n687), .A2(new_n911), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n756), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n931), .A2(new_n934), .B1(new_n663), .B2(new_n926), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n927), .B1(new_n928), .B2(new_n935), .ZN(G72));
  NOR2_X1   g750(.A1(new_n571), .A2(new_n563), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n920), .A2(new_n904), .A3(new_n922), .ZN(new_n939));
  NAND2_X1  g753(.A1(G472), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT63), .Z(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n930), .A2(new_n904), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(new_n934), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n681), .B1(new_n944), .B2(new_n941), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n681), .A2(new_n823), .A3(new_n941), .A4(new_n938), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n942), .A2(new_n945), .A3(new_n857), .A4(new_n946), .ZN(G57));
endmodule


