//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT68), .Z(G261));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n455), .A2(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(G2104), .ZN(new_n469));
  OAI22_X1  g044(.A1(new_n466), .A2(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n476), .A2(new_n478), .A3(new_n465), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT72), .Z(new_n484));
  NAND2_X1  g059(.A1(new_n464), .A2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT71), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n488), .A2(KEYINPUT73), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(KEYINPUT73), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n476), .A2(new_n478), .A3(G126), .A4(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n476), .A2(new_n478), .A3(G138), .A4(new_n465), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n464), .A2(new_n499), .A3(G138), .A4(new_n465), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  XOR2_X1   g076(.A(KEYINPUT74), .B(G651), .Z(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT78), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n502), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT75), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT74), .B(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n519), .B(KEYINPUT6), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n503), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(G50), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n523), .B2(G50), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n514), .B1(new_n502), .B2(KEYINPUT6), .ZN(new_n529));
  NOR3_X1   g104(.A1(new_n516), .A2(KEYINPUT75), .A3(new_n517), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n508), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT77), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(G543), .B1(new_n529), .B2(new_n530), .ZN(new_n535));
  INV_X1    g110(.A(G50), .ZN(new_n536));
  OAI21_X1  g111(.A(KEYINPUT76), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n533), .B1(new_n537), .B2(new_n525), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n512), .B1(new_n534), .B2(new_n540), .ZN(G166));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT7), .Z(new_n543));
  AOI21_X1  g118(.A(new_n507), .B1(new_n518), .B2(new_n522), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(G89), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n523), .A2(G51), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n502), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n544), .A2(G90), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n523), .A2(G52), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n502), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n544), .A2(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n523), .A2(G43), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT79), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n535), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n523), .A2(new_n571), .A3(G53), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n507), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT80), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G91), .B2(new_n544), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(new_n512), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n538), .A2(new_n539), .ZN(new_n581));
  AOI211_X1 g156(.A(KEYINPUT77), .B(new_n533), .C1(new_n537), .C2(new_n525), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(G303));
  NAND2_X1  g158(.A1(new_n544), .A2(G87), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT82), .B1(new_n535), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n523), .A2(new_n590), .A3(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(G288));
  AOI22_X1  g168(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n502), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n523), .A2(G48), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n544), .A2(G86), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n502), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n544), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n523), .A2(G47), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n531), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n507), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n523), .A2(G54), .B1(G651), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT10), .B1(new_n531), .B2(new_n605), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n606), .A2(KEYINPUT83), .A3(new_n610), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n604), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n604), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  XNOR2_X1  g197(.A(G280), .B(KEYINPUT84), .ZN(G297));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n560), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n616), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g205(.A1(new_n479), .A2(G135), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G111), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G2105), .ZN(new_n634));
  AOI211_X1 g209(.A(new_n631), .B(new_n634), .C1(new_n486), .C2(G123), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT85), .B(G2438), .Z(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G14), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n660), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n662), .B1(new_n661), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n665), .B(new_n668), .Z(G227));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n680), .B(new_n681), .C1(new_n679), .C2(new_n678), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  NAND3_X1  g265(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT25), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n479), .A2(G139), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n692), .B(new_n693), .C1(new_n465), .C2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G33), .B(new_n695), .S(G29), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2072), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT30), .B(G28), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(G26), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n486), .A2(G128), .B1(G140), .B2(new_n479), .ZN(new_n704));
  OR2_X1    g279(.A1(G104), .A2(G2105), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n705), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n707), .B2(G29), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G2067), .ZN(new_n709));
  OR2_X1    g284(.A1(KEYINPUT24), .A2(G34), .ZN(new_n710));
  NAND2_X1  g285(.A1(KEYINPUT24), .A2(G34), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(new_n698), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G160), .B2(new_n698), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2084), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT92), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n700), .A2(new_n709), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n489), .A2(G29), .A3(new_n490), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n718));
  INV_X1    g293(.A(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G29), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n698), .A2(KEYINPUT94), .A3(G35), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n717), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  INV_X1    g298(.A(G2090), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT29), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n717), .A2(new_n725), .A3(new_n720), .A4(new_n721), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT95), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n723), .A2(KEYINPUT95), .A3(new_n724), .A4(new_n726), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n716), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n724), .B1(new_n723), .B2(new_n726), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT96), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n734), .A2(KEYINPUT23), .A3(G20), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT23), .ZN(new_n736));
  INV_X1    g311(.A(G20), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G16), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n738), .C1(new_n621), .C2(new_n734), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  OR3_X1    g315(.A1(new_n732), .A2(new_n733), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G19), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n561), .B2(G16), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G1341), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G21), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G168), .B2(G16), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G1966), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n479), .A2(G141), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  INV_X1    g326(.A(G105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n751), .C1(new_n752), .C2(new_n469), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G129), .B2(new_n486), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  AOI211_X1 g331(.A(new_n744), .B(new_n747), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n733), .B1(new_n732), .B2(new_n740), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n731), .A2(new_n741), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n746), .A2(G1966), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n734), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n734), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT31), .B(G11), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n755), .B2(new_n756), .ZN(new_n767));
  NOR2_X1   g342(.A1(G27), .A2(G29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G164), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2078), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n743), .A2(G1341), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n761), .A2(new_n765), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n759), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n734), .A2(G4), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n617), .B2(new_n734), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT90), .B(G1348), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT34), .ZN(new_n780));
  INV_X1    g355(.A(G305), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G6), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT32), .B(G1981), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n592), .A2(new_n587), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n584), .B(KEYINPUT81), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G16), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT33), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G16), .B2(G23), .ZN(new_n792));
  OR3_X1    g367(.A1(new_n791), .A2(G16), .A3(G23), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n789), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n792), .B(new_n793), .C1(G288), .C2(new_n734), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(KEYINPUT33), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n794), .A2(new_n796), .A3(G1976), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(G1976), .B1(new_n794), .B2(new_n796), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n785), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n734), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n734), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1971), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n780), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n785), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n794), .A2(new_n796), .ZN(new_n806));
  INV_X1    g381(.A(G1976), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n805), .B1(new_n808), .B2(new_n797), .ZN(new_n809));
  INV_X1    g384(.A(new_n803), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n809), .A2(new_n810), .A3(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n698), .A2(G25), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n486), .A2(G119), .B1(G131), .B2(new_n479), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(new_n698), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT35), .B(G1991), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT88), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G290), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G16), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G16), .B2(G24), .ZN(new_n825));
  INV_X1    g400(.A(G1986), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n822), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n779), .B1(new_n812), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g406(.A(KEYINPUT36), .B(new_n829), .C1(new_n804), .C2(new_n811), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n774), .B(new_n778), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n713), .A2(G2084), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n635), .A2(G29), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(G311));
  OR2_X1    g412(.A1(new_n759), .A2(new_n773), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n812), .A2(new_n830), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n812), .A2(new_n779), .A3(new_n830), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n834), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n835), .A4(new_n778), .ZN(G150));
  NAND2_X1  g419(.A1(new_n523), .A2(G55), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT97), .B(G93), .Z(new_n847));
  OAI221_X1 g422(.A(new_n845), .B1(new_n502), .B2(new_n846), .C1(new_n531), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n617), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n561), .A2(new_n848), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n561), .A2(new_n848), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT39), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n852), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n850), .B1(new_n857), .B2(G860), .ZN(G145));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n707), .B(G164), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n695), .A2(KEYINPUT100), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n754), .B(KEYINPUT99), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n486), .A2(G130), .B1(G142), .B2(new_n479), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n465), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n638), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n817), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n863), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n862), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n870), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G160), .B(KEYINPUT98), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n635), .Z(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n873), .B(new_n880), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n859), .B(new_n879), .C1(new_n881), .C2(new_n878), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g458(.A(new_n823), .B1(new_n786), .B2(new_n787), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n586), .A2(new_n587), .A3(new_n592), .A4(G290), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT102), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(G303), .A2(G305), .ZN(new_n888));
  NOR2_X1   g463(.A1(G166), .A2(new_n781), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(G303), .A2(G305), .ZN(new_n891));
  NAND2_X1  g466(.A1(G166), .A2(new_n781), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT102), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n886), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n890), .B2(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n621), .A2(new_n612), .ZN(new_n899));
  NAND4_X1  g474(.A1(G299), .A2(new_n610), .A3(new_n611), .A4(new_n606), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT41), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n628), .A2(new_n854), .A3(new_n853), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n855), .B1(new_n616), .B2(G559), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n900), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n890), .A2(new_n894), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n898), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n909), .B1(new_n898), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n848), .A2(new_n626), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(G295));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n917), .ZN(G331));
  NOR2_X1   g496(.A1(new_n896), .A2(new_n897), .ZN(new_n922));
  NAND2_X1  g497(.A1(G168), .A2(G301), .ZN(new_n923));
  NAND2_X1  g498(.A1(G171), .A2(G286), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n855), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n853), .A2(new_n923), .A3(new_n854), .A4(new_n924), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n908), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n901), .B2(new_n902), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n922), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n910), .A2(KEYINPUT103), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n933), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n859), .B1(new_n938), .B2(new_n933), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n931), .A2(new_n928), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n896), .B2(new_n897), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n938), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n940), .B(new_n941), .C1(new_n948), .C2(KEYINPUT43), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT43), .B1(new_n935), .B2(new_n939), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n948), .B2(KEYINPUT43), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n951), .B2(new_n941), .ZN(G397));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G164), .B2(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(G160), .A2(G40), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n820), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n817), .B(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G2067), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n707), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n754), .B(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n959), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n826), .B2(new_n823), .ZN(new_n967));
  NOR2_X1   g542(.A1(G290), .A2(G1986), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT107), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n956), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g545(.A1(G288), .A2(KEYINPUT112), .A3(new_n807), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n498), .A2(new_n500), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n492), .A2(new_n495), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n955), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT112), .B1(G288), .B2(new_n807), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n971), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(G305), .B(G1981), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT113), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT49), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n979), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n981), .B(new_n982), .C1(G1976), .C2(new_n788), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n955), .B1(KEYINPUT50), .B2(new_n976), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n974), .A2(new_n992), .A3(new_n975), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT109), .B(G2090), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n994), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n991), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n974), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n999));
  INV_X1    g574(.A(G40), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n470), .A2(new_n473), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n954), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1971), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n978), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1006), .B(new_n1009), .C1(G166), .C2(new_n978), .ZN(new_n1010));
  NAND4_X1  g585(.A1(G303), .A2(new_n1007), .A3(new_n1008), .A4(G8), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1005), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT115), .Z(new_n1013));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n991), .A2(new_n993), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  INV_X1    g591(.A(G2078), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n954), .A2(new_n999), .A3(new_n1017), .A4(new_n1001), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1015), .A2(new_n764), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1018), .A2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G171), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT126), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1016), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1025));
  AOI21_X1  g600(.A(G301), .B1(new_n1025), .B2(new_n1019), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1014), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1021), .A2(G171), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1019), .A3(G301), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(KEYINPUT54), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT124), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(G286), .B2(G8), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(G286), .A2(new_n1031), .A3(G8), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(G8), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1966), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1002), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT116), .B(G2084), .Z(new_n1040));
  NAND4_X1  g615(.A1(new_n1039), .A2(new_n1001), .A3(new_n993), .A4(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT123), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1034), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n1032), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1037), .A2(new_n1041), .A3(new_n1038), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT125), .B(KEYINPUT51), .Z(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(G8), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1048), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1027), .A2(new_n1030), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n577), .A2(G651), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n544), .A2(G91), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n523), .A2(new_n571), .A3(G53), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n571), .B1(new_n523), .B2(G53), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT119), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n570), .A2(new_n1064), .A3(new_n572), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1060), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT57), .B(G299), .C1(new_n1066), .C2(KEYINPUT118), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT56), .B(G2072), .Z(new_n1068));
  NOR2_X1   g643(.A1(new_n1002), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n991), .A2(new_n995), .A3(new_n997), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT117), .B(G1956), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1067), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1072), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1057), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1996), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n954), .A2(new_n999), .A3(new_n1079), .A4(new_n1001), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(KEYINPUT121), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(KEYINPUT121), .ZN(new_n1082));
  INV_X1    g657(.A(new_n977), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT58), .B(G1341), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n561), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT59), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1089), .A3(new_n561), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n614), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT60), .B1(new_n614), .B2(new_n615), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1039), .A2(new_n1001), .A3(new_n993), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1093), .A2(G1348), .B1(new_n1083), .B2(G2067), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1015), .A2(new_n1096), .B1(new_n961), .B2(new_n977), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n617), .A2(KEYINPUT60), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1088), .A2(new_n1090), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1067), .A2(new_n1100), .A3(new_n1075), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1101), .A2(new_n1102), .A3(new_n1072), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1067), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT61), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1078), .B(new_n1099), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1076), .A2(new_n616), .A3(new_n1097), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1056), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1052), .A2(KEYINPUT62), .A3(new_n1055), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1026), .A3(new_n1113), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n1053), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1013), .B1(new_n1109), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1093), .A2(new_n996), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1004), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT110), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n990), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1053), .A2(G286), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n988), .A2(new_n1125), .A3(new_n1126), .A4(new_n989), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT63), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n987), .A2(new_n807), .A3(new_n788), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(G1981), .B2(G305), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n979), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n970), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n956), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n962), .B2(new_n754), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT46), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(KEYINPUT127), .B2(new_n1136), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1134), .A2(G1996), .B1(KEYINPUT127), .B2(new_n1136), .ZN(new_n1138));
  OR4_X1    g713(.A1(KEYINPUT127), .A2(new_n1134), .A3(new_n1136), .A4(G1996), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT47), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n962), .A2(new_n963), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n818), .A2(new_n957), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1142), .A2(new_n1143), .B1(G2067), .B2(new_n707), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n956), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n969), .A2(new_n956), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT48), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n966), .B2(new_n1134), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1141), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1133), .A2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g725(.A(new_n940), .B(G319), .C1(new_n948), .C2(KEYINPUT43), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n882), .A2(new_n655), .A3(new_n689), .ZN(new_n1153));
  NOR3_X1   g727(.A1(new_n1152), .A2(G227), .A3(new_n1153), .ZN(G308));
  AND3_X1   g728(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n939), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n945), .A2(new_n947), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1156), .A2(new_n935), .ZN(new_n1157));
  INV_X1    g731(.A(KEYINPUT43), .ZN(new_n1158));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g733(.A1(new_n882), .A2(new_n655), .A3(new_n689), .ZN(new_n1160));
  INV_X1    g734(.A(G227), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(G319), .A4(new_n1161), .ZN(G225));
endmodule


