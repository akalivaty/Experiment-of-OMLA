//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT7), .ZN(new_n203));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  INV_X1    g004(.A(G92gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(KEYINPUT8), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G99gat), .B(G106gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT93), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(KEYINPUT15), .A3(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n216), .B(KEYINPUT85), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n215), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT17), .ZN(new_n225));
  NAND2_X1  g024(.A1(G232gat), .A2(G233gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n212), .A2(new_n225), .B1(KEYINPUT41), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n210), .B(KEYINPUT93), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G190gat), .B(G218gat), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n232), .B(KEYINPUT94), .Z(new_n233));
  NOR2_X1   g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n227), .A2(KEYINPUT41), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT92), .ZN(new_n237));
  XOR2_X1   g036(.A(G134gat), .B(G162gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n239), .A2(KEYINPUT95), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n233), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n235), .A2(new_n241), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n239), .B(KEYINPUT95), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G57gat), .B(G64gat), .Z(new_n247));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G71gat), .B(G78gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT9), .ZN(new_n252));
  INV_X1    g051(.A(G71gat), .ZN(new_n253));
  INV_X1    g052(.A(G78gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n255), .A3(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n255), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(new_n249), .A3(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(KEYINPUT21), .ZN(new_n260));
  XOR2_X1   g059(.A(G127gat), .B(G155gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G15gat), .B(G22gat), .ZN(new_n263));
  INV_X1    g062(.A(G1gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT16), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n265), .B(new_n266), .C1(new_n264), .C2(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(KEYINPUT21), .B2(new_n259), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n262), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G231gat), .A2(G233gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT91), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G183gat), .B(G211gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n271), .B(new_n277), .Z(new_n278));
  NOR2_X1   g077(.A1(new_n246), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G230gat), .ZN(new_n280));
  INV_X1    g079(.A(G233gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n259), .A2(KEYINPUT10), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n212), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n210), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n259), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n210), .A2(new_n256), .A3(new_n258), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT10), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n282), .A3(new_n288), .ZN(new_n291));
  XNOR2_X1  g090(.A(G120gat), .B(G148gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G176gat), .B(G204gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  AND3_X1   g093(.A1(new_n290), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n290), .B2(new_n291), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n301));
  INV_X1    g100(.A(G211gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT22), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT70), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT22), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n299), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n316));
  OAI21_X1  g115(.A(G218gat), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(new_n312), .A3(new_n299), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  AND2_X1   g121(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n324));
  OAI21_X1  g123(.A(G155gat), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT2), .ZN(new_n326));
  XNOR2_X1  g125(.A(G141gat), .B(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G162gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n331), .A2(G162gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n329), .A2(G155gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT75), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n326), .A2(new_n328), .A3(new_n334), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339));
  OAI22_X1  g138(.A1(new_n327), .A2(KEYINPUT2), .B1(new_n335), .B2(new_n336), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n321), .B1(new_n322), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n337), .A2(new_n328), .A3(new_n334), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n325), .A2(KEYINPUT2), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n314), .B2(new_n320), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n345), .B1(new_n344), .B2(new_n350), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n312), .B1(new_n319), .B2(new_n299), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n314), .A2(KEYINPUT79), .A3(new_n320), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n356), .B2(new_n357), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT3), .ZN(new_n361));
  INV_X1    g160(.A(new_n348), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT81), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n357), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT80), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n339), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n368), .A3(new_n348), .ZN(new_n369));
  INV_X1    g168(.A(new_n342), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(G22gat), .B(new_n353), .C1(new_n371), .C2(new_n343), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT3), .B1(new_n364), .B2(KEYINPUT80), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n362), .B1(new_n374), .B2(new_n366), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n370), .B1(new_n375), .B2(new_n368), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n361), .A2(KEYINPUT81), .A3(new_n362), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n343), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n353), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n373), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381));
  INV_X1    g180(.A(G50gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n372), .A2(new_n380), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n343), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n348), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n342), .B1(new_n389), .B2(KEYINPUT81), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n390), .B2(new_n369), .ZN(new_n391));
  OAI21_X1  g190(.A(G22gat), .B1(new_n391), .B2(new_n353), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n378), .A2(new_n373), .A3(new_n379), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n385), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT35), .ZN(new_n396));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G183gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT27), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G183gat), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT64), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT28), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n400), .A2(new_n402), .A3(new_n405), .A4(new_n403), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n417));
  INV_X1    g216(.A(G169gat), .ZN(new_n418));
  INV_X1    g217(.A(G176gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT65), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n415), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT66), .B1(new_n413), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G113gat), .B(G120gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n429), .B1(new_n430), .B2(KEYINPUT1), .ZN(new_n431));
  INV_X1    g230(.A(new_n430), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT24), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n436), .A2(new_n437), .B1(G169gat), .B2(G176gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT23), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n418), .A3(new_n419), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n399), .A2(new_n403), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(KEYINPUT24), .A3(new_n411), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n438), .A2(new_n442), .A3(new_n444), .A4(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n412), .A2(new_n411), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n410), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n427), .A2(new_n435), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n434), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n449), .A2(new_n453), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n451), .B1(new_n459), .B2(new_n452), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n454), .A2(new_n455), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n398), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT68), .ZN(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n454), .A2(new_n455), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n473), .A2(new_n397), .A3(new_n461), .A4(new_n456), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT69), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n466), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n477), .B2(new_n471), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT32), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n472), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n480), .B2(new_n472), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n321), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT72), .B1(new_n458), .B2(new_n460), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n427), .A2(new_n486), .A3(new_n449), .A4(new_n453), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n322), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G226gat), .A2(G233gat), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n488), .A2(KEYINPUT73), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n449), .B1(new_n426), .B2(new_n413), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(G226gat), .A3(G233gat), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n488), .A2(new_n489), .B1(KEYINPUT73), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n484), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n322), .A3(new_n489), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n485), .A2(new_n487), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(new_n489), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n321), .ZN(new_n498));
  XOR2_X1   g297(.A(G8gat), .B(G36gat), .Z(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT74), .ZN(new_n500));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  NAND3_X1  g301(.A1(new_n494), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(new_n341), .A3(new_n457), .ZN(new_n507));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n348), .B2(new_n457), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n435), .A2(new_n338), .A3(KEYINPUT4), .A4(new_n340), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n507), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n508), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n348), .A2(new_n457), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n338), .A2(new_n340), .B1(new_n434), .B2(new_n431), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n510), .A2(new_n511), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT5), .A3(new_n508), .A4(new_n507), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G1gat), .B(G29gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT0), .ZN(new_n523));
  XNOR2_X1  g322(.A(G57gat), .B(G85gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n518), .A2(new_n525), .A3(new_n520), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n518), .A2(new_n520), .A3(KEYINPUT6), .A4(new_n525), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n498), .A4(new_n502), .ZN(new_n535));
  INV_X1    g334(.A(new_n502), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n488), .A2(new_n489), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n492), .A2(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n488), .A2(KEYINPUT73), .A3(new_n489), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n321), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n497), .A2(new_n321), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n505), .A2(new_n534), .A3(new_n535), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n395), .A2(new_n396), .A3(new_n483), .A4(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n386), .B1(new_n372), .B2(new_n380), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n392), .A2(new_n393), .A3(new_n385), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n483), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT35), .B1(new_n549), .B2(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n494), .A2(new_n498), .A3(new_n502), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n534), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n321), .B1(new_n490), .B2(new_n493), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n497), .B2(new_n484), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT38), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n502), .B1(new_n494), .B2(new_n498), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n502), .A2(new_n555), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n494), .B2(new_n498), .ZN(new_n561));
  INV_X1    g360(.A(new_n559), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n543), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT38), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n553), .B(new_n560), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n505), .A2(new_n535), .A3(new_n543), .ZN(new_n566));
  INV_X1    g365(.A(new_n529), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n519), .A2(new_n507), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n513), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n514), .A2(new_n515), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n569), .B(KEYINPUT39), .C1(new_n513), .C2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n571), .B(new_n526), .C1(new_n569), .C2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n567), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n566), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n395), .A2(new_n565), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n547), .A2(new_n548), .ZN(new_n580));
  INV_X1    g379(.A(new_n482), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n472), .A2(new_n476), .A3(new_n480), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT36), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n481), .B2(new_n482), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n580), .A2(new_n544), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n579), .B1(new_n586), .B2(KEYINPUT83), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n544), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n585), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n588), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n551), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n269), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n225), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n269), .A2(new_n224), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT87), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G197gat), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT11), .B(G169gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n594), .B(KEYINPUT13), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n269), .A2(new_n224), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n595), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n596), .B2(new_n597), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n593), .A2(KEYINPUT18), .A3(new_n594), .A4(new_n595), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n610), .B(new_n609), .C1(new_n598), .C2(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT88), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(KEYINPUT88), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n591), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT89), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n591), .A2(KEYINPUT89), .A3(new_n618), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n298), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n534), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G1gat), .ZN(G1324gat));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  INV_X1    g426(.A(new_n298), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n591), .A2(KEYINPUT89), .A3(new_n618), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT89), .B1(new_n591), .B2(new_n618), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n566), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n627), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g434(.A(KEYINPUT96), .B(new_n627), .C1(new_n631), .C2(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n632), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n623), .A2(KEYINPUT42), .A3(new_n566), .A4(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n631), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n642), .A2(KEYINPUT97), .A3(KEYINPUT42), .A4(new_n638), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n631), .A2(G8gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n644), .A3(new_n645), .ZN(G1325gat));
  INV_X1    g445(.A(new_n623), .ZN(new_n647));
  OAI21_X1  g446(.A(G15gat), .B1(new_n647), .B2(new_n589), .ZN(new_n648));
  INV_X1    g447(.A(new_n483), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(G15gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n647), .B2(new_n650), .ZN(G1326gat));
  OAI211_X1 g450(.A(new_n580), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n653), .B2(new_n654), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(G1327gat));
  NAND2_X1  g457(.A1(new_n621), .A2(new_n622), .ZN(new_n659));
  INV_X1    g458(.A(new_n278), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n295), .A2(new_n296), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n245), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n666));
  INV_X1    g465(.A(G29gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n624), .A2(new_n667), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n579), .A2(new_n586), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n245), .B1(new_n551), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT44), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n591), .A2(KEYINPUT44), .A3(new_n246), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n614), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n663), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G29gat), .B1(new_n677), .B2(new_n534), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n666), .B1(new_n665), .B2(new_n668), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n669), .A2(new_n678), .A3(new_n679), .ZN(G1328gat));
  INV_X1    g479(.A(new_n566), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(G36gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n659), .A2(new_n664), .A3(new_n682), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n683), .A2(KEYINPUT99), .A3(KEYINPUT46), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT99), .B1(new_n683), .B2(KEYINPUT46), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n677), .B2(new_n681), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .A4(new_n687), .ZN(G1329gat));
  INV_X1    g487(.A(new_n589), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n673), .A3(new_n689), .A4(new_n676), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G43gat), .ZN(new_n691));
  OR2_X1    g490(.A1(KEYINPUT100), .A2(KEYINPUT47), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n649), .A2(G43gat), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n691), .B(new_n692), .C1(new_n665), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(KEYINPUT100), .A2(KEYINPUT47), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1330gat));
  NAND4_X1  g495(.A1(new_n672), .A2(new_n673), .A3(new_n580), .A4(new_n676), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G50gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n580), .A2(new_n382), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n665), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1331gat));
  NAND3_X1  g501(.A1(new_n279), .A2(new_n675), .A3(new_n661), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT101), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n551), .A2(new_n670), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n624), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT102), .B(G57gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n681), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT104), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  NAND3_X1  g516(.A1(new_n706), .A2(new_n253), .A3(new_n483), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n704), .A2(new_n705), .A3(new_n589), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n253), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n580), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT105), .B(G78gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1335gat));
  NOR3_X1   g523(.A1(new_n660), .A2(new_n614), .A3(new_n297), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n674), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n534), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n660), .A2(new_n614), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n671), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT51), .Z(new_n730));
  NAND4_X1  g529(.A1(new_n730), .A2(new_n205), .A3(new_n624), .A4(new_n661), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(G1336gat));
  NOR3_X1   g531(.A1(new_n681), .A2(G92gat), .A3(new_n297), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT52), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n674), .A2(new_n566), .A3(new_n725), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G92gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(KEYINPUT51), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n729), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n729), .A2(new_n739), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n735), .A2(G92gat), .B1(new_n742), .B2(new_n733), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n737), .B1(new_n743), .B2(new_n744), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n726), .B2(new_n589), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n649), .A2(G99gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n661), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1338gat));
  NOR3_X1   g548(.A1(new_n395), .A2(G106gat), .A3(new_n297), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n740), .B2(new_n741), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT107), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n672), .A2(new_n673), .A3(new_n580), .A4(new_n725), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n755), .B(new_n750), .C1(new_n740), .C2(new_n741), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT53), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT53), .B1(new_n730), .B2(new_n750), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n754), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1339gat));
  NOR4_X1   g560(.A1(new_n246), .A2(new_n278), .A3(new_n614), .A4(new_n661), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n607), .A2(new_n595), .A3(new_n606), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n602), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n609), .A2(new_n603), .A3(new_n610), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n661), .A2(KEYINPUT109), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n765), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n297), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n259), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n287), .A2(new_n288), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT10), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n775), .A3(new_n282), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n290), .A2(new_n776), .A3(KEYINPUT54), .ZN(new_n777));
  INV_X1    g576(.A(new_n294), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n290), .B2(KEYINPUT54), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n771), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n295), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n282), .B1(new_n772), .B2(new_n775), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n294), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n290), .A2(new_n776), .A3(KEYINPUT54), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n780), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n767), .B(new_n770), .C1(new_n675), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n245), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n245), .A2(new_n787), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n769), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n762), .B1(new_n794), .B2(new_n278), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n549), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n566), .A2(new_n534), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n618), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n675), .A2(G113gat), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT110), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n799), .B2(new_n803), .ZN(G1340gat));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n661), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT111), .B(G120gat), .Z(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1341gat));
  NAND2_X1  g606(.A1(new_n798), .A2(new_n660), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G127gat), .ZN(G1342gat));
  INV_X1    g608(.A(G134gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n798), .B2(new_n246), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n246), .A2(new_n681), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT112), .Z(new_n813));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n810), .A3(new_n624), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT113), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n811), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n816), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n814), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(KEYINPUT56), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n817), .B1(new_n818), .B2(new_n822), .ZN(G1343gat));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n589), .A2(new_n797), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n787), .B1(new_n616), .B2(new_n617), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n769), .A2(new_n297), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n245), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n660), .B1(new_n828), .B2(new_n793), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT57), .B(new_n580), .C1(new_n829), .C2(new_n762), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n279), .A2(new_n675), .A3(new_n297), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n788), .A2(new_n245), .B1(new_n790), .B2(new_n792), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n660), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT57), .B1(new_n833), .B2(new_n580), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT115), .B(KEYINPUT57), .C1(new_n833), .C2(new_n580), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n825), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n824), .B(G141gat), .C1(new_n838), .C2(new_n800), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n589), .A2(new_n580), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n833), .A2(new_n624), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n566), .ZN(new_n844));
  INV_X1    g643(.A(G141gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n618), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n839), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n614), .B(new_n825), .C1(new_n836), .C2(new_n837), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(G141gat), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n824), .B2(new_n851), .ZN(G1344gat));
  OAI211_X1 g651(.A(new_n661), .B(new_n825), .C1(new_n836), .C2(new_n837), .ZN(new_n853));
  INV_X1    g652(.A(G148gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(KEYINPUT59), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n795), .B2(new_n395), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n395), .A2(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n298), .A2(new_n618), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n829), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n825), .A2(new_n661), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G148gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT59), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n854), .A3(new_n661), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(KEYINPUT118), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n853), .A2(new_n855), .B1(KEYINPUT59), .B2(new_n863), .ZN(new_n869));
  INV_X1    g668(.A(new_n866), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n871), .ZN(G1345gat));
  OAI21_X1  g671(.A(G155gat), .B1(new_n838), .B2(new_n278), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n844), .A2(new_n331), .A3(new_n660), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  OR2_X1    g674(.A1(new_n323), .A2(new_n324), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n838), .B2(new_n245), .ZN(new_n877));
  INV_X1    g676(.A(new_n813), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n843), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT119), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n877), .A2(new_n882), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n681), .A2(new_n624), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n795), .A2(new_n549), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n418), .B1(new_n887), .B2(new_n618), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT120), .Z(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n418), .A3(new_n614), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1348gat));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n661), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(G176gat), .ZN(G1349gat));
  INV_X1    g692(.A(new_n549), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n833), .A2(new_n894), .A3(new_n660), .A4(new_n885), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n399), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n400), .A2(new_n402), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(KEYINPUT121), .B2(new_n399), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n897), .B(KEYINPUT122), .C1(new_n895), .C2(new_n899), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT60), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT123), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT123), .A4(KEYINPUT60), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1350gat));
  NOR2_X1   g708(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n887), .B2(new_n246), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n911), .B(new_n912), .Z(G1351gat));
  NAND3_X1  g712(.A1(new_n589), .A2(new_n580), .A3(new_n566), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n833), .B(new_n534), .C1(KEYINPUT124), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(KEYINPUT124), .B2(new_n914), .ZN(new_n916));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n614), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n886), .A2(new_n689), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n857), .A2(new_n860), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n618), .A2(G197gat), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1352gat));
  XNOR2_X1  g720(.A(KEYINPUT125), .B(G204gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n916), .A2(new_n661), .A3(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n919), .A2(new_n661), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n924), .B(new_n925), .C1(new_n926), .C2(new_n922), .ZN(G1353gat));
  NAND4_X1  g726(.A1(new_n916), .A2(new_n303), .A3(new_n304), .A4(new_n660), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n857), .A2(new_n860), .A3(new_n660), .A4(new_n918), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT126), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n300), .A3(new_n246), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n919), .A2(new_n246), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n300), .ZN(G1355gat));
endmodule


