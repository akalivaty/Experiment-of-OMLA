//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G77), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G87), .A2(G250), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G226), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(KEYINPUT9), .ZN(new_n244));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n214), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n206), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT69), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n206), .A2(KEYINPUT69), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT8), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT68), .ZN(new_n254));
  INV_X1    g0054(.A(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT8), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT67), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n251), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n259), .A2(new_n261), .B1(new_n201), .B2(new_n206), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n246), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT70), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G50), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n246), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n205), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n268), .B1(new_n271), .B2(new_n267), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n263), .B2(KEYINPUT70), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n244), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n264), .A2(new_n244), .A3(new_n273), .ZN(new_n276));
  OR2_X1    g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G222), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n279), .B(new_n281), .C1(new_n282), .C2(new_n280), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n283), .B(new_n286), .C1(G77), .C2(new_n279), .ZN(new_n287));
  AND2_X1   g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT66), .B1(new_n288), .B2(new_n214), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT66), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n284), .A2(new_n290), .A3(G1), .A4(G13), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G226), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n289), .A2(G274), .A3(new_n291), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n287), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n275), .A2(new_n276), .B1(G190), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(G200), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n301), .B(new_n302), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(G190), .ZN(new_n304));
  INV_X1    g0104(.A(new_n276), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n302), .B(new_n304), .C1(new_n305), .C2(new_n274), .ZN(new_n306));
  OAI211_X1 g0106(.A(KEYINPUT72), .B(new_n304), .C1(new_n305), .C2(new_n274), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n299), .A2(G179), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n299), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n264), .A2(new_n273), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n303), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n269), .A2(G68), .A3(new_n270), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT12), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n265), .B2(G68), .ZN(new_n318));
  INV_X1    g0118(.A(G68), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n266), .A2(KEYINPUT12), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n249), .A2(G77), .A3(new_n250), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n319), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n269), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n321), .B1(new_n324), .B2(KEYINPUT11), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n324), .A2(KEYINPUT11), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n280), .A2(G226), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G232), .A2(G1698), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n277), .A2(new_n278), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n286), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n289), .A2(G238), .A3(new_n291), .A4(new_n293), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n298), .A4(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n336), .A2(G190), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n328), .A2(new_n329), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n279), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n335), .B(new_n298), .C1(new_n339), .C2(new_n285), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n327), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(KEYINPUT73), .A3(new_n336), .ZN(new_n343));
  OR3_X1    g0143(.A1(new_n340), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(G200), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n344), .A3(G169), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT14), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n343), .A2(new_n344), .A3(new_n349), .A4(G169), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n341), .A2(G179), .A3(new_n336), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n325), .A2(new_n326), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n346), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G238), .A2(G1698), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n279), .B(new_n358), .C1(new_n230), .C2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n286), .C1(G107), .C2(new_n279), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n292), .A2(new_n217), .A3(new_n293), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n298), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n311), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n364), .A2(new_n247), .B1(new_n206), .B2(new_n202), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n261), .B1(new_n253), .B2(new_n256), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n246), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n266), .A2(new_n202), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(new_n202), .C2(new_n271), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n362), .A2(G179), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n363), .A2(KEYINPUT71), .A3(new_n369), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n369), .B1(new_n362), .B2(G200), .ZN(new_n376));
  INV_X1    g0176(.A(G190), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n362), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  XNOR2_X1  g0182(.A(G58), .B(G68), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(G20), .ZN(new_n384));
  AND2_X1   g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n382), .B(G20), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n384), .A2(new_n388), .B1(new_n389), .B2(new_n261), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n277), .A2(new_n206), .A3(new_n278), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  NOR2_X1   g0194(.A1(KEYINPUT3), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n319), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n381), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n396), .B2(new_n206), .ZN(new_n400));
  NOR4_X1   g0200(.A1(new_n394), .A2(new_n395), .A3(new_n392), .A4(G20), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n385), .B2(new_n386), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT75), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(new_n387), .B1(G159), .B2(new_n260), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT16), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(new_n246), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n254), .A2(new_n257), .ZN(new_n408));
  INV_X1    g0208(.A(new_n271), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n408), .B2(new_n265), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n205), .B(G274), .C1(G41), .C2(G45), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n297), .B2(new_n230), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n415), .A2(new_n289), .A3(new_n291), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n282), .A2(new_n280), .ZN(new_n417));
  INV_X1    g0217(.A(G226), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n419), .C1(new_n394), .C2(new_n395), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n285), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n413), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n286), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n289), .A3(new_n291), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n377), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n407), .A2(new_n412), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT17), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  INV_X1    g0231(.A(G179), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n416), .A2(new_n432), .A3(new_n422), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n311), .B1(new_n425), .B2(new_n426), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(G169), .B1(new_n416), .B2(new_n422), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n425), .A2(G179), .A3(new_n426), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT76), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n402), .A2(new_n405), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n269), .B1(new_n441), .B2(new_n381), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n411), .B1(new_n442), .B2(new_n406), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n431), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n435), .B1(new_n433), .B2(new_n434), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n437), .A2(KEYINPUT76), .A3(new_n438), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n407), .A2(new_n412), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT18), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n357), .A2(new_n380), .A3(new_n430), .A4(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n315), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n205), .A2(G33), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n265), .A2(new_n454), .A3(new_n214), .A4(new_n245), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT80), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n455), .A2(new_n456), .B1(new_n265), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(new_n459), .A3(G20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n246), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT84), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT84), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n466), .A3(new_n246), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n206), .C1(G33), .C2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n463), .A2(new_n466), .A3(new_n246), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n466), .B1(new_n463), .B2(new_n246), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT20), .B(new_n471), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n462), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT5), .B(G41), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n289), .A2(new_n478), .A3(new_n480), .A4(new_n291), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n296), .A2(G1), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n292), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n485), .B2(G270), .ZN(new_n486));
  OAI211_X1 g0286(.A(G257), .B(new_n280), .C1(new_n394), .C2(new_n395), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n277), .A2(G303), .A3(new_n278), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(G264), .A2(G1698), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n394), .B2(new_n395), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT82), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(KEYINPUT82), .B(new_n490), .C1(new_n394), .C2(new_n395), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n286), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n494), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n487), .A2(new_n488), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n486), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n477), .A2(new_n502), .A3(KEYINPUT21), .A4(G169), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n292), .A2(new_n484), .ZN(new_n504));
  INV_X1    g0304(.A(G270), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n481), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n499), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n285), .B1(new_n507), .B2(KEYINPUT83), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(new_n500), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n477), .A2(new_n509), .A3(G179), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g0311(.A(KEYINPUT85), .B(KEYINPUT21), .Z(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(KEYINPUT83), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n286), .A3(new_n500), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n311), .B1(new_n514), .B2(new_n486), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n512), .B1(new_n515), .B2(new_n477), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n477), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(G190), .A3(new_n486), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n413), .C2(new_n509), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n484), .A2(G257), .A3(new_n289), .A4(new_n291), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n481), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT79), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(KEYINPUT79), .A3(new_n481), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(G1698), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n527), .B(G244), .C1(new_n395), .C2(new_n394), .ZN(new_n528));
  INV_X1    g0328(.A(G244), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n277), .B2(new_n278), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(new_n469), .C1(new_n530), .C2(KEYINPUT4), .ZN(new_n531));
  OAI21_X1  g0331(.A(G250), .B1(new_n394), .B2(new_n395), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n280), .B1(new_n532), .B2(KEYINPUT4), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n286), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n524), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(KEYINPUT6), .B2(G97), .ZN(new_n538));
  XNOR2_X1  g0338(.A(KEYINPUT77), .B(G107), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  OAI21_X1  g0341(.A(G20), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n260), .A2(G77), .ZN(new_n543));
  OAI21_X1  g0343(.A(G107), .B1(new_n400), .B2(new_n401), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n246), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n269), .A2(KEYINPUT78), .A3(new_n265), .A4(new_n454), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n455), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n549), .A3(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n266), .A2(new_n470), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n521), .A2(new_n481), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n534), .A3(G190), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n546), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n534), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n546), .A2(new_n553), .B1(new_n557), .B2(new_n311), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n524), .A2(new_n432), .A3(new_n525), .A4(new_n534), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n536), .A2(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n364), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n547), .A2(new_n549), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G87), .ZN(new_n563));
  INV_X1    g0363(.A(G107), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n470), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n331), .A2(new_n206), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT19), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n206), .B(G68), .C1(new_n394), .C2(new_n395), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n247), .B2(new_n470), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n246), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n364), .A2(new_n266), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n562), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n460), .A2(G33), .ZN(new_n575));
  OR2_X1    g0375(.A1(G238), .A2(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n529), .A2(G1698), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n394), .C2(new_n395), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n285), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G250), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n479), .B1(new_n483), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n581), .A2(new_n289), .A3(new_n291), .ZN(new_n582));
  OAI21_X1  g0382(.A(G169), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n289), .A3(new_n291), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n576), .A2(new_n577), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(new_n279), .B1(new_n460), .B2(G33), .ZN(new_n586));
  OAI211_X1 g0386(.A(G179), .B(new_n584), .C1(new_n586), .C2(new_n285), .ZN(new_n587));
  AOI22_X1  g0387(.A1(KEYINPUT81), .A2(new_n574), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n574), .A2(KEYINPUT81), .ZN(new_n589));
  OAI21_X1  g0389(.A(G200), .B1(new_n579), .B2(new_n582), .ZN(new_n590));
  OAI211_X1 g0390(.A(G190), .B(new_n584), .C1(new_n586), .C2(new_n285), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n547), .A2(new_n549), .A3(G87), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n593), .A2(new_n572), .A3(new_n573), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n588), .A2(new_n589), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G257), .B(G1698), .C1(new_n394), .C2(new_n395), .ZN(new_n596));
  OAI211_X1 g0396(.A(G250), .B(new_n280), .C1(new_n394), .C2(new_n395), .ZN(new_n597));
  NAND2_X1  g0397(.A1(G33), .A2(G294), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n286), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n484), .A2(G264), .A3(new_n289), .A4(new_n291), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n481), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n602), .A2(G179), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n311), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n206), .B(G87), .C1(new_n394), .C2(new_n395), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT22), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT22), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n279), .A2(new_n607), .A3(new_n206), .A4(G87), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n247), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT23), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n206), .A2(G107), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n460), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT86), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n612), .B2(new_n611), .ZN(new_n615));
  OAI211_X1 g0415(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n206), .C2(G107), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT24), .B1(new_n609), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n613), .A2(new_n617), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT24), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n606), .A2(new_n608), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n269), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n547), .A2(new_n549), .A3(G107), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n265), .A2(G107), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT25), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n603), .B(new_n604), .C1(new_n624), .C2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n609), .A2(new_n618), .A3(KEYINPUT24), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n246), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n602), .A2(new_n413), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n600), .A2(new_n377), .A3(new_n481), .A4(new_n601), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n628), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n595), .A2(new_n629), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n517), .A2(new_n520), .A3(new_n560), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n453), .A2(new_n639), .ZN(G372));
  NOR2_X1   g0440(.A1(new_n433), .A2(new_n434), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n443), .A2(KEYINPUT18), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n641), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n431), .B1(new_n448), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n374), .A2(new_n373), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT71), .B1(new_n363), .B2(new_n369), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n342), .A2(new_n345), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n356), .A2(new_n352), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(KEYINPUT89), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n430), .B1(new_n650), .B2(KEYINPUT89), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n645), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n303), .A2(new_n309), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n313), .B2(new_n312), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n546), .A2(new_n553), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n557), .A2(new_n311), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n656), .A2(new_n559), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n595), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n656), .A2(new_n559), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n592), .A2(new_n594), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n583), .A2(new_n587), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n574), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n659), .B(KEYINPUT88), .C1(KEYINPUT26), .C2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n658), .A2(new_n667), .A3(KEYINPUT26), .A4(new_n595), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n477), .A2(new_n502), .A3(G169), .ZN(new_n670));
  INV_X1    g0470(.A(new_n512), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n503), .A3(new_n510), .A4(new_n629), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT87), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n552), .B1(new_n545), .B2(new_n246), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n536), .A2(new_n675), .A3(new_n555), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(new_n660), .A3(new_n637), .A4(new_n661), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n673), .B2(KEYINPUT87), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n669), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n655), .B1(new_n453), .B2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n672), .A2(new_n503), .A3(new_n510), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n518), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n520), .A2(new_n672), .A3(new_n503), .A4(new_n510), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n687), .B1(new_n624), .B2(new_n628), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n629), .A2(new_n637), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n632), .A2(new_n636), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(new_n603), .A3(new_n604), .A4(new_n687), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT90), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n629), .A2(new_n687), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n688), .B1(new_n511), .B2(new_n516), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT91), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(new_n688), .C1(new_n511), .C2(new_n516), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n705), .B1(new_n710), .B2(new_n703), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n209), .ZN(new_n713));
  OR3_X1    g0513(.A1(new_n713), .A2(KEYINPUT92), .A3(G41), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT92), .B1(new_n713), .B2(G41), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n565), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n212), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT26), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n658), .A2(new_n721), .A3(new_n595), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT26), .B1(new_n660), .B2(new_n664), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n722), .A2(new_n723), .A3(new_n663), .ZN(new_n724));
  AND4_X1   g0524(.A1(new_n660), .A2(new_n676), .A3(new_n661), .A4(new_n637), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n673), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n687), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n674), .A2(new_n678), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n668), .A2(new_n663), .ZN(new_n730));
  INV_X1    g0530(.A(new_n665), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n667), .B1(new_n731), .B2(new_n721), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n730), .B1(new_n732), .B2(new_n659), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n687), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n728), .B1(new_n734), .B2(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(G330), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n560), .A2(new_n595), .A3(new_n629), .A4(new_n637), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT31), .B1(new_n737), .B2(new_n691), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n600), .A2(new_n601), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n557), .A2(new_n587), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n509), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n584), .B1(new_n586), .B2(new_n285), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n602), .A2(new_n432), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n502), .A2(new_n743), .A3(new_n535), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n509), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n747), .A2(KEYINPUT93), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n587), .ZN(new_n750));
  INV_X1    g0550(.A(new_n739), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(new_n554), .A4(new_n534), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n748), .B1(new_n752), .B2(new_n502), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n745), .A2(new_n746), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n687), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n738), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n745), .A2(new_n753), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n736), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n735), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n720), .B1(new_n763), .B2(G1), .ZN(G364));
  INV_X1    g0564(.A(new_n716), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n206), .A2(G13), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n205), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n214), .B1(G20), .B2(new_n311), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n377), .A2(G200), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n206), .B1(new_n773), .B2(new_n432), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT98), .Z(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G97), .ZN(new_n776));
  NAND2_X1  g0576(.A1(G20), .A2(G179), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n377), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n413), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(KEYINPUT97), .B1(new_n377), .B2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n377), .A2(KEYINPUT97), .A3(G20), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n413), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n776), .B1(new_n319), .B2(new_n781), .C1(new_n564), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n779), .A2(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n790), .A2(KEYINPUT96), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(KEYINPUT96), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n788), .B1(new_n794), .B2(G77), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n377), .A2(new_n413), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(G20), .A3(new_n432), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n396), .B1(new_n798), .B2(G87), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n778), .A2(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n778), .A2(new_n773), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n267), .C1(new_n255), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n785), .A2(G200), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G159), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n802), .B1(KEYINPUT32), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n795), .B(new_n805), .C1(KEYINPUT32), .C2(new_n804), .ZN(new_n806));
  INV_X1    g0606(.A(new_n800), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G326), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n774), .C1(new_n790), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT99), .ZN(new_n812));
  INV_X1    g0612(.A(G322), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n396), .B1(new_n801), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n797), .B(KEYINPUT100), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G303), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n780), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G283), .A2(new_n786), .B1(new_n803), .B2(G329), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n812), .A2(new_n816), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n772), .B1(new_n806), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G13), .A2(G33), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n771), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT94), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n242), .A2(G45), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n713), .A2(new_n279), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G45), .C2(new_n212), .ZN(new_n829));
  INV_X1    g0629(.A(G355), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n209), .A2(new_n279), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(G116), .B2(new_n209), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n770), .B(new_n821), .C1(new_n826), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT101), .Z(new_n834));
  INV_X1    g0634(.A(new_n824), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n692), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n694), .A2(new_n769), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(G330), .B2(new_n692), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  NAND2_X1  g0640(.A1(new_n369), .A2(new_n687), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n375), .A2(new_n378), .A3(new_n841), .ZN(new_n842));
  OR3_X1    g0642(.A1(new_n646), .A2(new_n647), .A3(new_n841), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n380), .A2(new_n688), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n734), .A2(new_n844), .B1(new_n679), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n769), .B1(new_n846), .B2(new_n762), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n762), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n771), .A2(new_n822), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n770), .B1(new_n202), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n279), .B1(new_n815), .B2(G107), .ZN(new_n851));
  INV_X1    g0651(.A(G303), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n809), .B2(new_n801), .C1(new_n852), .C2(new_n800), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n787), .A2(new_n563), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G283), .B2(new_n780), .ZN(new_n855));
  INV_X1    g0655(.A(new_n803), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n855), .B(new_n776), .C1(new_n810), .C2(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n853), .B(new_n857), .C1(new_n460), .C2(new_n794), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n807), .A2(G137), .ZN(new_n859));
  INV_X1    g0659(.A(G143), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n860), .B2(new_n801), .C1(new_n781), .C2(new_n259), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n794), .B2(G159), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT34), .Z(new_n863));
  OAI21_X1  g0663(.A(new_n279), .B1(new_n774), .B2(new_n255), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n815), .A2(G50), .B1(new_n786), .B2(G68), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT102), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(G132), .C2(new_n803), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n858), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n850), .B1(new_n823), .B2(new_n844), .C1(new_n868), .C2(new_n772), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n848), .A2(new_n869), .ZN(G384));
  NOR2_X1   g0670(.A1(new_n540), .A2(new_n541), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(KEYINPUT35), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(KEYINPUT35), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n873), .A2(G116), .A3(new_n215), .A4(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT36), .Z(new_n876));
  OAI211_X1 g0676(.A(new_n213), .B(G77), .C1(new_n255), .C2(new_n319), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n267), .A2(G68), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n205), .B(G13), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n352), .A2(new_n356), .A3(new_n688), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  INV_X1    g0683(.A(new_n685), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n448), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n450), .B2(new_n430), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n448), .A2(new_n643), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n885), .A3(new_n429), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT37), .B1(new_n443), .B2(new_n428), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n448), .B1(new_n447), .B2(new_n884), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n888), .A2(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n886), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n886), .B2(new_n891), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(KEYINPUT104), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT104), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n896), .B(new_n892), .C1(new_n886), .C2(new_n891), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n883), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n885), .B1(new_n645), .B2(new_n430), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n892), .B1(new_n899), .B2(new_n891), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT18), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT18), .B1(new_n447), .B2(new_n448), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT17), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n443), .B2(new_n428), .ZN(new_n904));
  AND4_X1   g0704(.A1(new_n903), .A2(new_n407), .A3(new_n412), .A4(new_n428), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n901), .A2(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n443), .A2(new_n685), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n429), .B1(new_n443), .B2(new_n641), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n909), .B2(new_n907), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n890), .A2(new_n889), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n900), .A2(new_n913), .A3(new_n883), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n900), .A2(new_n913), .A3(KEYINPUT105), .A4(new_n883), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n882), .B1(new_n898), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n648), .A2(new_n688), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n679), .B2(new_n845), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n906), .A2(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT104), .B1(new_n925), .B2(KEYINPUT38), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n897), .A3(new_n913), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n353), .A2(new_n355), .A3(new_n687), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n928), .B(new_n346), .C1(new_n352), .C2(new_n356), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n356), .B(new_n687), .C1(new_n352), .C2(new_n346), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n924), .A2(new_n927), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n645), .A2(new_n884), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n919), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n452), .B(new_n728), .C1(new_n734), .C2(KEYINPUT29), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n655), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n687), .A2(KEYINPUT31), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT93), .B1(new_n747), .B2(new_n748), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n741), .A2(new_n744), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n944), .B2(new_n749), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n738), .B2(new_n757), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n844), .B1(new_n929), .B2(new_n931), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT40), .B1(new_n948), .B2(new_n927), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n904), .A2(new_n905), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT18), .B1(new_n443), .B2(new_n641), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n448), .A2(new_n431), .A3(new_n643), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n907), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n954), .B2(new_n912), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT40), .B1(new_n893), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n949), .B1(new_n948), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n453), .A2(new_n946), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n736), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n940), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n205), .B2(new_n766), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n940), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n880), .B1(new_n963), .B2(new_n964), .ZN(G367));
  INV_X1    g0765(.A(new_n763), .ZN(new_n966));
  INV_X1    g0766(.A(new_n704), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n656), .A2(new_n687), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n560), .A2(KEYINPUT106), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n676), .A2(new_n660), .A3(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT106), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n969), .B(new_n972), .C1(new_n660), .C2(new_n688), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT113), .B1(new_n711), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT113), .ZN(new_n975));
  INV_X1    g0775(.A(new_n973), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n707), .A2(new_n709), .B1(new_n700), .B2(new_n702), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(new_n705), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(KEYINPUT44), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n709), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n708), .B1(new_n681), .B2(new_n688), .ZN(new_n981));
  INV_X1    g0781(.A(new_n702), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n701), .B1(new_n696), .B2(new_n698), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n980), .A2(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n705), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(new_n973), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n987), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n711), .A2(new_n973), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n979), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT44), .B1(new_n974), .B2(new_n978), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n967), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n710), .A2(new_n703), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n984), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n693), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n694), .A3(new_n984), .ZN(new_n998));
  AND4_X1   g0798(.A1(new_n762), .A2(new_n997), .A3(new_n735), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n974), .A2(new_n978), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n1002), .A2(new_n704), .A3(new_n979), .A4(new_n991), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n994), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT114), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n994), .A2(new_n1003), .A3(KEYINPUT114), .A4(new_n999), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n966), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n716), .B(KEYINPUT41), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n767), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n967), .A2(new_n973), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT111), .Z(new_n1012));
  INV_X1    g0812(.A(KEYINPUT42), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n710), .A2(new_n1013), .A3(new_n703), .A4(new_n973), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT107), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n710), .A2(new_n703), .A3(new_n973), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT42), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n977), .A2(KEYINPUT107), .A3(new_n1013), .A4(new_n973), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n969), .A2(new_n972), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n660), .B1(new_n1020), .B2(new_n629), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n688), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT108), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1017), .A2(KEYINPUT42), .B1(new_n1021), .B2(new_n688), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT108), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1025), .A2(new_n1026), .A3(new_n1019), .A4(new_n1016), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n594), .A2(new_n688), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1028), .A2(new_n574), .A3(new_n662), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n664), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(KEYINPUT43), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1024), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT109), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1024), .A2(KEYINPUT109), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1030), .B(KEYINPUT43), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT110), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT110), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1036), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1041));
  AOI221_X4 g0841(.A(new_n1012), .B1(new_n1034), .B2(new_n1035), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1012), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1010), .A2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n793), .A2(new_n267), .B1(new_n389), .B2(new_n781), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n396), .B1(new_n798), .B2(G58), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n800), .B2(new_n860), .C1(new_n259), .C2(new_n801), .ZN(new_n1053));
  INV_X1    g0853(.A(G137), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n202), .A2(new_n787), .B1(new_n856), .B2(new_n1054), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(G68), .C2(new_n775), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1050), .A2(new_n1051), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(G283), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n793), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT115), .B(KEYINPUT46), .Z(new_n1060));
  INV_X1    g0860(.A(new_n460), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n797), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n396), .C1(new_n564), .C2(new_n774), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G97), .B2(new_n786), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n852), .A2(new_n801), .B1(new_n800), .B2(new_n810), .ZN(new_n1065));
  AND2_X1   g0865(.A1(KEYINPUT46), .A2(G116), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n815), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n780), .A2(G294), .B1(new_n803), .B2(G317), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1057), .B1(new_n1059), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT47), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n772), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n828), .A2(new_n234), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n825), .B1(new_n209), .B2(new_n364), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n769), .B1(new_n1075), .B2(new_n1076), .C1(new_n1030), .C2(new_n835), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1048), .A2(new_n1079), .ZN(G387));
  NOR2_X1   g0880(.A1(new_n999), .A2(new_n716), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n997), .A2(new_n998), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1081), .B1(new_n763), .B2(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n279), .B1(new_n202), .B2(new_n797), .C1(new_n801), .C2(new_n267), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G159), .B2(new_n807), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n780), .A2(new_n408), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n789), .A2(G68), .B1(new_n803), .B2(G150), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n775), .A2(new_n561), .B1(G97), .B2(new_n786), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n279), .B1(new_n803), .B2(G326), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1058), .A2(new_n774), .B1(new_n797), .B2(new_n809), .ZN(new_n1091));
  INV_X1    g0891(.A(G317), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1092), .A2(new_n801), .B1(new_n800), .B2(new_n813), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G311), .B2(new_n780), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n793), .B2(new_n852), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT48), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT49), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1090), .B1(new_n1061), .B2(new_n787), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1089), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(new_n771), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n231), .A2(G45), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT117), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n253), .A2(new_n256), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n267), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT50), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n717), .B(new_n296), .C1(new_n319), .C2(new_n202), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1105), .B(new_n828), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(G107), .B2(new_n209), .C1(new_n717), .C2(new_n831), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n770), .B(new_n1103), .C1(new_n826), .C2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n700), .A2(new_n702), .A3(new_n824), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1112), .A2(new_n1113), .B1(new_n768), .B2(new_n1082), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1083), .A2(new_n1114), .ZN(G393));
  NAND3_X1  g0915(.A1(new_n994), .A2(new_n768), .A3(new_n1003), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n825), .B1(new_n470), .B2(new_n209), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n828), .B2(new_n238), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n794), .A2(new_n1106), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n396), .B(new_n854), .C1(G68), .C2(new_n798), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n775), .A2(G77), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n267), .B2(new_n781), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G143), .B2(new_n803), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n259), .A2(new_n800), .B1(new_n801), .B2(new_n389), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT51), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1119), .A2(new_n1120), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n810), .A2(new_n801), .B1(new_n800), .B2(new_n1092), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT118), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT52), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n279), .B1(new_n798), .B2(G283), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1061), .B2(new_n774), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G107), .B2(new_n786), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G294), .A2(new_n789), .B1(new_n780), .B2(G303), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n813), .C2(new_n856), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1126), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n770), .B(new_n1118), .C1(new_n1135), .C2(new_n771), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n835), .B2(new_n973), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT119), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n999), .B1(new_n994), .B2(new_n1003), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n716), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1116), .B(new_n1137), .C1(new_n1143), .C2(new_n1144), .ZN(G390));
  INV_X1    g0945(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n724), .A2(new_n726), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n688), .A3(new_n844), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n932), .B1(new_n1148), .B2(new_n923), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT120), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n881), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n893), .B2(new_n955), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1146), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n900), .A2(new_n913), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n922), .B1(new_n727), .B2(new_n844), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(KEYINPUT121), .C1(new_n1157), .C2(new_n932), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n761), .A2(new_n844), .A3(new_n933), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n927), .A2(KEYINPUT39), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n917), .A3(new_n916), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n882), .B1(new_n924), .B2(new_n933), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1159), .B(new_n1160), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n946), .A2(new_n736), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n452), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n938), .A2(new_n655), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n933), .B1(new_n761), .B2(new_n844), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n946), .A2(new_n947), .A3(new_n736), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n924), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n842), .A2(new_n843), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n946), .A2(new_n736), .A3(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1160), .B(new_n1157), .C1(new_n933), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1167), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n898), .A2(new_n918), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n845), .B1(new_n729), .B2(new_n733), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n922), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n881), .B1(new_n1177), .B2(new_n932), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1175), .A2(new_n1178), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1169), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1164), .B(new_n1174), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n765), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(KEYINPUT122), .A3(new_n765), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1174), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1164), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1184), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n767), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1175), .A2(new_n822), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n849), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n769), .B1(new_n408), .B2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT54), .B(G143), .Z(new_n1195));
  NAND2_X1  g0995(.A1(new_n794), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n798), .A2(G150), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT53), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n396), .B(new_n1198), .C1(G137), .C2(new_n780), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n775), .A2(G159), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n267), .B2(new_n787), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G125), .B2(new_n803), .ZN(new_n1202));
  INV_X1    g1002(.A(G128), .ZN(new_n1203));
  INV_X1    g1003(.A(G132), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1203), .A2(new_n800), .B1(new_n801), .B2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT123), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1196), .A2(new_n1199), .A3(new_n1202), .A4(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n793), .A2(new_n470), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n456), .A2(new_n801), .B1(new_n800), .B2(new_n1058), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n279), .B(new_n1209), .C1(G87), .C2(new_n815), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n786), .A2(G68), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n780), .A2(G107), .B1(new_n803), .B2(G294), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1121), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1194), .B1(new_n1214), .B2(new_n771), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1191), .B1(new_n1192), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1190), .A2(new_n1216), .ZN(G378));
  INV_X1    g1017(.A(new_n1167), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1181), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n928), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n357), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1171), .B1(new_n1221), .B2(new_n930), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n639), .A2(KEYINPUT31), .B1(new_n687), .B2(new_n756), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(new_n945), .ZN(new_n1224));
  OAI21_X1  g1024(.A(G330), .B1(new_n1224), .B2(new_n956), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n949), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n315), .B(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n313), .A2(new_n884), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1229), .B(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1226), .B1(new_n949), .B2(new_n1225), .ZN(new_n1234));
  AND4_X1   g1034(.A1(new_n934), .A2(new_n1234), .A3(new_n919), .A4(new_n936), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n935), .B1(new_n1162), .B2(new_n882), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1236), .B2(new_n934), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1233), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n949), .A2(new_n1225), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n937), .A2(new_n1226), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1236), .A2(new_n934), .A3(new_n1234), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1232), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1219), .A2(new_n1238), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1219), .A2(new_n1238), .A3(new_n1242), .A4(KEYINPUT57), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n765), .A3(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1238), .A2(new_n1242), .A3(new_n768), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n769), .B1(G50), .B2(new_n1193), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G50), .B1(new_n278), .B2(new_n295), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n470), .A2(new_n781), .B1(new_n790), .B2(new_n364), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G283), .B2(new_n803), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n295), .B(new_n396), .C1(new_n797), .C2(new_n202), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n801), .A2(new_n564), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(G116), .C2(new_n807), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n775), .A2(G68), .B1(G58), .B2(new_n786), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT58), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1250), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n798), .A2(new_n1195), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1203), .B2(new_n801), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n775), .A2(G150), .B1(G137), .B2(new_n789), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1204), .B2(new_n781), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1261), .B(new_n1263), .C1(G125), .C2(new_n807), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(KEYINPUT59), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n803), .A2(G124), .ZN(new_n1267));
  AOI211_X1 g1067(.A(G33), .B(G41), .C1(new_n786), .C2(G159), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT59), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1267), .B(new_n1268), .C1(new_n1264), .C2(new_n1269), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1259), .B1(new_n1258), .B2(new_n1257), .C1(new_n1266), .C2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1249), .B1(new_n1271), .B2(new_n771), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1231), .B2(new_n823), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1248), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1247), .A2(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n932), .A2(new_n822), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n769), .B1(G68), .B2(new_n1193), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n801), .A2(new_n1054), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n279), .B1(new_n800), .B2(new_n1204), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1279), .B(new_n1280), .C1(G159), .C2(new_n815), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n775), .A2(G50), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n789), .A2(G150), .B1(new_n803), .B2(G128), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n780), .A2(new_n1195), .B1(new_n786), .B2(G58), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1058), .A2(new_n801), .B1(new_n800), .B2(new_n809), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n279), .B(new_n1286), .C1(G97), .C2(new_n815), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n775), .A2(new_n561), .B1(G77), .B2(new_n786), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n780), .A2(new_n460), .B1(new_n803), .B2(G303), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n793), .A2(new_n564), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1285), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1278), .B1(new_n1292), .B2(new_n771), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1276), .A2(new_n768), .B1(new_n1277), .B2(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1174), .A2(new_n1009), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1276), .A2(new_n1218), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(G381));
  NOR2_X1   g1097(.A1(G375), .A2(G378), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1078), .B1(new_n1010), .B2(new_n1047), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1116), .A2(new_n1137), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT119), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1302), .B2(new_n1142), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  NOR4_X1   g1104(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1298), .A2(new_n1304), .A3(new_n1305), .ZN(G407));
  NAND2_X1  g1106(.A1(new_n686), .A2(G213), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1298), .A2(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(KEYINPUT125), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1111(.A1(G387), .A2(G390), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(G393), .B(G396), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1247), .A2(G378), .A3(new_n1274), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1248), .B(new_n1273), .C1(new_n1243), .C2(new_n1009), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1190), .A3(new_n1216), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1307), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1170), .A2(new_n1173), .A3(new_n1167), .A4(KEYINPUT60), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1186), .A2(new_n765), .A3(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1296), .A2(KEYINPUT60), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1294), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(new_n848), .A3(new_n869), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G384), .B(new_n1294), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1318), .B1(new_n1323), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1308), .A2(KEYINPUT126), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1328), .A2(new_n1329), .A3(new_n1332), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1308), .A2(G2897), .ZN(new_n1334));
  XOR2_X1   g1134(.A(new_n1333), .B(new_n1334), .Z(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1308), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1330), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(KEYINPUT63), .A3(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1317), .A2(new_n1331), .A3(new_n1336), .A4(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1337), .A2(new_n1341), .A3(new_n1338), .ZN(new_n1342));
  XOR2_X1   g1142(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1343));
  XNOR2_X1  g1143(.A(new_n1333), .B(new_n1334), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1343), .B1(new_n1337), .B2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1341), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1342), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1340), .B1(new_n1347), .B2(new_n1317), .ZN(G405));
  NAND3_X1  g1148(.A1(G375), .A2(new_n1190), .A3(new_n1216), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1319), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1314), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1351), .B1(new_n1304), .B2(new_n1352), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1353), .A2(new_n1354), .A3(new_n1330), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1330), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1350), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1338), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1353), .A2(new_n1354), .A3(new_n1330), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1358), .A2(new_n1319), .A3(new_n1349), .A4(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1357), .A2(new_n1360), .ZN(G402));
endmodule


