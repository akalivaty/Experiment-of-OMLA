//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n223), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n219), .A2(new_n220), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G58), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  AND2_X1   g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OR2_X1    g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT66), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G222), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n254), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n251), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n248), .B2(new_n249), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n251), .A2(new_n269), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(G226), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  XOR2_X1   g0075(.A(KEYINPUT8), .B(G58), .Z(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n276), .A2(new_n278), .B1(G150), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n280), .A2(new_n281), .B1(G20), .B2(new_n203), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(new_n281), .B2(new_n280), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n224), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n225), .A3(G1), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n285), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n202), .B1(new_n267), .B2(G20), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(new_n290), .B1(new_n202), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(G169), .B1(new_n264), .B2(new_n273), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n275), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G200), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n264), .B2(new_n273), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT9), .B1(new_n286), .B2(new_n291), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n274), .A2(new_n300), .B1(new_n301), .B2(new_n292), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n264), .A2(new_n273), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n304), .A2(G190), .B1(new_n293), .B2(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n297), .A2(new_n298), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n295), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT16), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n252), .A2(new_n225), .A3(new_n253), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT7), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n253), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n208), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G58), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n208), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n317), .B2(new_n201), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n279), .A2(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n310), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT7), .B1(new_n324), .B2(new_n225), .ZN(new_n325));
  NOR4_X1   g0125(.A1(new_n322), .A2(new_n323), .A3(new_n312), .A4(G20), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n320), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n321), .A2(new_n329), .A3(new_n285), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n267), .A2(G20), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n276), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT71), .ZN(new_n333));
  INV_X1    g0133(.A(new_n285), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n287), .A2(G1), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G20), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n332), .B2(KEYINPUT71), .ZN(new_n338));
  INV_X1    g0138(.A(new_n276), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n333), .A2(new_n338), .B1(new_n288), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT18), .ZN(new_n342));
  INV_X1    g0142(.A(G226), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G1698), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n344), .B1(G223), .B2(G1698), .C1(new_n322), .C2(new_n323), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G87), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n251), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n250), .A2(G232), .A3(new_n268), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n270), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(G169), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n250), .B1(new_n345), .B2(new_n346), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n270), .A2(new_n349), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n352), .A2(new_n353), .A3(G179), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n341), .A2(new_n342), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n342), .B1(new_n341), .B2(new_n355), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n348), .A2(new_n300), .A3(new_n350), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n296), .B1(new_n352), .B2(new_n353), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n330), .A2(new_n340), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n330), .A2(new_n361), .A3(KEYINPUT17), .A4(new_n340), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n364), .A2(KEYINPUT72), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT72), .B1(new_n364), .B2(new_n365), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n358), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n278), .A2(G77), .B1(G20), .B2(new_n208), .ZN(new_n370));
  INV_X1    g0170(.A(new_n279), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n202), .B2(new_n371), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n372), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT11), .B1(new_n372), .B2(new_n285), .ZN(new_n374));
  OR3_X1    g0174(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT69), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n288), .A2(new_n208), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT12), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT69), .B1(new_n373), .B2(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n337), .A2(KEYINPUT68), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n289), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(G68), .A3(new_n331), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n375), .A2(new_n377), .A3(new_n378), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G97), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n254), .A2(G232), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n386), .B1(new_n387), .B2(new_n259), .C1(new_n343), .C2(new_n260), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n251), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n271), .B1(G238), .B2(new_n272), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n389), .B2(new_n391), .ZN(new_n393));
  OAI21_X1  g0193(.A(G200), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(G190), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n385), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G169), .B1(new_n392), .B2(new_n393), .ZN(new_n401));
  NAND2_X1  g0201(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n396), .A2(new_n397), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(G169), .A3(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n396), .A2(G179), .A3(new_n397), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n400), .B1(new_n408), .B2(new_n384), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n382), .A2(G77), .A3(new_n331), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n288), .A2(new_n262), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n339), .A2(new_n371), .B1(new_n225), .B2(new_n262), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n225), .A2(G33), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n285), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n410), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n387), .A2(G1698), .B1(new_n418), .B2(new_n254), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n257), .B2(G238), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(new_n250), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n271), .B1(G244), .B2(new_n272), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G169), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n417), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G179), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n426), .A3(new_n422), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n296), .B1(new_n421), .B2(new_n422), .ZN(new_n430));
  OAI211_X1 g0230(.A(G190), .B(new_n422), .C1(new_n420), .C2(new_n250), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n417), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n309), .A2(new_n369), .A3(new_n409), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n267), .A2(G33), .ZN(new_n437));
  AND4_X1   g0237(.A1(G116), .A2(new_n379), .A3(new_n381), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G283), .ZN(new_n439));
  INV_X1    g0239(.A(G97), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n225), .C1(G33), .C2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G20), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n285), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT20), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n444), .A2(new_n445), .ZN(new_n447));
  INV_X1    g0247(.A(new_n335), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n446), .A2(new_n447), .B1(new_n448), .B2(new_n443), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n438), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G41), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n267), .B(G45), .C1(new_n451), .C2(KEYINPUT5), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G41), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT74), .A3(new_n267), .A4(G45), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(KEYINPUT5), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(G270), .A3(new_n250), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n452), .A2(new_n453), .B1(KEYINPUT5), .B2(new_n451), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(new_n266), .A3(new_n457), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT77), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n259), .A2(G257), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G264), .A2(G1698), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n252), .A2(new_n253), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G303), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n322), .A2(new_n323), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n465), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G257), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1698), .ZN(new_n473));
  INV_X1    g0273(.A(new_n467), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n473), .A2(new_n474), .B1(new_n322), .B2(new_n323), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n252), .A2(G303), .A3(new_n253), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(KEYINPUT77), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT78), .B1(new_n478), .B2(new_n251), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT78), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n480), .B(new_n250), .C1(new_n471), .C2(new_n477), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n464), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n450), .B1(new_n482), .B2(new_n300), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n468), .A2(new_n470), .A3(new_n465), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT77), .B1(new_n475), .B2(new_n476), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n251), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n480), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n478), .A2(KEYINPUT78), .A3(new_n251), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n463), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n296), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n436), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n438), .A2(new_n449), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n489), .B2(G190), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n482), .A2(G200), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n487), .A2(new_n488), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n497), .A3(G179), .A4(new_n464), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n482), .A2(new_n492), .A3(G169), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT21), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n482), .A2(new_n492), .A3(new_n502), .A4(G169), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  AND2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT73), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT6), .A2(G97), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(G107), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n418), .A2(KEYINPUT73), .A3(KEYINPUT6), .A4(G97), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n515));
  OAI21_X1  g0315(.A(G107), .B1(new_n325), .B2(new_n326), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n334), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n288), .A2(new_n440), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n289), .A2(new_n437), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n440), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G244), .B(new_n259), .C1(new_n322), .C2(new_n323), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n439), .A4(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(new_n251), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n459), .A2(G257), .A3(new_n250), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n462), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n424), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n529), .A2(new_n462), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n251), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n426), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n521), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n517), .A2(new_n520), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(G190), .A3(new_n533), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n296), .B1(new_n532), .B2(new_n533), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(KEYINPUT75), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(new_n259), .C1(new_n322), .C2(new_n323), .ZN(new_n542));
  OAI211_X1 g0342(.A(G257), .B(G1698), .C1(new_n322), .C2(new_n323), .ZN(new_n543));
  INV_X1    g0343(.A(G294), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n543), .C1(new_n277), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n251), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n459), .A2(G264), .A3(new_n250), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(new_n462), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n424), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n251), .B1(new_n461), .B2(new_n457), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G264), .B1(new_n545), .B2(new_n251), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n426), .A3(new_n462), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n225), .A2(KEYINPUT80), .A3(G87), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT22), .B1(new_n324), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n553), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n254), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n278), .A2(G116), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT82), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(KEYINPUT23), .B1(new_n561), .B2(KEYINPUT24), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n560), .A2(KEYINPUT23), .B1(new_n225), .B2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(new_n418), .A3(KEYINPUT81), .A4(G20), .ZN(new_n565));
  AND4_X1   g0365(.A1(new_n559), .A2(new_n562), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n558), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n561), .A2(KEYINPUT24), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n558), .A2(new_n568), .A3(new_n566), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n334), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n519), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT25), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n336), .B2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n418), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n573), .A2(G107), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n549), .B(new_n552), .C1(new_n572), .C2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n571), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n568), .B1(new_n558), .B2(new_n566), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n285), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(G200), .B1(new_n551), .B2(new_n462), .ZN(new_n583));
  AND4_X1   g0383(.A1(new_n300), .A2(new_n546), .A3(new_n547), .A4(new_n462), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n577), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n267), .A2(new_n265), .A3(G45), .ZN(new_n586));
  INV_X1    g0386(.A(G45), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n211), .B1(new_n587), .B2(G1), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n250), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n209), .A2(G1698), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n322), .B2(new_n323), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT76), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n254), .A2(G244), .A3(G1698), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT76), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n254), .A2(new_n595), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G116), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n590), .B1(new_n598), .B2(new_n251), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(G169), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n426), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n254), .A2(new_n225), .A3(G68), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n225), .B1(new_n386), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n508), .A2(new_n210), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n414), .B2(new_n440), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n285), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n413), .A2(new_n288), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n609), .B(new_n610), .C1(new_n413), .C2(new_n519), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n600), .A2(new_n601), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n599), .A2(G190), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n289), .A2(G87), .A3(new_n437), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n609), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n613), .B(new_n615), .C1(new_n296), .C2(new_n599), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n579), .A2(new_n585), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n435), .A2(new_n505), .A3(new_n541), .A4(new_n617), .ZN(G372));
  OAI21_X1  g0418(.A(new_n407), .B1(new_n401), .B2(new_n403), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n402), .B1(new_n405), .B2(G169), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n384), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n400), .B2(new_n428), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n367), .B2(new_n366), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n358), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n303), .A2(new_n308), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n295), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n435), .ZN(new_n627));
  INV_X1    g0427(.A(new_n612), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n504), .A2(new_n579), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n615), .B1(new_n296), .B2(new_n599), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT83), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n615), .B(KEYINPUT83), .C1(new_n296), .C2(new_n599), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n613), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n585), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n541), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n628), .B1(new_n629), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n521), .A2(new_n531), .A3(new_n534), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n634), .A2(new_n638), .A3(new_n612), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n612), .A2(new_n616), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n535), .ZN(new_n641));
  MUX2_X1   g0441(.A(new_n639), .B(new_n641), .S(KEYINPUT26), .Z(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n627), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n626), .A2(new_n644), .ZN(G369));
  INV_X1    g0445(.A(KEYINPUT84), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n335), .A2(new_n225), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(KEYINPUT27), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(new_n646), .A3(KEYINPUT27), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(G213), .B1(new_n647), .B2(KEYINPUT27), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n505), .B1(new_n492), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n655), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n504), .A2(new_n450), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT85), .Z(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n572), .B2(new_n578), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n579), .A2(new_n585), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n579), .A2(new_n657), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n664), .A2(KEYINPUT87), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n661), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n504), .A2(new_n655), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n579), .A2(new_n655), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n673), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n221), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n605), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n228), .B2(new_n682), .ZN(new_n685));
  XOR2_X1   g0485(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n686));
  XNOR2_X1  g0486(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n655), .B1(new_n637), .B2(new_n642), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n640), .A2(KEYINPUT26), .A3(new_n535), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n655), .B1(new_n637), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n689), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n537), .A2(new_n536), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n638), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n579), .A2(new_n585), .A3(new_n612), .A4(new_n616), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n657), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n551), .B(new_n599), .C1(new_n479), .C2(new_n481), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n464), .A2(new_n532), .A3(G179), .A4(new_n533), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n460), .A2(G179), .A3(new_n462), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n528), .A2(new_n706), .A3(new_n530), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n599), .A2(new_n551), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n497), .A3(new_n708), .A4(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n532), .A2(new_n533), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n599), .A2(G179), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n482), .A2(new_n710), .A3(new_n548), .A4(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n705), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n713), .A2(new_n714), .A3(new_n655), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n713), .B2(new_n655), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n505), .A2(new_n701), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT89), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n718), .B1(new_n717), .B2(G330), .ZN(new_n721));
  NOR4_X1   g0521(.A1(new_n690), .A2(new_n694), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n687), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n287), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n267), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n681), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n224), .B1(G20), .B2(new_n424), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n426), .A2(new_n296), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT95), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n225), .B1(new_n735), .B2(G190), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(KEYINPUT98), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(KEYINPUT98), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n440), .ZN(new_n740));
  NAND3_X1  g0540(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT94), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n208), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n300), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n202), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n426), .A2(G200), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G20), .A3(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n225), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n749), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n750), .A2(new_n316), .B1(new_n752), .B2(new_n262), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT93), .Z(new_n754));
  NOR4_X1   g0554(.A1(new_n740), .A2(new_n745), .A3(new_n748), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n735), .A2(new_n751), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G159), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n225), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G87), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n300), .A3(G200), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n764), .B(new_n254), .C1(new_n418), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n760), .B1(new_n767), .B2(KEYINPUT97), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n755), .B(new_n768), .C1(KEYINPUT97), .C2(new_n767), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT99), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT33), .B(G317), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G326), .A2(new_n746), .B1(new_n743), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n757), .A2(G329), .ZN(new_n773));
  INV_X1    g0573(.A(G322), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n324), .B1(new_n750), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n752), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(G311), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n765), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n763), .A2(G303), .B1(new_n778), .B2(G283), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n772), .A2(new_n773), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n739), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(G294), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n769), .B2(KEYINPUT99), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n733), .B1(new_n770), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n732), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n254), .A2(new_n221), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT90), .Z(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G355), .B1(new_n442), .B2(new_n680), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n680), .A2(new_n254), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT91), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n228), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n246), .A2(new_n587), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n728), .B(new_n784), .C1(new_n788), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT100), .ZN(new_n798));
  INV_X1    g0598(.A(new_n787), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n659), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT101), .Z(new_n801));
  XNOR2_X1  g0601(.A(new_n660), .B(KEYINPUT85), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n728), .B1(new_n659), .B2(G330), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(G396));
  OAI22_X1  g0604(.A1(new_n430), .A2(new_n432), .B1(new_n417), .B2(new_n657), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n428), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n425), .A2(new_n427), .A3(new_n657), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n688), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n720), .A2(new_n721), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n727), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n733), .A2(new_n786), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n727), .B1(new_n814), .B2(G77), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n778), .A2(G68), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n816), .B(new_n254), .C1(new_n202), .C2(new_n762), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G132), .B2(new_n757), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n739), .B2(new_n316), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT102), .Z(new_n820));
  INV_X1    g0620(.A(new_n750), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G143), .B1(new_n776), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(G150), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n744), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G137), .B2(new_n746), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT34), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n210), .A2(new_n765), .B1(new_n762), .B2(new_n418), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n324), .B1(new_n752), .B2(new_n442), .C1(new_n544), .C2(new_n750), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G311), .C2(new_n757), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n744), .C1(new_n469), .C2(new_n747), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n820), .A2(new_n826), .B1(new_n740), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n815), .B1(new_n832), .B2(new_n732), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n809), .B2(new_n786), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n813), .A2(new_n834), .ZN(G384));
  AOI21_X1  g0635(.A(new_n653), .B1(new_n330), .B2(new_n340), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n368), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT104), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n341), .A2(new_n355), .B1(new_n838), .B2(KEYINPUT37), .ZN(new_n839));
  INV_X1    g0639(.A(new_n653), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n341), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AND4_X1   g0643(.A1(new_n362), .A2(new_n839), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n330), .A2(new_n340), .A3(new_n361), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n836), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n843), .B1(new_n846), .B2(new_n839), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n837), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT38), .B1(new_n837), .B2(new_n848), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT105), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n364), .A2(new_n854), .A3(new_n365), .ZN(new_n855));
  INV_X1    g0655(.A(new_n357), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n341), .A2(new_n342), .A3(new_n355), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n854), .B1(new_n364), .B2(new_n365), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n836), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n848), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n837), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n851), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n853), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n408), .A2(new_n384), .A3(new_n657), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n358), .A2(new_n840), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n384), .A2(new_n655), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n621), .A2(new_n399), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n384), .B(new_n655), .C1(new_n408), .C2(new_n400), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n643), .A2(new_n657), .A3(new_n809), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n807), .B(KEYINPUT103), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n849), .A2(new_n850), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n872), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n627), .B1(new_n690), .B2(new_n694), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n626), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n884), .B(new_n886), .Z(new_n887));
  NAND2_X1  g0687(.A1(new_n713), .A2(new_n655), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT31), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n713), .A2(new_n714), .A3(new_n655), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT106), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n541), .A2(new_n617), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(new_n496), .A3(new_n504), .A4(new_n657), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n892), .B1(new_n891), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n627), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT107), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n717), .A2(KEYINPUT106), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n808), .B1(new_n874), .B2(new_n875), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n904), .B2(new_n881), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n900), .B1(new_n863), .B2(new_n864), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n897), .A2(new_n906), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(G330), .B1(new_n899), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n908), .B2(new_n899), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n887), .A2(new_n910), .B1(new_n267), .B2(new_n724), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n887), .B2(new_n910), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(G116), .A3(new_n226), .A4(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OR3_X1    g0716(.A1(new_n228), .A2(new_n262), .A3(new_n317), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n202), .A2(G68), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n267), .B(G13), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OR3_X1    g0719(.A1(new_n912), .A2(new_n916), .A3(new_n919), .ZN(G367));
  OAI21_X1  g0720(.A(new_n699), .B1(new_n536), .B2(new_n657), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n638), .A2(new_n655), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n671), .A2(new_n674), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n535), .B1(new_n921), .B2(new_n579), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n924), .A2(KEYINPUT42), .B1(new_n657), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n657), .A2(new_n615), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(new_n612), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n612), .A3(new_n634), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n928), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n925), .A2(new_n927), .A3(new_n934), .A4(new_n933), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n673), .A2(new_n923), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n939), .B(new_n940), .Z(new_n941));
  XOR2_X1   g0741(.A(new_n681), .B(KEYINPUT41), .Z(new_n942));
  NAND3_X1  g0742(.A1(new_n675), .A2(new_n677), .A3(new_n923), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  INV_X1    g0746(.A(new_n923), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n678), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT44), .B1(new_n678), .B2(new_n947), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n945), .A2(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(new_n673), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n673), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n671), .A2(new_n674), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n675), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n661), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n802), .A2(new_n675), .A3(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n951), .A2(new_n952), .A3(new_n722), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n942), .B1(new_n959), .B2(new_n722), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n725), .B(KEYINPUT108), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n941), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n788), .ZN(new_n964));
  INV_X1    g0764(.A(new_n413), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n680), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n793), .A2(new_n238), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n728), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n781), .A2(G68), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n823), .B2(new_n750), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT110), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n324), .B1(new_n776), .B2(G50), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n316), .B2(new_n762), .C1(new_n262), .C2(new_n765), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT111), .B(G137), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n757), .B2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G143), .A2(new_n746), .B1(new_n743), .B2(G159), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT112), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT46), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n762), .B2(new_n442), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n744), .C2(new_n544), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT109), .Z(new_n984));
  INV_X1    g0784(.A(G311), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n747), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n254), .B1(new_n776), .B2(G283), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n440), .B2(new_n765), .C1(new_n469), .C2(new_n750), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(G317), .C2(new_n757), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n984), .B(new_n989), .C1(new_n418), .C2(new_n739), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n979), .A2(KEYINPUT47), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n732), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT47), .B1(new_n979), .B2(new_n990), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n968), .B1(new_n799), .B2(new_n932), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n963), .A2(new_n994), .ZN(G387));
  NAND2_X1  g0795(.A1(new_n672), .A2(new_n787), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n793), .B1(new_n235), .B2(new_n587), .ZN(new_n997));
  INV_X1    g0797(.A(new_n790), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n683), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n339), .B2(G50), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n276), .A2(new_n1000), .A3(new_n202), .ZN(new_n1003));
  AOI21_X1  g0803(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1002), .A2(new_n683), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n999), .A2(new_n1005), .B1(new_n418), .B2(new_n680), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n727), .B1(new_n1006), .B2(new_n964), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n781), .A2(new_n965), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n262), .A2(new_n762), .B1(new_n765), .B2(new_n440), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n254), .B1(new_n752), .B2(new_n208), .C1(new_n202), .C2(new_n750), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G150), .C2(new_n757), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G159), .A2(new_n746), .B1(new_n743), .B2(new_n276), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n821), .A2(G317), .B1(new_n776), .B2(G303), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n744), .B2(new_n985), .C1(new_n774), .C2(new_n747), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT48), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n781), .A2(G283), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n763), .A2(G294), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT49), .Z(new_n1022));
  INV_X1    g0822(.A(G326), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n324), .B1(new_n442), .B2(new_n765), .C1(new_n756), .C2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1013), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1007), .B1(new_n1025), .B2(new_n732), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n958), .A2(new_n962), .B1(new_n996), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n958), .A2(new_n722), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n681), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n958), .A2(new_n722), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(G393));
  NAND2_X1  g0831(.A1(new_n951), .A2(new_n952), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n1028), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n681), .A3(new_n959), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n951), .A2(new_n952), .A3(new_n962), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n788), .B1(new_n440), .B2(new_n221), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n243), .B2(new_n793), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n781), .A2(G77), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n202), .B2(new_n744), .C1(new_n339), .C2(new_n752), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT114), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n746), .A2(G150), .B1(G159), .B2(new_n821), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT51), .Z(new_n1042));
  OAI221_X1 g0842(.A(new_n254), .B1(new_n765), .B2(new_n210), .C1(new_n208), .C2(new_n762), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n757), .B2(G143), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n746), .A2(G317), .B1(G311), .B2(new_n821), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n254), .B1(new_n776), .B2(G294), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n418), .B2(new_n765), .C1(new_n830), .C2(new_n762), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G322), .B2(new_n757), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n442), .B2(new_n739), .C1(new_n469), .C2(new_n744), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1045), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n728), .B(new_n1037), .C1(new_n1052), .C2(new_n732), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n799), .B2(new_n923), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1035), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1034), .A2(new_n1055), .ZN(G390));
  AND3_X1   g0856(.A1(new_n901), .A2(G330), .A3(new_n903), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n902), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n878), .A2(new_n879), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n876), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1061), .A2(new_n869), .B1(new_n853), .B2(new_n866), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n865), .A2(new_n869), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n637), .A2(new_n692), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(new_n657), .A3(new_n806), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n807), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1063), .B1(new_n1066), .B2(new_n876), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1059), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n867), .B1(new_n870), .B2(new_n880), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1067), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n809), .B(new_n876), .C1(new_n720), .C2(new_n721), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n901), .A2(G330), .A3(new_n809), .A4(new_n903), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n877), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1071), .A2(new_n1076), .A3(new_n807), .A4(new_n1065), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n809), .B1(new_n720), .B2(new_n721), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1078), .A2(new_n877), .B1(new_n1057), .B2(new_n902), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1060), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1057), .A2(new_n627), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n885), .A2(new_n626), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1074), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1068), .A2(new_n1072), .A3(new_n1084), .A4(new_n1081), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n681), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1073), .A2(new_n962), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n727), .B1(new_n814), .B2(new_n276), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT115), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1038), .B1(new_n442), .B2(new_n750), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT116), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n254), .B1(new_n776), .B2(G97), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n764), .A3(new_n816), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G294), .B2(new_n757), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G107), .A2(new_n743), .B1(new_n746), .B2(G283), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n781), .A2(G159), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n324), .B1(new_n776), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(G132), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1102), .B1(new_n202), .B2(new_n765), .C1(new_n1103), .C2(new_n750), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G125), .B2(new_n757), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n762), .A2(new_n823), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G128), .A2(new_n746), .B1(new_n743), .B2(new_n975), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1099), .A2(new_n1105), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1098), .A2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1091), .B1(new_n733), .B2(new_n1110), .C1(new_n868), .C2(new_n786), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1089), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(KEYINPUT117), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(KEYINPUT117), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1088), .B1(new_n1113), .B2(new_n1114), .ZN(G378));
  INV_X1    g0915(.A(KEYINPUT57), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1087), .B2(new_n1084), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT121), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n905), .A2(new_n907), .A3(G330), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT120), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n905), .A2(new_n907), .A3(new_n1121), .A4(G330), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n293), .A2(new_n653), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n309), .A2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n295), .B(new_n1125), .C1(new_n303), .C2(new_n308), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n295), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n299), .A2(KEYINPUT10), .A3(new_n302), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1125), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n309), .A2(new_n1126), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n1123), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1129), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AND4_X1   g0938(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .A4(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n905), .A2(new_n907), .A3(G330), .A4(new_n1137), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1137), .B1(new_n1119), .B2(KEYINPUT120), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n1122), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n884), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1139), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1120), .A2(new_n1122), .A3(new_n1138), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1141), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n884), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1117), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT122), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1117), .B(KEYINPUT122), .C1(new_n1145), .C2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1144), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1148), .A2(new_n884), .A3(new_n1149), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1156), .A2(new_n1157), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n681), .B1(new_n1158), .B2(KEYINPUT57), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n961), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1138), .A2(new_n785), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n727), .B1(new_n814), .B2(G50), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n316), .A2(new_n765), .B1(new_n762), .B2(new_n262), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n254), .A2(G41), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n418), .B2(new_n750), .C1(new_n413), .C2(new_n752), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G283), .C2(new_n757), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G97), .A2(new_n743), .B1(new_n746), .B2(G116), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n969), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT58), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n778), .C2(G159), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT118), .B(G124), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n744), .A2(new_n1103), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n746), .A2(G125), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n821), .A2(G128), .B1(new_n776), .B2(G137), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n762), .C2(new_n1100), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1174), .B(new_n1177), .C1(new_n781), .C2(G150), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1172), .B1(new_n756), .B2(new_n1173), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1178), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1170), .B1(new_n1165), .B2(new_n1171), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(new_n733), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1163), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1161), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1160), .A2(new_n1191), .ZN(G375));
  INV_X1    g0992(.A(new_n942), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1083), .B(new_n1077), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1085), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n877), .A2(new_n785), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n727), .B1(new_n814), .B2(G68), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n781), .A2(G50), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n743), .A2(new_n1101), .B1(new_n821), .B2(new_n975), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1103), .B2(new_n747), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT123), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n324), .B1(new_n776), .B2(G150), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n763), .A2(G159), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n316), .C2(new_n765), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G128), .B2(new_n757), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1198), .A2(new_n1202), .A3(new_n1203), .A4(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n262), .A2(new_n765), .B1(new_n762), .B2(new_n440), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n324), .B1(new_n752), .B2(new_n418), .C1(new_n830), .C2(new_n750), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G303), .C2(new_n757), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G116), .A2(new_n743), .B1(new_n746), .B2(G294), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1008), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1208), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1197), .B1(new_n1214), .B2(new_n732), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1081), .A2(new_n962), .B1(new_n1196), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1195), .A2(new_n1216), .ZN(G381));
  NOR4_X1   g1017(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1218));
  INV_X1    g1018(.A(G390), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1088), .A2(new_n1089), .A3(new_n1111), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OR3_X1    g1021(.A1(G375), .A2(new_n1221), .A3(G387), .ZN(G407));
  NAND2_X1  g1022(.A1(new_n654), .A2(G213), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G375), .C2(new_n1225), .ZN(G409));
  AOI21_X1  g1026(.A(new_n682), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1194), .A2(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT125), .B1(new_n1194), .B2(new_n1228), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n721), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n808), .B1(new_n1232), .B2(new_n719), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1058), .B1(new_n1233), .B2(new_n876), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1066), .B1(new_n877), .B2(new_n1075), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1234), .A2(new_n1060), .B1(new_n1071), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(KEYINPUT60), .A4(new_n1083), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1231), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1230), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G384), .B1(new_n1240), .B2(new_n1216), .ZN(new_n1241));
  INV_X1    g1041(.A(G384), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1216), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(new_n1230), .C2(new_n1239), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT126), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1224), .B1(new_n1245), .B2(G2897), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1245), .B2(G2897), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1241), .A2(new_n1244), .A3(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1231), .A2(new_n1238), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1229), .A2(new_n1085), .A3(new_n681), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1216), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1242), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1240), .A2(G384), .A3(new_n1216), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1224), .A2(G2897), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT127), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(KEYINPUT127), .B(new_n1255), .C1(new_n1241), .C2(new_n1244), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1248), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1191), .C1(new_n1155), .C2(new_n1159), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n962), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(KEYINPUT124), .A3(new_n1189), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1161), .B2(new_n1190), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1158), .A2(new_n1193), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1220), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1261), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1223), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1260), .B2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G396), .B(G393), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n963), .A2(new_n994), .A3(G390), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G390), .B1(new_n963), .B2(new_n994), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(new_n1219), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1272), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n963), .A2(G390), .A3(new_n994), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1270), .B2(new_n1254), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1224), .B1(new_n1261), .B2(new_n1268), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1254), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1271), .A2(new_n1280), .A3(new_n1282), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1283), .A2(new_n1287), .A3(new_n1284), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1283), .B2(new_n1259), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1286), .B1(new_n1292), .B2(new_n1280), .ZN(G405));
  NAND2_X1  g1093(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1220), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1261), .A3(new_n1254), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1254), .B1(new_n1295), .B2(new_n1261), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1294), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1298), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1280), .A3(new_n1296), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(G402));
endmodule


