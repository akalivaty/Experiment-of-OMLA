//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT66), .B(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n202), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G250), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n209), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G257), .ZN(new_n231));
  INV_X1    g0031(.A(G264), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n228), .B(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n227), .B1(new_n233), .B2(KEYINPUT0), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n219), .B(new_n234), .C1(KEYINPUT0), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n240), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n202), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n225), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n206), .B2(G20), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n260), .B2(new_n202), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G58), .ZN(new_n265));
  OR3_X1    g0065(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT8), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n207), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n259), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT9), .B(new_n261), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n271), .B2(new_n273), .ZN(new_n278));
  INV_X1    g0078(.A(new_n261), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G1), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT69), .B(G45), .Z(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n282), .B1(new_n284), .B2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n285), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT71), .B(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT70), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n293), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G222), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(new_n301), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G223), .A3(G1698), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n305), .C1(new_n211), .C2(new_n304), .ZN(new_n306));
  INV_X1    g0106(.A(new_n289), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n292), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n276), .B(new_n280), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(G190), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT75), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  INV_X1    g0118(.A(new_n316), .ZN(new_n319));
  NOR4_X1   g0119(.A1(new_n310), .A2(new_n312), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n315), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n308), .A2(G179), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n308), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n278), .A2(new_n279), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n272), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n269), .A2(new_n211), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n259), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT11), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n260), .A2(G68), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT78), .ZN(new_n334));
  INV_X1    g0134(.A(G68), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n255), .A2(G20), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(KEYINPUT12), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n336), .A2(KEYINPUT12), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(KEYINPUT79), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(KEYINPUT79), .B2(new_n338), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n332), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n291), .A2(KEYINPUT76), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT76), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n289), .A2(new_n343), .A3(new_n290), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G238), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT77), .B(new_n285), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n346), .B1(new_n342), .B2(new_n344), .ZN(new_n349));
  AOI211_X1 g0149(.A(G1), .B(new_n281), .C1(new_n283), .C2(new_n288), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G97), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n287), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n239), .B1(new_n297), .B2(new_n301), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n302), .A2(G226), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n289), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT13), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n358), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n351), .A4(new_n347), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n362), .A3(G179), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n323), .B1(new_n359), .B2(new_n362), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT14), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g0166(.A(KEYINPUT14), .B(new_n323), .C1(new_n359), .C2(new_n362), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n341), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n341), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n359), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(G200), .B1(new_n359), .B2(new_n362), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n321), .A2(new_n327), .A3(new_n368), .A4(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT80), .B1(new_n294), .B2(G33), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT80), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n287), .A3(KEYINPUT3), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n375), .A2(G33), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G223), .ZN(new_n380));
  INV_X1    g0180(.A(G1698), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n293), .A2(new_n380), .B1(new_n286), .B2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n379), .A2(new_n382), .B1(G33), .B2(G87), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n289), .ZN(new_n384));
  INV_X1    g0184(.A(new_n291), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G232), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n285), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G200), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n285), .A2(new_n386), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(G190), .C1(new_n289), .C2(new_n383), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT84), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n272), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n304), .B2(G20), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(G20), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n296), .B(KEYINPUT82), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n375), .A2(G33), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n398), .B1(new_n405), .B2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT83), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT83), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n335), .B1(new_n400), .B2(new_n404), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n398), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT7), .B1(new_n379), .B2(G20), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n379), .A2(KEYINPUT7), .A3(G20), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT16), .B(new_n397), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n407), .A2(new_n411), .A3(new_n259), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n267), .A2(new_n256), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n267), .B2(new_n260), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n395), .A2(KEYINPUT17), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n411), .A2(new_n259), .A3(new_n415), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n405), .A2(G68), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n397), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n408), .B1(new_n423), .B2(new_n409), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n418), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n392), .A2(new_n394), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n420), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n384), .A2(new_n387), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(G169), .ZN(new_n431));
  INV_X1    g0231(.A(G179), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n430), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n425), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n429), .B1(new_n425), .B2(new_n433), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n262), .A2(new_n328), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n275), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n260), .A2(G77), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G77), .B2(new_n256), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n285), .B1(new_n210), .B2(new_n291), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n355), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n304), .A2(G238), .A3(G1698), .ZN(new_n450));
  INV_X1    g0250(.A(G107), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n449), .B(new_n450), .C1(new_n451), .C2(new_n304), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n445), .B1(new_n452), .B2(new_n307), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n444), .B1(new_n454), .B2(new_n323), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n432), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT73), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n456), .A2(KEYINPUT73), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n454), .A2(G190), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n453), .A2(G200), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n444), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n428), .A2(new_n436), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n374), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n451), .B1(new_n400), .B2(new_n404), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT6), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n353), .A2(new_n451), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n451), .A2(KEYINPUT6), .A3(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n211), .B2(new_n328), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n259), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n256), .A2(new_n353), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n275), .B(new_n256), .C1(G1), .C2(new_n287), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n479), .B2(new_n353), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT86), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n288), .A3(KEYINPUT5), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(KEYINPUT86), .B2(G41), .ZN(new_n485));
  INV_X1    g0285(.A(G45), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G1), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n483), .A2(new_n485), .A3(new_n487), .A4(G274), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n289), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n492), .B2(G257), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n300), .B1(new_n298), .B2(new_n299), .ZN(new_n496));
  OAI211_X1 g0296(.A(G250), .B(G1698), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(KEYINPUT4), .A2(G244), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n302), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n376), .A2(new_n378), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n294), .A2(KEYINPUT81), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT81), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT3), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n505), .A3(G33), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n502), .A2(new_n506), .A3(G244), .A4(new_n448), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT85), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT4), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n507), .B2(new_n509), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n497), .B(new_n501), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n494), .B1(new_n512), .B2(new_n307), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n481), .B1(G190), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n448), .B(new_n500), .C1(new_n495), .C2(new_n496), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n497), .A2(new_n515), .A3(new_n498), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n507), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT85), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n493), .B1(new_n520), .B2(new_n289), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT87), .B1(new_n521), .B2(G200), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT87), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n513), .A2(new_n523), .A3(new_n309), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n514), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n519), .A2(new_n517), .ZN(new_n526));
  INV_X1    g0326(.A(new_n516), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n289), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(G169), .B1(new_n528), .B2(new_n494), .ZN(new_n529));
  OAI211_X1 g0329(.A(G179), .B(new_n493), .C1(new_n520), .C2(new_n289), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n529), .A2(new_n530), .B1(new_n476), .B2(new_n480), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(G250), .B1(new_n486), .B2(G1), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n282), .A2(G45), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n307), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n502), .A2(new_n506), .A3(G244), .A4(G1698), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n502), .A2(new_n506), .A3(G238), .A4(new_n448), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n535), .B1(new_n539), .B2(new_n307), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  AOI211_X1 g0341(.A(G190), .B(new_n535), .C1(new_n539), .C2(new_n307), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT19), .B1(new_n354), .B2(new_n207), .ZN(new_n544));
  NAND3_X1  g0344(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n207), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G87), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n451), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT88), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT88), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n544), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n379), .A2(KEYINPUT89), .A3(new_n207), .A4(G68), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n502), .A2(new_n506), .A3(new_n207), .A4(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT89), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n259), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n438), .A2(new_n256), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G87), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n559), .B(new_n561), .C1(new_n562), .C2(new_n478), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n543), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n479), .A2(new_n438), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n559), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT90), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n560), .B1(new_n558), .B2(new_n259), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(KEYINPUT90), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n540), .A2(G179), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n323), .B2(new_n540), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n564), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n525), .A2(new_n532), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n490), .A2(G270), .A3(new_n289), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n488), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT91), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(KEYINPUT91), .A3(new_n488), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n446), .A2(new_n447), .A3(new_n231), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n232), .A2(new_n381), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n506), .B(new_n502), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT92), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n297), .A2(G303), .A3(new_n301), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n307), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n581), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n287), .A2(G97), .ZN(new_n591));
  AOI21_X1  g0391(.A(G20), .B1(new_n591), .B2(new_n498), .ZN(new_n592));
  INV_X1    g0392(.A(G116), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n207), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n259), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n256), .A2(new_n593), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n479), .B2(new_n593), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n323), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n590), .A2(KEYINPUT21), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n584), .A2(new_n586), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT92), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n307), .A3(new_n587), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(new_n599), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(G179), .A4(new_n581), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT21), .B1(new_n590), .B2(new_n600), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n255), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n451), .A2(G20), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g0412(.A(new_n612), .B(KEYINPUT25), .Z(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(G107), .B2(new_n479), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n611), .B(KEYINPUT23), .ZN(new_n615));
  INV_X1    g0415(.A(new_n538), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n207), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n502), .A2(new_n506), .A3(new_n207), .A4(G87), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT93), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT22), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n562), .A2(KEYINPUT22), .A3(G20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n304), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n619), .B1(new_n618), .B2(KEYINPUT22), .ZN(new_n624));
  OAI211_X1 g0424(.A(KEYINPUT24), .B(new_n617), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n259), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n618), .A2(KEYINPUT22), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT93), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n620), .A3(new_n622), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT24), .B1(new_n629), .B2(new_n617), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n614), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n293), .A2(new_n228), .B1(new_n231), .B2(new_n381), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n379), .A2(new_n632), .B1(G33), .B2(G294), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT94), .B1(new_n633), .B2(new_n289), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n448), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n502), .A2(new_n506), .ZN(new_n636));
  INV_X1    g0436(.A(G294), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n635), .A2(new_n636), .B1(new_n287), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT94), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(new_n307), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n491), .A2(new_n232), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(new_n489), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n634), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n638), .A2(new_n307), .ZN(new_n644));
  INV_X1    g0444(.A(new_n641), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n488), .A3(new_n645), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n643), .A2(new_n323), .B1(new_n432), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n631), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n309), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n634), .A2(new_n370), .A3(new_n640), .A4(new_n642), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n651), .B(new_n614), .C1(new_n630), .C2(new_n626), .ZN(new_n652));
  INV_X1    g0452(.A(new_n605), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n581), .B(new_n370), .C1(new_n588), .C2(new_n589), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(G200), .B1(new_n604), .B2(new_n581), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n609), .A2(new_n648), .A3(new_n652), .A4(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n466), .A2(new_n575), .A3(new_n658), .ZN(G372));
  INV_X1    g0459(.A(new_n327), .ZN(new_n660));
  INV_X1    g0460(.A(new_n321), .ZN(new_n661));
  INV_X1    g0461(.A(new_n435), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n425), .A2(new_n429), .A3(new_n433), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n368), .A2(new_n460), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n419), .A2(new_n427), .A3(new_n373), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n661), .B1(new_n667), .B2(KEYINPUT95), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT95), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n419), .A2(new_n427), .A3(new_n373), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n460), .B2(new_n368), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n671), .B2(new_n664), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n660), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n609), .A2(new_n648), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n652), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n575), .A2(new_n675), .ZN(new_n676));
  AND4_X1   g0476(.A1(KEYINPUT90), .A2(new_n559), .A3(new_n561), .A4(new_n565), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT90), .B1(new_n569), .B2(new_n565), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n573), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI221_X1 g0479(.A(new_n569), .B1(new_n562), .B2(new_n478), .C1(new_n541), .C2(new_n542), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n530), .B1(new_n323), .B2(new_n513), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .A4(new_n481), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT26), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n531), .A2(new_n684), .A3(new_n679), .A4(new_n680), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n465), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n673), .A2(new_n687), .ZN(G369));
  OR3_X1    g0488(.A1(new_n610), .A2(KEYINPUT27), .A3(G20), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT27), .B1(new_n610), .B2(G20), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n653), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n609), .B2(new_n657), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n609), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n631), .A2(new_n693), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n648), .A2(new_n699), .A3(new_n652), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n631), .A2(new_n647), .A3(new_n693), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n652), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n648), .B2(new_n609), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n694), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(new_n708), .ZN(G399));
  NOR2_X1   g0509(.A1(new_n230), .A2(G41), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n547), .A2(new_n451), .A3(new_n593), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n206), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n224), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n581), .B(G179), .C1(new_n588), .C2(new_n589), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n540), .A2(new_n644), .A3(new_n645), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n718), .A2(new_n513), .A3(KEYINPUT30), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n539), .A2(new_n307), .ZN(new_n722));
  INV_X1    g0522(.A(new_n535), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n646), .A2(new_n724), .A3(new_n432), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n521), .A3(new_n590), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n717), .A2(new_n719), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT30), .B1(new_n728), .B2(new_n513), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n716), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n718), .A2(new_n513), .A3(new_n720), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(KEYINPUT96), .A3(new_n721), .A4(new_n726), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n693), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n575), .A2(new_n658), .A3(new_n693), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT31), .B(new_n693), .C1(new_n727), .C2(new_n729), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n715), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n685), .A2(new_n679), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n684), .B1(new_n574), .B2(new_n531), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT97), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n523), .B1(new_n513), .B2(new_n309), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n521), .A2(KEYINPUT87), .A3(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n531), .B1(new_n748), .B2(new_n514), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n707), .A2(new_n574), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT97), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n683), .A2(new_n751), .A3(new_n679), .A4(new_n685), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n745), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n694), .B1(new_n676), .B2(new_n686), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n742), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n714), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(new_n710), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n254), .A2(G20), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G45), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT98), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(G1), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n225), .B1(G20), .B2(new_n323), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n207), .A2(new_n370), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n432), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT100), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(G190), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n265), .B1(new_n211), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT101), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n432), .A2(new_n309), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n769), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(G50), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n780), .B2(new_n779), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT102), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n777), .B(KEYINPUT103), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(G179), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT104), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT104), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  OAI21_X1  g0593(.A(KEYINPUT32), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OR3_X1    g0594(.A1(new_n792), .A2(KEYINPUT32), .A3(new_n793), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n309), .A2(G179), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n769), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n562), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n781), .A2(new_n777), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(G68), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n370), .A2(G179), .A3(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n207), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G97), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n801), .A2(new_n304), .A3(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n787), .A2(G179), .A3(new_n309), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G107), .B2(new_n807), .ZN(new_n808));
  AND4_X1   g0608(.A1(new_n786), .A2(new_n794), .A3(new_n795), .A4(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT33), .B(G317), .Z(new_n810));
  INV_X1    g0610(.A(G303), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n799), .B1(new_n797), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G326), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n782), .A2(new_n813), .B1(new_n778), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n495), .A2(new_n496), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(new_n637), .C2(new_n803), .ZN(new_n818));
  INV_X1    g0618(.A(new_n807), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  INV_X1    g0620(.A(G322), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n819), .A2(new_n820), .B1(new_n821), .B2(new_n776), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n792), .A2(KEYINPUT105), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n792), .A2(KEYINPUT105), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n818), .B(new_n822), .C1(new_n825), .C2(G329), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n768), .B1(new_n809), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(G13), .A2(G33), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(G20), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n229), .A2(G355), .A3(new_n304), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n230), .A2(new_n379), .ZN(new_n832));
  INV_X1    g0632(.A(new_n224), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n284), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n249), .A2(new_n486), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n831), .B1(G116), .B2(new_n229), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n830), .B(new_n768), .C1(new_n836), .C2(KEYINPUT99), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT99), .B2(new_n836), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n827), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n830), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n697), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n767), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n698), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n697), .A2(G330), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n766), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  NOR2_X1   g0647(.A1(new_n768), .A2(new_n828), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT106), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n766), .B1(new_n211), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n817), .B1(new_n451), .B2(new_n797), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT107), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n819), .A2(new_n562), .ZN(new_n854));
  INV_X1    g0654(.A(new_n778), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G283), .A2(new_n800), .B1(new_n855), .B2(G116), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n805), .C1(new_n811), .C2(new_n782), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n776), .A2(new_n637), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n853), .A2(new_n854), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n825), .A2(G311), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n825), .A2(G132), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G137), .A2(new_n783), .B1(new_n855), .B2(G159), .ZN(new_n862));
  INV_X1    g0662(.A(G150), .ZN(new_n863));
  INV_X1    g0663(.A(G143), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n863), .B2(new_n799), .C1(new_n776), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(KEYINPUT108), .B(KEYINPUT34), .Z(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n819), .A2(new_n335), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n379), .B1(new_n202), .B2(new_n797), .C1(new_n265), .C2(new_n803), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n859), .A2(new_n860), .B1(new_n861), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n768), .ZN(new_n873));
  AND4_X1   g0673(.A1(new_n459), .A2(new_n457), .A3(new_n455), .A4(new_n694), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n693), .B1(new_n441), .B2(new_n443), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n463), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n460), .B2(new_n876), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n851), .B1(new_n872), .B2(new_n873), .C1(new_n877), .C2(new_n829), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n755), .B(new_n877), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n767), .B1(new_n879), .B2(new_n741), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n879), .A2(new_n741), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(G384));
  OAI211_X1 g0683(.A(G116), .B(new_n226), .C1(new_n473), .C2(KEYINPUT35), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(KEYINPUT35), .B2(new_n473), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT36), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n224), .B(G77), .C1(new_n265), .C2(new_n335), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n202), .A2(G68), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n206), .B(G13), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  OR3_X1    g0690(.A1(new_n368), .A2(KEYINPUT110), .A3(new_n694), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n368), .B(new_n373), .C1(new_n369), .C2(new_n694), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT110), .B1(new_n368), .B2(new_n694), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n397), .B1(new_n413), .B2(new_n414), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n896), .A2(new_n409), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n415), .A2(new_n259), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n418), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n691), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n428), .B2(new_n436), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n416), .A2(new_n418), .A3(new_n394), .A4(new_n392), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n899), .B1(new_n433), .B2(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n425), .A2(new_n433), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n425), .A2(new_n900), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n903), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n895), .B1(new_n902), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n662), .A2(new_n663), .A3(new_n427), .A4(new_n419), .ZN(new_n913));
  INV_X1    g0713(.A(new_n901), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n906), .A2(new_n910), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n694), .B(new_n877), .C1(new_n676), .C2(new_n686), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT109), .ZN(new_n920));
  INV_X1    g0720(.A(new_n874), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n894), .B(new_n918), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT111), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n664), .A2(new_n691), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n902), .A2(new_n911), .A3(new_n895), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n915), .B2(new_n916), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT39), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  INV_X1    g0731(.A(new_n908), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n907), .A2(new_n908), .A3(new_n903), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n913), .A2(new_n932), .B1(new_n934), .B2(new_n910), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n917), .B(new_n931), .C1(new_n935), .C2(KEYINPUT38), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n368), .A2(new_n693), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT112), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n927), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n754), .A2(new_n465), .A3(new_n757), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n673), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n944), .B(new_n946), .Z(new_n947));
  AOI21_X1  g0747(.A(new_n694), .B1(new_n730), .B2(new_n734), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT31), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n739), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(new_n877), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n894), .A3(new_n918), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT40), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n917), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n951), .A2(KEYINPUT40), .A3(new_n894), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n950), .A2(new_n465), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n957), .B(new_n958), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(G330), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n947), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n206), .B2(new_n763), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n947), .A2(new_n960), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n890), .B1(new_n962), .B2(new_n963), .ZN(G367));
  INV_X1    g0764(.A(new_n832), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n244), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n830), .A2(new_n768), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n229), .B2(new_n437), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G294), .A2(new_n800), .B1(new_n855), .B2(G283), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n814), .B2(new_n782), .C1(new_n819), .C2(new_n353), .ZN(new_n970));
  INV_X1    g0770(.A(new_n776), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(G303), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n797), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n974), .A2(new_n975), .B1(new_n451), .B2(new_n803), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n379), .B(new_n976), .C1(new_n975), .C2(new_n974), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n972), .B(new_n977), .C1(new_n978), .C2(new_n792), .ZN(new_n979));
  INV_X1    g0779(.A(G137), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n792), .A2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n971), .A2(G150), .B1(new_n807), .B2(G77), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n265), .A2(new_n797), .B1(new_n799), .B2(new_n793), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n782), .A2(new_n864), .B1(new_n778), .B2(new_n202), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n803), .A2(new_n335), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n817), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n982), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n979), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT47), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n768), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n767), .B1(new_n966), .B2(new_n968), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT114), .Z(new_n994));
  INV_X1    g0794(.A(new_n679), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n563), .A2(new_n693), .ZN(new_n996));
  MUX2_X1   g0796(.A(new_n995), .B(new_n574), .S(new_n996), .Z(new_n997));
  OAI21_X1  g0797(.A(new_n994), .B1(new_n840), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n481), .B1(new_n681), .B2(new_n693), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n525), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n532), .B2(new_n694), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n609), .A2(new_n693), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(new_n702), .A3(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT42), .Z(new_n1004));
  OAI21_X1  g0804(.A(new_n532), .B1(new_n1000), .B2(new_n648), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n694), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT113), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n997), .B(KEYINPUT43), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n704), .A2(new_n1001), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n765), .A2(G1), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1001), .A2(new_n708), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT44), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n1001), .A2(new_n708), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT45), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n704), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n698), .A2(new_n703), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n705), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(new_n1002), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n760), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n760), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n710), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1015), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n998), .B1(new_n1014), .B2(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n1024), .A2(new_n1015), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n240), .A2(new_n284), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT115), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n262), .A2(G50), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  AOI211_X1 g0835(.A(G45), .B(new_n711), .C1(G68), .C2(G77), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n965), .B(new_n1033), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n229), .A2(new_n304), .A3(new_n711), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(G107), .B2(new_n229), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n967), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n792), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT116), .B(G150), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n803), .A2(new_n437), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n778), .A2(new_n335), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n797), .A2(new_n211), .ZN(new_n1046));
  NOR4_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n636), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n807), .A2(G97), .B1(new_n268), .B2(new_n800), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n782), .A2(KEYINPUT117), .A3(new_n793), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT117), .B1(new_n782), .B2(new_n793), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n971), .A2(G50), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1043), .A2(new_n1047), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n379), .B1(new_n807), .B2(G116), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n803), .A2(new_n820), .B1(new_n797), .B2(new_n637), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G322), .A2(new_n783), .B1(new_n855), .B2(G303), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n814), .B2(new_n799), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G317), .B2(new_n971), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1057), .B2(KEYINPUT48), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(KEYINPUT48), .B2(new_n1057), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT49), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1053), .B1(new_n813), .B2(new_n792), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1052), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n766), .B1(new_n1063), .B2(new_n768), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1040), .B(new_n1064), .C1(new_n702), .C2(new_n840), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1024), .A2(new_n760), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n710), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1024), .A2(new_n760), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1031), .B(new_n1065), .C1(new_n1067), .C2(new_n1068), .ZN(G393));
  XNOR2_X1  g0869(.A(new_n1020), .B(new_n705), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n1066), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1025), .A2(new_n710), .A3(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1001), .A2(new_n840), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n967), .B1(new_n229), .B2(new_n353), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n832), .B2(new_n252), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n817), .B1(new_n593), .B2(new_n803), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n973), .A2(G283), .B1(new_n800), .B2(G303), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n637), .B2(new_n778), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(G107), .C2(new_n807), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n792), .B2(new_n821), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n776), .A2(new_n814), .B1(new_n978), .B2(new_n782), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT52), .Z(new_n1084));
  AOI22_X1  g0884(.A1(new_n973), .A2(G68), .B1(new_n800), .B2(G50), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n262), .B2(new_n778), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n379), .B1(new_n211), .B2(new_n803), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n854), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n792), .B2(new_n864), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n776), .A2(new_n793), .B1(new_n863), .B2(new_n782), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT51), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n1082), .A2(new_n1084), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n766), .B(new_n1077), .C1(new_n1092), .C2(new_n768), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1021), .A2(new_n1015), .B1(new_n1075), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1073), .A2(new_n1074), .A3(new_n1094), .ZN(G390));
  OAI21_X1  g0895(.A(new_n767), .B1(new_n268), .B2(new_n849), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n825), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n637), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n869), .B1(G116), .B2(new_n971), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n799), .A2(new_n451), .B1(new_n778), .B2(new_n353), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n798), .B(new_n1100), .C1(G283), .C2(new_n783), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n304), .B1(G77), .B2(new_n804), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(G125), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n973), .A2(new_n1042), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G50), .B2(new_n807), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n782), .A2(new_n1109), .B1(new_n799), .B2(new_n980), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n817), .B(new_n1110), .C1(G159), .C2(new_n804), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT120), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n971), .A2(G132), .B1(new_n855), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1108), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1098), .A2(new_n1103), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1096), .B1(new_n1116), .B2(new_n768), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n937), .B2(new_n829), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT121), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n460), .A2(new_n876), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n753), .A2(new_n694), .A3(new_n1120), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1121), .A2(new_n921), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n894), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n939), .B(new_n955), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n919), .A2(new_n921), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT109), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n940), .B1(new_n1128), .B2(new_n894), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1124), .B1(new_n1129), .B2(new_n937), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n950), .A2(G330), .A3(new_n894), .A4(new_n877), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n739), .A2(new_n740), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(G330), .A3(new_n894), .A4(new_n877), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1124), .B(new_n1135), .C1(new_n1129), .C2(new_n937), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1015), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n950), .A2(G330), .A3(new_n465), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n673), .A2(new_n945), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n648), .A2(new_n652), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n608), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n657), .A2(new_n1142), .A3(new_n601), .A4(new_n606), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(new_n574), .A3(new_n749), .A4(new_n694), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n948), .B1(new_n1145), .B2(KEYINPUT31), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n949), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n877), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1123), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1122), .A2(new_n1149), .A3(new_n1135), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n740), .ZN(new_n1151));
  OAI211_X1 g0951(.A(G330), .B(new_n877), .C1(new_n1146), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1123), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1153), .A2(new_n1131), .B1(new_n1127), .B2(new_n1126), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1140), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1157), .B(new_n1140), .C1(new_n1150), .C2(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n710), .B1(new_n1137), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1153), .A2(new_n1131), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1128), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1122), .A2(new_n1149), .A3(new_n1135), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1157), .B1(new_n1164), .B2(new_n1140), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n673), .A2(new_n945), .A3(new_n1139), .ZN(new_n1166));
  AOI211_X1 g0966(.A(KEYINPUT119), .B(new_n1166), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1133), .B(new_n1136), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1119), .B(new_n1138), .C1(new_n1160), .C2(new_n1169), .ZN(G378));
  OAI211_X1 g0970(.A(new_n326), .B(new_n900), .C1(new_n661), .C2(new_n324), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n321), .B(new_n327), .C1(new_n325), .C2(new_n691), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n942), .B2(new_n943), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n954), .A2(G330), .A3(new_n956), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n924), .A2(new_n926), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT111), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1181), .A2(new_n927), .A3(new_n941), .A4(new_n1176), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1179), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1166), .B1(new_n1137), .B2(new_n1159), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT57), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1179), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1168), .A2(new_n1140), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1188), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n710), .B1(new_n1187), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1015), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n766), .B1(new_n202), .B2(new_n848), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G97), .A2(new_n800), .B1(new_n855), .B2(new_n438), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n593), .B2(new_n782), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G58), .B2(new_n807), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n986), .A2(new_n379), .A3(new_n1046), .A4(G41), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n451), .C2(new_n776), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n825), .B2(G283), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT58), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n288), .B1(new_n636), .B2(new_n287), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n202), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n971), .A2(G128), .B1(new_n973), .B2(new_n1113), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n804), .A2(G150), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n855), .A2(G137), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G125), .A2(new_n783), .B1(new_n800), .B2(G132), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1041), .A2(G124), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n807), .C2(G159), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1205), .A2(new_n1207), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(KEYINPUT58), .B2(new_n1204), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1198), .B1(new_n873), .B2(new_n1219), .C1(new_n1177), .C2(new_n829), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1197), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1196), .A2(new_n1222), .ZN(G375));
  XNOR2_X1  g1023(.A(new_n1015), .B(KEYINPUT122), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1123), .A2(new_n828), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n767), .B1(G68), .B2(new_n849), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1097), .A2(new_n811), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n782), .A2(new_n637), .B1(new_n799), .B2(new_n593), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n797), .A2(new_n353), .B1(new_n778), .B2(new_n451), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1044), .A4(new_n304), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n211), .B2(new_n819), .C1(new_n820), .C2(new_n776), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1097), .A2(new_n1109), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G132), .A2(new_n783), .B1(new_n855), .B2(G150), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n793), .B2(new_n797), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n636), .B(new_n1235), .C1(G50), .C2(new_n804), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n807), .A2(G58), .B1(new_n1113), .B2(new_n800), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n980), .C2(new_n776), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n1228), .A2(new_n1232), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1227), .B1(new_n1239), .B2(new_n768), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1164), .A2(new_n1225), .B1(new_n1226), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1164), .A2(new_n1140), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1028), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1241), .B1(new_n1244), .B2(new_n1159), .ZN(G381));
  INV_X1    g1045(.A(G378), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1196), .A2(new_n1246), .A3(new_n1222), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(G387), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(G390), .A2(G381), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(G407));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G343), .C2(new_n1247), .ZN(G409));
  NAND3_X1  g1052(.A1(new_n1156), .A2(KEYINPUT60), .A3(new_n1158), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1243), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n762), .B1(new_n1242), .B2(KEYINPUT60), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1254), .B1(new_n1253), .B2(new_n1243), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1241), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G384), .B(new_n1241), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1265));
  INV_X1    g1065(.A(G213), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(G343), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(G2897), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1264), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1225), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1220), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT123), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT123), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1274), .A2(new_n1277), .A3(new_n1220), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1191), .A2(new_n1192), .B1(new_n1168), .B2(new_n1140), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1028), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1246), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1196), .A2(G378), .A3(new_n1222), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1267), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT63), .B1(new_n1273), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1267), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1193), .A2(new_n1188), .A3(new_n1194), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n762), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1289), .A2(new_n1246), .A3(new_n1221), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1275), .A2(KEYINPUT123), .B1(new_n1028), .B2(new_n1279), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G378), .B1(new_n1291), .B2(new_n1278), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1286), .B(new_n1271), .C1(new_n1290), .C2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1285), .A2(new_n1293), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1073), .A2(new_n1074), .A3(new_n1094), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1013), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1012), .B(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1015), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(G390), .A2(new_n1302), .A3(new_n998), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1296), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(new_n846), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1296), .B(new_n1303), .C1(new_n1305), .C2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1293), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1314), .B2(KEYINPUT63), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1294), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1286), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1286), .A4(new_n1271), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1318), .A2(new_n1319), .A3(new_n1312), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1311), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1316), .A2(new_n1325), .ZN(G405));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1246), .B1(new_n1196), .B2(new_n1222), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1271), .B1(new_n1248), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1328), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1271), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1247), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1327), .B1(new_n1333), .B2(new_n1324), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1329), .A2(new_n1332), .A3(KEYINPUT127), .A4(new_n1311), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1324), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .ZN(G402));
endmodule


