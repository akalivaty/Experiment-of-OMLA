//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT68), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n455), .A2(G2106), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(G567), .B2(new_n458), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT70), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n468), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n473), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n467), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n476), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n475), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n472), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n471), .A2(new_n473), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(G2105), .A3(new_n468), .ZN(new_n492));
  OAI221_X1 g067(.A(new_n487), .B1(new_n488), .B2(new_n489), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT71), .ZN(G162));
  AND4_X1   g069(.A1(G138), .A2(new_n478), .A3(new_n473), .A4(new_n472), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  OAI22_X1  g071(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n474), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT72), .B(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(new_n472), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n468), .A2(new_n471), .A3(new_n473), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n497), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n510), .A2(KEYINPUT74), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n510), .A2(KEYINPUT74), .B1(G75), .B2(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n506), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G543), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n509), .A3(new_n520), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n514), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n513), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(new_n522), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  INV_X1    g102(.A(new_n521), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n509), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  XNOR2_X1  g111(.A(KEYINPUT75), .B(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n528), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n506), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n526), .A2(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n544), .A2(new_n521), .B1(new_n522), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  OAI221_X1 g123(.A(new_n548), .B1(new_n522), .B2(new_n545), .C1(new_n544), .C2(new_n521), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n506), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n550), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(G860), .A3(new_n556), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n519), .A2(G53), .A3(G543), .A4(new_n520), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n507), .B2(new_n508), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n507), .A2(new_n566), .A3(new_n508), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n526), .A2(G91), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n564), .A2(new_n573), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND2_X1  g151(.A1(new_n528), .A2(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n526), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n506), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n526), .A2(G86), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n517), .A2(new_n518), .B1(new_n516), .B2(G651), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  AND2_X1   g161(.A1(G48), .A2(G543), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n583), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n526), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n528), .A2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n506), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n526), .A2(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT10), .Z(new_n597));
  INV_X1    g172(.A(new_n569), .ZN(new_n598));
  OAI21_X1  g173(.A(G66), .B1(new_n598), .B2(new_n567), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n506), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(G54), .B2(new_n528), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G284));
  XNOR2_X1  g180(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  XNOR2_X1  g184(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n554), .A2(new_n556), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n603), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g192(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n618));
  XNOR2_X1  g193(.A(G323), .B(new_n618), .ZN(G282));
  NAND2_X1  g194(.A1(new_n475), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n472), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(new_n492), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(new_n624), .A3(G123), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n624), .B1(new_n623), .B2(G123), .ZN(new_n627));
  OAI221_X1 g202(.A(new_n620), .B1(new_n621), .B2(new_n622), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n630));
  NOR3_X1   g205(.A1(new_n470), .A2(new_n467), .A3(G2105), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2100), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n628), .A2(G2096), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(G156));
  INV_X1    g211(.A(G14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  AOI211_X1 g227(.A(new_n637), .B(new_n652), .C1(new_n650), .C2(new_n649), .ZN(G401));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT87), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT17), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n655), .B2(new_n657), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n656), .B2(new_n657), .ZN(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(new_n658), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2096), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  INV_X1    g251(.A(new_n671), .ZN(new_n677));
  INV_X1    g252(.A(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n680), .C1(new_n677), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G6), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G22), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G166), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n689), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n689), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n694), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT34), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n475), .A2(G131), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  INV_X1    g285(.A(G107), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G2105), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n623), .B2(G119), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n707), .B1(new_n715), .B2(new_n706), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT90), .Z(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(G290), .A2(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n689), .A2(G24), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1986), .Z(new_n726));
  NOR4_X1   g301(.A1(new_n705), .A2(new_n719), .A3(new_n720), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT36), .ZN(new_n728));
  INV_X1    g303(.A(G32), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G105), .B2(new_n483), .ZN(new_n734));
  INV_X1    g309(.A(G129), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n492), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n475), .A2(G141), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n730), .B1(new_n739), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT97), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n706), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n706), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT98), .Z(new_n746));
  OAI21_X1  g321(.A(new_n743), .B1(G2078), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G162), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G2090), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n706), .A2(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n475), .A2(G139), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g329(.A1(G115), .A2(G2104), .ZN(new_n755));
  INV_X1    g330(.A(G127), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n479), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n758));
  NAND2_X1  g333(.A1(G103), .A2(G2104), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G2105), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n757), .A2(G2105), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n752), .B1(new_n763), .B2(new_n706), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2072), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n689), .A2(G20), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT23), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n608), .B2(new_n689), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1956), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n747), .A2(new_n751), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n750), .A2(G2090), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT99), .Z(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  NOR2_X1   g348(.A1(G168), .A2(new_n689), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n689), .B2(G21), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n740), .A2(new_n741), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n773), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n689), .A2(G5), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G171), .B2(new_n689), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G28), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT30), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n782), .B2(KEYINPUT30), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n788), .B2(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(KEYINPUT24), .B2(new_n788), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n485), .B2(new_n706), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n628), .A2(new_n706), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n793), .B(new_n794), .C1(new_n792), .C2(new_n791), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n777), .A2(new_n781), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n689), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n604), .B2(new_n689), .ZN(new_n798));
  INV_X1    g373(.A(G1348), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n746), .A2(G2078), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n706), .A2(G26), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT28), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n475), .A2(G140), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT93), .B1(G104), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(KEYINPUT93), .A2(G104), .A3(G2105), .ZN(new_n808));
  OAI221_X1 g383(.A(G2104), .B1(G116), .B2(new_n472), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G128), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n805), .B(new_n809), .C1(new_n492), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT94), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n804), .B1(new_n812), .B2(G29), .ZN(new_n813));
  INV_X1    g388(.A(G2067), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n796), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G19), .B(new_n613), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1341), .Z(new_n818));
  NAND4_X1  g393(.A1(new_n770), .A2(new_n772), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n728), .A2(new_n819), .ZN(G150));
  XNOR2_X1  g395(.A(G150), .B(KEYINPUT100), .ZN(G311));
  NAND2_X1  g396(.A1(new_n526), .A2(G93), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n506), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n528), .A2(G55), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n554), .A2(new_n556), .A3(new_n826), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n550), .A2(new_n552), .ZN(new_n831));
  OAI21_X1  g406(.A(KEYINPUT102), .B1(new_n831), .B2(new_n826), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n826), .B1(new_n550), .B2(new_n552), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n833), .B(KEYINPUT102), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n839), .A2(KEYINPUT103), .A3(new_n830), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n604), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n829), .B1(new_n846), .B2(new_n848), .ZN(G145));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n763), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n739), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n714), .B(new_n632), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n496), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT4), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n478), .A2(new_n473), .A3(G138), .A4(new_n472), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n475), .A2(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n859));
  INV_X1    g434(.A(new_n503), .ZN(new_n860));
  INV_X1    g435(.A(G114), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT72), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT72), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G114), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n498), .B1(new_n865), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n859), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n501), .A2(KEYINPUT105), .A3(new_n503), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n858), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n812), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n623), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n472), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n475), .A2(KEYINPUT107), .A3(G142), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT107), .B1(new_n475), .B2(G142), .ZN(new_n875));
  OAI221_X1 g450(.A(new_n871), .B1(new_n872), .B2(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n870), .B(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n854), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(G162), .B(G160), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n628), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n854), .A2(new_n877), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT108), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n878), .A2(new_n881), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n883), .B(new_n884), .C1(new_n880), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g462(.A1(new_n826), .A2(new_n614), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n603), .A2(G299), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n597), .A2(new_n608), .A3(new_n602), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n891), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n891), .B(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n894), .B2(KEYINPUT109), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n841), .A2(new_n616), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n838), .B(new_n840), .C1(G559), .C2(new_n603), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n898), .B(KEYINPUT110), .C1(new_n899), .C2(new_n891), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n901), .A3(new_n895), .ZN(new_n902));
  XOR2_X1   g477(.A(G305), .B(G290), .Z(new_n903));
  XNOR2_X1  g478(.A(G166), .B(G288), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT42), .Z(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT112), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n900), .A2(KEYINPUT112), .A3(new_n902), .A4(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI211_X1 g486(.A(KEYINPUT111), .B(new_n906), .C1(new_n900), .C2(new_n902), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n906), .B1(new_n900), .B2(new_n902), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT111), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n888), .B1(new_n916), .B2(new_n614), .ZN(G295));
  OAI21_X1  g492(.A(new_n888), .B1(new_n916), .B2(new_n614), .ZN(G331));
  XNOR2_X1  g493(.A(G301), .B(G286), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n838), .A2(new_n840), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n891), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n838), .B2(new_n840), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(KEYINPUT113), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT113), .ZN(new_n926));
  AOI211_X1 g501(.A(new_n926), .B(new_n919), .C1(new_n838), .C2(new_n840), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n920), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n928), .B2(new_n895), .ZN(new_n929));
  AOI21_X1  g504(.A(G37), .B1(new_n929), .B2(new_n905), .ZN(new_n930));
  INV_X1    g505(.A(new_n905), .ZN(new_n931));
  INV_X1    g506(.A(new_n919), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n836), .A2(new_n837), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT103), .B1(new_n839), .B2(new_n830), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n926), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n923), .A2(KEYINPUT113), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n922), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n894), .B1(new_n935), .B2(new_n920), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n931), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT114), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(KEYINPUT114), .B(new_n931), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n930), .A2(KEYINPUT43), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(new_n924), .ZN(new_n946));
  INV_X1    g521(.A(new_n920), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n936), .B2(new_n937), .ZN(new_n948));
  INV_X1    g523(.A(new_n895), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n905), .B(new_n946), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n884), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n929), .A2(new_n905), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n944), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT44), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n930), .A2(new_n945), .A3(new_n942), .A4(new_n943), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n951), .B2(new_n952), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n960), .ZN(G397));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT45), .B1(new_n869), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n485), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n812), .B(G2067), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n967), .B2(new_n739), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT116), .Z(new_n971));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n966), .A2(new_n739), .A3(G1996), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT117), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n966), .B2(new_n967), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n971), .A2(new_n738), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n718), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n981), .A2(new_n982), .A3(new_n714), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n812), .A2(G2067), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n966), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n715), .B(new_n718), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n981), .B1(new_n966), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(G290), .A2(G1986), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n966), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n976), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n962), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT118), .B1(new_n869), .B2(new_n962), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT50), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n962), .B1(new_n497), .B2(new_n504), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n965), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1956), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT124), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT57), .B1(new_n564), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G299), .ZN(new_n1005));
  OAI21_X1  g580(.A(G65), .B1(new_n598), .B2(new_n567), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n571), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1007), .A2(G651), .B1(G91), .B2(new_n526), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n564), .C1(new_n1003), .C2(KEYINPUT57), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n869), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n996), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n965), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1002), .A2(new_n1011), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT125), .ZN(new_n1021));
  INV_X1    g596(.A(new_n965), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n993), .A2(new_n994), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n501), .A2(KEYINPUT105), .A3(new_n503), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT105), .B1(new_n501), .B2(new_n503), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n497), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(new_n1027), .B2(G1384), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n962), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n998), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n965), .A3(new_n1031), .ZN(new_n1032));
  AOI221_X4 g607(.A(new_n1021), .B1(new_n1023), .B2(new_n814), .C1(new_n1032), .C2(new_n799), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n799), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1023), .A2(new_n814), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT125), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1033), .A2(new_n1036), .A3(new_n603), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1011), .B1(new_n1002), .B2(new_n1019), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1020), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1021), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(KEYINPUT125), .A3(new_n1035), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT60), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n604), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT60), .B(new_n603), .C1(new_n1033), .C2(new_n1036), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT61), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1018), .B(new_n1010), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1038), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n999), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1956), .B1(new_n1053), .B2(new_n965), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1010), .B1(new_n1054), .B2(new_n1018), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(KEYINPUT61), .A3(new_n1020), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1015), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1028), .A2(new_n965), .A3(new_n1029), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT58), .B(G1341), .Z(new_n1059));
  AOI22_X1  g634(.A1(new_n969), .A2(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OR3_X1    g635(.A1(new_n1060), .A2(KEYINPUT59), .A3(new_n613), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT59), .B1(new_n1060), .B2(new_n613), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1047), .A2(new_n1050), .A3(new_n1056), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1039), .B1(new_n1046), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1032), .A2(new_n780), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1052), .A2(new_n1013), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G2078), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n965), .B1(new_n1013), .B2(new_n996), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1067), .A2(new_n1073), .A3(KEYINPUT126), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT126), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1069), .B1(new_n1015), .B2(G2078), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1012), .A2(new_n965), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n963), .A2(new_n1069), .A3(G2078), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1067), .B(new_n1077), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1066), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT45), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n773), .B1(new_n1084), .B2(new_n1071), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1030), .A2(new_n792), .A3(new_n965), .A4(new_n1031), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(G168), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(G168), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT51), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(KEYINPUT51), .B2(new_n1088), .ZN(new_n1091));
  OAI211_X1 g666(.A(G301), .B(new_n1077), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1066), .B1(new_n1081), .B2(G171), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1015), .A2(new_n697), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT119), .B(G2090), .Z(new_n1100));
  NOR2_X1   g675(.A1(new_n1022), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1099), .B1(new_n1053), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT122), .B1(G305), .B2(G1981), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT121), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n584), .B(new_n1108), .C1(new_n589), .C2(new_n588), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1109), .A3(new_n583), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1105), .B1(new_n1110), .B2(G1981), .ZN(new_n1111));
  INV_X1    g686(.A(G1981), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n582), .B1(new_n1106), .B2(KEYINPUT121), .ZN(new_n1113));
  AOI211_X1 g688(.A(KEYINPUT122), .B(new_n1112), .C1(new_n1113), .C2(new_n1109), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT49), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1023), .A2(new_n1103), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(new_n1117), .A3(G1981), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT49), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1112), .B1(new_n1113), .B2(new_n1109), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n1105), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n700), .A2(G1976), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1058), .A2(G8), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT52), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT120), .B(G1976), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT52), .B1(G288), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1058), .A2(G8), .A3(new_n1123), .A4(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1030), .A2(new_n1031), .A3(new_n1101), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1015), .A2(new_n697), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1103), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1098), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1104), .A2(new_n1122), .A3(new_n1129), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1091), .A2(new_n1094), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1065), .A2(new_n1083), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G288), .A2(G1976), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1122), .A2(new_n1140), .B1(new_n1112), .B2(new_n691), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1116), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1129), .A2(new_n1122), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n1134), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1103), .B(G286), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT123), .B1(new_n1135), .B2(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n995), .A2(new_n999), .A3(new_n1101), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1131), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1133), .B1(new_n1150), .B2(G8), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1129), .A2(new_n1122), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1145), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1147), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1143), .A2(new_n1146), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(KEYINPUT63), .A3(new_n1134), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1144), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1138), .A2(new_n1139), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1139), .B1(new_n1138), .B2(new_n1161), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1091), .A2(KEYINPUT62), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(new_n1078), .A3(new_n1136), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1091), .A2(KEYINPUT62), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1162), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n989), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT115), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n987), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n992), .B1(new_n1168), .B2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g748(.A1(G401), .A2(new_n465), .A3(G227), .A4(G229), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n958), .A2(new_n1175), .A3(new_n886), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


