//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n451, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  INV_X1    g025(.A(G567), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g029(.A1(G221), .A2(G218), .A3(G220), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT69), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2106), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n458), .A2(new_n451), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT71), .B(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G137), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n469), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n479), .ZN(G160));
  INV_X1    g055(.A(new_n468), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n469), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n482), .B1(new_n483), .B2(G136), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT72), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT73), .B1(new_n471), .B2(G114), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n489), .A2(new_n493), .A3(new_n492), .A4(KEYINPUT74), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n471), .A2(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n502), .B(new_n504), .C1(new_n475), .C2(new_n476), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n468), .A2(new_n469), .A3(G138), .A4(new_n499), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n498), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n517), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n518), .A2(G89), .ZN(new_n526));
  INV_X1    g101(.A(G63), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(new_n516), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n518), .A2(G543), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(new_n514), .B1(new_n529), .B2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT76), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n512), .A2(new_n513), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n516), .B1(new_n539), .B2(KEYINPUT77), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(KEYINPUT77), .B2(new_n539), .ZN(new_n541));
  INV_X1    g116(.A(new_n519), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G90), .B1(new_n529), .B2(G52), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n542), .A2(G81), .B1(new_n529), .B2(G43), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n516), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n537), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n542), .B2(G91), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n518), .A2(G53), .A3(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(new_n542), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n529), .A2(G49), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  NAND3_X1  g141(.A1(new_n514), .A2(new_n518), .A3(G86), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT79), .ZN(new_n568));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n512), .B2(new_n513), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT78), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n573), .B1(new_n570), .B2(KEYINPUT78), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(G48), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT80), .B1(new_n518), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(KEYINPUT6), .A2(G651), .ZN(new_n578));
  NOR2_X1   g153(.A1(KEYINPUT6), .A2(G651), .ZN(new_n579));
  OAI211_X1 g154(.A(KEYINPUT80), .B(new_n576), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n568), .A2(new_n575), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n529), .A2(G47), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT81), .B(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n519), .B2(new_n585), .C1(new_n516), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n519), .A2(KEYINPUT82), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT82), .B1(new_n519), .B2(new_n589), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT83), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n537), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n594), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n468), .A2(new_n472), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n483), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n469), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n482), .A2(G123), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n622), .A2(KEYINPUT84), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(KEYINPUT84), .ZN(new_n624));
  OAI221_X1 g199(.A(new_n619), .B1(new_n620), .B2(new_n621), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(G2100), .A2(new_n618), .B1(new_n625), .B2(G2096), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(G2096), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(G2100), .C2(new_n618), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n641), .A2(G14), .A3(new_n642), .ZN(G401));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NOR2_X1   g219(.A1(G2072), .A2(G2078), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n444), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n647), .B2(KEYINPUT85), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(KEYINPUT85), .B2(new_n647), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n646), .B(KEYINPUT17), .ZN(new_n652));
  INV_X1    g227(.A(new_n644), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n649), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n651), .A2(new_n646), .A3(new_n653), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n652), .A2(new_n653), .A3(new_n650), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  NOR2_X1   g252(.A1(G29), .A2(G35), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(G162), .B2(G29), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G2090), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT97), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n482), .A2(G129), .ZN(new_n685));
  NAND3_X1  g260(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT26), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT92), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G29), .B2(G32), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n691), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT27), .B(G1996), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT24), .ZN(new_n697));
  INV_X1    g272(.A(G34), .ZN(new_n698));
  AOI21_X1  g273(.A(G29), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G160), .B2(new_n689), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n696), .B1(G2084), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1961), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(G171), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G5), .B2(new_n704), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n702), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT94), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n689), .A2(G26), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n483), .A2(G140), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n482), .A2(G128), .ZN(new_n712));
  OAI221_X1 g287(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n710), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(G2067), .Z(new_n716));
  INV_X1    g291(.A(G1966), .ZN(new_n717));
  NOR2_X1   g292(.A1(G168), .A2(new_n704), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n704), .B2(G21), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n720), .B1(new_n717), .B2(new_n719), .C1(new_n695), .C2(new_n694), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n550), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G16), .B2(G19), .ZN(new_n723));
  INV_X1    g298(.A(G1341), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n625), .A2(new_n689), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G28), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n689), .B1(new_n727), .B2(G28), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT31), .B(G11), .Z(new_n733));
  NOR4_X1   g308(.A1(new_n725), .A2(new_n726), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n723), .A2(new_n724), .B1(G2084), .B2(new_n701), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(new_n703), .C2(new_n706), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n704), .A2(G20), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT23), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n606), .B2(new_n704), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1956), .Z(new_n740));
  NAND2_X1  g315(.A1(G164), .A2(G29), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G27), .B2(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(new_n443), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n443), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n721), .A2(new_n736), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n683), .A2(new_n708), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n681), .A2(G2090), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n689), .A2(G33), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n483), .A2(G139), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n753), .B(new_n754), .C1(new_n469), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT90), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(new_n689), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G2072), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT91), .Z(new_n761));
  NOR2_X1   g336(.A1(new_n602), .A2(new_n704), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G4), .B2(new_n704), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G2072), .B2(new_n759), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n764), .B2(new_n763), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n747), .A2(new_n749), .A3(new_n761), .A4(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G6), .B(G305), .S(G16), .Z(new_n769));
  XOR2_X1   g344(.A(KEYINPUT32), .B(G1981), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n704), .A2(G22), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G166), .B2(new_n704), .ZN(new_n776));
  INV_X1    g351(.A(G1971), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n704), .A2(G23), .ZN(new_n779));
  INV_X1    g354(.A(G288), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n704), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n773), .A2(new_n774), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT34), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n689), .A2(G25), .ZN(new_n787));
  AOI22_X1  g362(.A1(G119), .A2(new_n482), .B1(new_n483), .B2(G131), .ZN(new_n788));
  OAI221_X1 g363(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n787), .B1(new_n791), .B2(new_n689), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT86), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n798));
  MUX2_X1   g373(.A(G24), .B(G290), .S(G16), .Z(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G1986), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G1986), .B2(new_n799), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n796), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n785), .A2(new_n786), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(KEYINPUT89), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n768), .A2(new_n805), .A3(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  AOI22_X1  g383(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(new_n516), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  INV_X1    g386(.A(G55), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n519), .A2(new_n811), .B1(new_n521), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(new_n550), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n814), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(new_n549), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n601), .A2(new_n609), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(G860), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g401(.A(G860), .B1(new_n810), .B2(new_n813), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  XNOR2_X1  g404(.A(new_n790), .B(new_n616), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n757), .A2(new_n688), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n757), .A2(new_n688), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n833), .ZN(new_n835));
  INV_X1    g410(.A(new_n830), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n510), .B(new_n714), .ZN(new_n839));
  AOI22_X1  g414(.A1(G130), .A2(new_n482), .B1(new_n483), .B2(G142), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT99), .B1(new_n469), .B2(G118), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n469), .A2(KEYINPUT99), .A3(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n839), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n838), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n625), .B(G160), .Z(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(G162), .Z(new_n849));
  NAND3_X1  g424(.A1(new_n834), .A2(new_n837), .A3(new_n845), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n849), .B1(new_n847), .B2(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT100), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n856), .A2(new_n857), .A3(new_n852), .A4(new_n851), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g435(.A1(new_n602), .A2(new_n606), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n601), .A2(G299), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT41), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n866), .A2(KEYINPUT101), .A3(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n820), .B(new_n611), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n863), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT42), .ZN(new_n875));
  XNOR2_X1  g450(.A(G305), .B(G290), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n780), .B(G303), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(KEYINPUT42), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n875), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n875), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n814), .A2(G868), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(G295));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n885), .ZN(G331));
  XNOR2_X1  g462(.A(G301), .B(G286), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n820), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n816), .A2(new_n819), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n888), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(KEYINPUT103), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n894), .A3(new_n888), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n866), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n865), .A2(new_n867), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(KEYINPUT104), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n891), .A2(new_n900), .A3(new_n888), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n890), .A3(new_n901), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n893), .A2(new_n895), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT105), .B1(new_n904), .B2(new_n866), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n879), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n868), .A2(new_n893), .A3(new_n869), .A4(new_n895), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n899), .A2(new_n863), .A3(new_n890), .A4(new_n901), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n879), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n852), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n909), .A2(new_n852), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n908), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n878), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT43), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT44), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n906), .A2(new_n910), .A3(KEYINPUT43), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n920), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g496(.A(new_n714), .B(G2067), .Z(new_n922));
  INV_X1    g497(.A(G1996), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n688), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n790), .B(new_n795), .Z(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G290), .A2(G1986), .ZN(new_n929));
  AND2_X1   g504(.A1(G290), .A2(G1986), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n496), .A2(new_n497), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n479), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT106), .B(G40), .Z(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n938), .A2(new_n473), .A3(new_n470), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n931), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(G288), .A2(G1976), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n474), .A2(new_n479), .A3(new_n939), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n510), .A2(new_n932), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(G8), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n567), .B1(new_n577), .B2(new_n581), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT108), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(new_n567), .C1(new_n577), .C2(new_n581), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n575), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G1981), .ZN(new_n953));
  INV_X1    g528(.A(G1981), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n568), .A2(new_n575), .A3(new_n954), .A4(new_n582), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(KEYINPUT49), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT49), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n947), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n944), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n955), .B(KEYINPUT110), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n780), .A2(G1976), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n946), .A3(G8), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT52), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(G288), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n964), .A2(new_n946), .A3(new_n968), .A4(G8), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n959), .B2(new_n960), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n974));
  NOR2_X1   g549(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n933), .B2(new_n934), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n945), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n510), .B2(new_n932), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n977), .A2(new_n979), .A3(G2090), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n936), .A2(G1384), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n941), .B1(new_n510), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G1971), .B1(new_n937), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n974), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT55), .Z(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n933), .B2(new_n934), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n945), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n510), .B2(new_n932), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n777), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n935), .A2(KEYINPUT50), .ZN(new_n991));
  INV_X1    g566(.A(G2090), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n941), .B1(new_n510), .B2(new_n975), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(KEYINPUT107), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n984), .A2(G8), .A3(new_n986), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n963), .A2(new_n947), .B1(new_n973), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(G8), .B1(new_n980), .B2(new_n983), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n985), .B(KEYINPUT55), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n972), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n971), .B(KEYINPUT111), .C1(new_n959), .C2(new_n960), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n937), .A2(new_n443), .A3(new_n982), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT121), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(KEYINPUT121), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(KEYINPUT53), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n991), .A2(new_n993), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT122), .B(G1961), .Z(new_n1012));
  AOI22_X1  g587(.A1(new_n1006), .A2(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G301), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n717), .B1(new_n988), .B2(new_n989), .ZN(new_n1016));
  INV_X1    g591(.A(G2084), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n991), .A2(new_n1017), .A3(new_n993), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(G168), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n1020));
  AND2_X1   g595(.A1(KEYINPUT119), .A2(G8), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(G8), .A3(G286), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1020), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT62), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT51), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT62), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n1024), .A4(new_n1022), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n998), .B1(new_n1015), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT117), .B(KEYINPUT61), .Z(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT113), .B(G1956), .Z(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n977), .B2(new_n979), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n1037));
  XNOR2_X1  g612(.A(G299), .B(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(new_n442), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n937), .A2(new_n982), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1036), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1034), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT118), .B(new_n1034), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n937), .A2(new_n923), .A3(new_n982), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT58), .B(G1341), .Z(new_n1051));
  NAND2_X1  g626(.A1(new_n946), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n550), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT59), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1056), .A3(new_n550), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1049), .A2(KEYINPUT61), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n764), .B1(new_n977), .B2(new_n979), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n946), .A2(G2067), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT60), .B(new_n601), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT60), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1348), .B1(new_n991), .B2(new_n993), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n946), .A2(G2067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT115), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n602), .A3(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1048), .A2(new_n1058), .A3(new_n1065), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1062), .A3(new_n602), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1043), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1042), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n474), .A2(KEYINPUT123), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n470), .A2(new_n1082), .A3(new_n473), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1081), .A2(G40), .A3(new_n938), .A4(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT124), .B1(new_n989), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n937), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1010), .B(G2078), .C1(new_n510), .C2(new_n981), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1013), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1008), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT53), .B1(new_n1006), .B2(KEYINPUT121), .ZN(new_n1094));
  OAI211_X1 g669(.A(G301), .B(new_n1013), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(KEYINPUT54), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1029), .A2(new_n1024), .A3(new_n1022), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n1099));
  OAI21_X1  g674(.A(new_n1013), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1013), .A2(G301), .A3(new_n1090), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1080), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1033), .B1(new_n1079), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT112), .B(KEYINPUT63), .Z(new_n1106));
  INV_X1    g681(.A(G8), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1107), .B(G286), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1106), .B1(new_n1080), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n984), .A2(G8), .A3(new_n995), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1000), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1108), .A2(KEYINPUT63), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n973), .A2(new_n1112), .A3(new_n996), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n943), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n942), .A2(new_n923), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT46), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT126), .Z(new_n1120));
  INV_X1    g695(.A(new_n688), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n922), .A2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n942), .A2(new_n1122), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT47), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n942), .A2(new_n929), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n928), .A2(new_n942), .B1(KEYINPUT48), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1127), .A2(KEYINPUT48), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n791), .A2(new_n795), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT125), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1131), .A2(new_n925), .B1(G2067), .B2(new_n714), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1128), .A2(new_n1129), .B1(new_n942), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT127), .B1(new_n1116), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1079), .A2(new_n1104), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1033), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1115), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n943), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1134), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1135), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g719(.A1(G229), .A2(new_n466), .A3(G401), .A4(G227), .ZN(new_n1146));
  NAND2_X1  g720(.A1(new_n859), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n1147), .ZN(G308));
  OR2_X1    g722(.A1(new_n920), .A2(new_n1147), .ZN(G225));
endmodule


