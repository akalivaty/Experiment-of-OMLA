//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(G183gat), .B2(G190gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n213), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n223), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n222), .B(KEYINPUT65), .C1(new_n226), .C2(new_n227), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n219), .B1(new_n233), .B2(new_n218), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n237), .A2(KEYINPUT28), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n237), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n210), .A2(KEYINPUT66), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT66), .B1(new_n210), .B2(new_n241), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n212), .B(new_n240), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n238), .A2(new_n239), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n234), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  INV_X1    g046(.A(G113gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G120gat), .ZN(new_n249));
  INV_X1    g048(.A(G120gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(G113gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G134gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G127gat), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G134gat), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT67), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n254), .B2(new_n256), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n252), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT68), .B1(new_n250), .B2(G113gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(new_n248), .A3(G120gat), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n260), .B(new_n262), .C1(new_n248), .C2(G120gat), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n254), .A2(new_n256), .A3(new_n247), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n238), .A2(new_n239), .A3(new_n244), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n213), .B1(new_n228), .B2(new_n229), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT25), .B1(new_n269), .B2(new_n231), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n267), .B(new_n268), .C1(new_n270), .C2(new_n219), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n246), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n268), .B1(new_n270), .B2(new_n219), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n256), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(new_n252), .B1(new_n263), .B2(new_n264), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n273), .A2(KEYINPUT69), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n204), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n204), .B(new_n282), .C1(new_n272), .C2(new_n280), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n272), .A2(new_n204), .A3(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT70), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n291), .A3(KEYINPUT32), .ZN(new_n292));
  XNOR2_X1  g091(.A(G15gat), .B(G43gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G71gat), .B(G99gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n290), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT33), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n288), .A2(KEYINPUT32), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n288), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n287), .B1(new_n298), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n292), .A3(new_n297), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n286), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n307), .A2(KEYINPUT36), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT36), .B1(new_n307), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G155gat), .B(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n320), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(new_n266), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n323), .B2(new_n324), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n320), .A2(new_n322), .ZN(new_n333));
  INV_X1    g132(.A(new_n321), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n337), .A3(new_n266), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT75), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n332), .A2(new_n337), .A3(new_n340), .A4(new_n266), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n325), .B2(new_n266), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n335), .A2(new_n336), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n279), .A2(new_n345), .A3(KEYINPUT4), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND4_X1   g149(.A1(new_n327), .A2(new_n342), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n347), .B1(new_n339), .B2(new_n341), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n352), .B2(new_n327), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n330), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n359), .B(new_n330), .C1(new_n351), .C2(new_n353), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n342), .A2(new_n348), .A3(new_n327), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n349), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n352), .A2(new_n327), .A3(new_n350), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n359), .A4(new_n330), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(KEYINPUT22), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G226gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(new_n203), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n273), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n223), .A2(new_n225), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT64), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n216), .A2(new_n224), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n215), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n232), .B1(new_n384), .B2(KEYINPUT65), .ZN(new_n385));
  INV_X1    g184(.A(new_n231), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n218), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n219), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n245), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n378), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n376), .B1(new_n380), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n374), .B(new_n375), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n273), .A2(new_n378), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  NAND4_X1  g199(.A1(new_n392), .A2(new_n396), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n380), .A2(new_n391), .A3(new_n376), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n394), .B1(new_n393), .B2(new_n395), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n392), .A2(new_n396), .A3(new_n400), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n364), .A2(new_n369), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n376), .A2(KEYINPUT29), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n331), .B1(new_n409), .B2(KEYINPUT78), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n394), .A2(KEYINPUT78), .A3(new_n379), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n325), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n394), .B1(new_n379), .B2(new_n332), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(G228gat), .B2(G233gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n379), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n345), .B1(new_n416), .B2(new_n331), .ZN(new_n417));
  OAI211_X1 g216(.A(G228gat), .B(G233gat), .C1(new_n417), .C2(new_n413), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n415), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n415), .B2(new_n418), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G22gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OR3_X1    g224(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n421), .B2(new_n422), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n408), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n327), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n326), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n432), .A2(KEYINPUT39), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n342), .A2(new_n348), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n431), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n352), .A2(KEYINPUT39), .A3(new_n327), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(new_n438), .A3(new_n359), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT39), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(new_n440), .A3(new_n431), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT79), .B1(new_n441), .B2(new_n360), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT40), .B(new_n436), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n363), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n438), .B1(new_n437), .B2(new_n359), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT79), .A3(new_n360), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT40), .B1(new_n447), .B2(new_n436), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n407), .A2(new_n401), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n428), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT37), .B1(new_n403), .B2(new_n404), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT37), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n392), .A2(new_n396), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n402), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT38), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT38), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n453), .A2(new_n458), .A3(new_n402), .A4(new_n455), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n457), .A2(new_n406), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n363), .A2(new_n362), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n359), .B1(new_n368), .B2(new_n330), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n369), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT80), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT80), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n369), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n460), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n430), .B1(new_n452), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT81), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n286), .B1(new_n308), .B2(new_n309), .ZN(new_n470));
  AND4_X1   g269(.A1(new_n309), .A2(new_n304), .A3(new_n305), .A4(new_n286), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT35), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n450), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n464), .B2(new_n466), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT81), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n472), .A2(new_n475), .A3(new_n429), .A4(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n429), .B(new_n408), .C1(new_n470), .C2(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n313), .A2(new_n468), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n481), .A2(G1gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n484), .B2(G1gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n486), .A3(G8gat), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n482), .B(new_n485), .C1(KEYINPUT82), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n492));
  INV_X1    g291(.A(G29gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n495));
  AOI21_X1  g294(.A(G36gat), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n492), .A2(new_n497), .A3(G29gat), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n496), .A2(KEYINPUT15), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT15), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n500), .A2(new_n501), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n491), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n502), .A2(new_n503), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT18), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G113gat), .B(G141gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(G197gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT11), .B(G169gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(KEYINPUT12), .Z(new_n518));
  NAND4_X1  g317(.A1(new_n507), .A2(KEYINPUT18), .A3(new_n508), .A4(new_n510), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n490), .B(new_n509), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(new_n508), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n513), .A2(new_n518), .A3(new_n519), .A4(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n511), .A2(new_n512), .B1(new_n520), .B2(new_n523), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(KEYINPUT84), .A3(new_n518), .A4(new_n519), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n519), .ZN(new_n531));
  INV_X1    g330(.A(new_n518), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n480), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G183gat), .B(G211gat), .Z(new_n537));
  OR2_X1    g336(.A1(G57gat), .A2(G64gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(G57gat), .A2(G64gat), .ZN(new_n539));
  AND2_X1   g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(KEYINPUT9), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT85), .B1(G71gat), .B2(G78gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT21), .ZN(new_n550));
  INV_X1    g349(.A(G231gat), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n203), .ZN(new_n552));
  XNOR2_X1  g351(.A(G127gat), .B(G155gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT86), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(G231gat), .B(G233gat), .C1(new_n548), .C2(KEYINPUT21), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n552), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n537), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  INV_X1    g360(.A(new_n537), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n557), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n490), .B1(KEYINPUT21), .B2(new_n548), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n560), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n566), .B1(new_n560), .B2(new_n563), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  INV_X1    g373(.A(G85gat), .ZN(new_n575));
  INV_X1    g374(.A(G92gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(KEYINPUT8), .A2(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT8), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(G99gat), .B2(G106gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n581), .A2(KEYINPUT87), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n573), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G99gat), .B(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT88), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(KEYINPUT90), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT87), .B1(new_n581), .B2(new_n582), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n577), .A2(new_n578), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n572), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n585), .B(KEYINPUT88), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT89), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT89), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n598), .A3(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n595), .B2(new_n600), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n603), .A2(new_n604), .B1(new_n506), .B2(new_n505), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n595), .A2(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT91), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(new_n509), .A3(new_n602), .ZN(new_n608));
  AND2_X1   g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G190gat), .B(G218gat), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n612), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n605), .A2(new_n617), .A3(new_n608), .A4(new_n610), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n616), .B1(new_n613), .B2(new_n618), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n569), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n569), .B(KEYINPUT92), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT94), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n549), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n607), .A2(new_n602), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n631), .A2(KEYINPUT93), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n584), .A2(new_n587), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n548), .A2(new_n596), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n606), .B2(new_n549), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n629), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT93), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n607), .A2(new_n637), .A3(new_n602), .A4(new_n630), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n628), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n635), .A2(new_n628), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT95), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  AND3_X1   g444(.A1(new_n640), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n640), .B2(new_n642), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n625), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n536), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n463), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT96), .B(G1gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1324gat));
  AND2_X1   g453(.A1(new_n536), .A2(new_n650), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT97), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G8gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n451), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(G8gat), .B1(new_n651), .B2(new_n450), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n660), .A2(new_n662), .A3(KEYINPUT98), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT98), .B1(new_n660), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n311), .B2(new_n312), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT36), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n470), .B2(new_n471), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT36), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(KEYINPUT99), .A3(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(G15gat), .B1(new_n651), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n472), .A2(new_n476), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n480), .A2(new_n674), .A3(new_n535), .ZN(new_n675));
  INV_X1    g474(.A(G15gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n650), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n651), .A2(new_n429), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT43), .B(G22gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n452), .A2(new_n467), .ZN(new_n682));
  INV_X1    g481(.A(new_n430), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n313), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n477), .A2(new_n479), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n613), .A2(new_n618), .ZN(new_n687));
  INV_X1    g486(.A(new_n616), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n649), .A2(new_n535), .A3(new_n569), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n686), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n463), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n493), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n468), .A2(new_n667), .A3(new_n671), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n685), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n692), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n480), .B2(new_n691), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n693), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n463), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n697), .A2(new_n705), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n694), .A2(new_n497), .A3(new_n451), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT101), .B(KEYINPUT46), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G36gat), .B1(new_n704), .B2(new_n450), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1329gat));
  NOR4_X1   g510(.A1(new_n649), .A2(G43gat), .A3(new_n569), .A4(new_n691), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n675), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n704), .A2(new_n672), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n715));
  OAI21_X1  g514(.A(G43gat), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n704), .A2(KEYINPUT103), .A3(new_n672), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT47), .B(new_n713), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n719));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n675), .A2(new_n712), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(G1330gat));
  INV_X1    g523(.A(new_n700), .ZN(new_n725));
  AOI211_X1 g524(.A(new_n691), .B(new_n725), .C1(new_n698), .C2(new_n685), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n686), .B2(new_n692), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n428), .B(new_n693), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n703), .A2(KEYINPUT104), .A3(new_n428), .A4(new_n693), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(G50gat), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n429), .A2(G50gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n694), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT48), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n729), .A2(G50gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n735), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(G50gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n729), .B2(new_n730), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n736), .B1(new_n746), .B2(new_n732), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT48), .B1(new_n739), .B2(new_n735), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT105), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n749), .ZN(G1331gat));
  NAND4_X1  g549(.A1(new_n649), .A2(new_n623), .A3(new_n535), .A4(new_n624), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT106), .B1(new_n699), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n754), .B(new_n751), .C1(new_n698), .C2(new_n685), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n695), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n699), .A2(new_n752), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n754), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n699), .A2(KEYINPUT106), .A3(new_n752), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(KEYINPUT107), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n753), .B2(new_n755), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n450), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT108), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n762), .A2(new_n764), .A3(new_n768), .A4(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771));
  INV_X1    g570(.A(G64gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n767), .A2(new_n771), .A3(new_n772), .A4(new_n769), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1333gat));
  INV_X1    g575(.A(new_n672), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n764), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G71gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n674), .A2(G71gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n756), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n779), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(G1334gat));
  NAND3_X1  g584(.A1(new_n762), .A2(new_n764), .A3(new_n428), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT109), .B(G78gat), .Z(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1335gat));
  INV_X1    g587(.A(new_n569), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n535), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT110), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n648), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n703), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT111), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n703), .A2(new_n795), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797), .B2(new_n463), .ZN(new_n798));
  INV_X1    g597(.A(new_n791), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n699), .A2(new_n692), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n692), .A4(new_n799), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n648), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n575), .A3(new_n695), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n805), .ZN(G1336gat));
  OAI21_X1  g605(.A(G92gat), .B1(new_n793), .B2(new_n450), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n450), .A2(G92gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n451), .A3(new_n796), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n812), .A2(G92gat), .B1(new_n804), .B2(new_n808), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n810), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n797), .B2(new_n672), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n674), .A2(G99gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n804), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1338gat));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n648), .A2(new_n429), .A3(G106gat), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT112), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n794), .A2(new_n428), .A3(new_n796), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(G106gat), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  OAI21_X1  g624(.A(G106gat), .B1(new_n793), .B2(new_n429), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT53), .B1(new_n819), .B2(new_n821), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n826), .B2(new_n827), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n824), .A2(new_n825), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  NAND2_X1  g630(.A1(new_n631), .A2(KEYINPUT93), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(new_n627), .A3(new_n636), .A4(new_n638), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n640), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n645), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n628), .C1(new_n632), .C2(new_n639), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n837), .A2(new_n835), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT55), .A4(new_n834), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n534), .B1(new_n619), .B2(new_n620), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n507), .A2(new_n510), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(G229gat), .A3(G233gat), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n520), .A2(new_n523), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n517), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n527), .B2(new_n529), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n689), .B(new_n690), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n840), .B2(new_n834), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n646), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n843), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n649), .A2(new_n691), .A3(new_n849), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n569), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n623), .A2(new_n648), .A3(new_n535), .A4(new_n624), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n428), .A3(new_n674), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n451), .A2(new_n463), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n248), .A3(new_n535), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n861), .A2(new_n463), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n428), .B1(new_n307), .B2(new_n310), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n450), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n534), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n865), .B1(new_n872), .B2(new_n248), .ZN(G1340gat));
  NOR3_X1   g672(.A1(new_n864), .A2(new_n250), .A3(new_n648), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n649), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n250), .ZN(G1341gat));
  OAI21_X1  g675(.A(G127gat), .B1(new_n864), .B2(new_n789), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n789), .A2(G127gat), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n870), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT116), .ZN(G1342gat));
  NOR2_X1   g680(.A1(new_n691), .A2(new_n451), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n869), .A2(new_n253), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n864), .B2(new_n691), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G1343gat));
  NAND2_X1  g686(.A1(new_n672), .A2(new_n863), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n428), .C1(new_n858), .C2(new_n860), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n861), .B2(new_n429), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n892), .B(new_n894), .C1(new_n861), .C2(new_n429), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n316), .B1(new_n898), .B2(new_n534), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n777), .A2(new_n429), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n866), .A2(new_n900), .ZN(new_n901));
  NOR4_X1   g700(.A1(new_n901), .A2(G141gat), .A3(new_n451), .A4(new_n535), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT58), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n902), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n535), .B(new_n890), .C1(new_n896), .C2(new_n897), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n316), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(G1344gat));
  NOR3_X1   g707(.A1(new_n901), .A2(new_n451), .A3(new_n648), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n317), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n897), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n890), .A2(new_n648), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n856), .A2(new_n857), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n789), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n859), .B(KEYINPUT119), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n429), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n919), .B2(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n859), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n428), .B1(new_n922), .B2(new_n858), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(KEYINPUT120), .A3(new_n894), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n891), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n913), .ZN(new_n926));
  NAND2_X1  g725(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n911), .B(new_n914), .C1(new_n926), .C2(new_n927), .ZN(G1345gat));
  INV_X1    g727(.A(G155gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n898), .B2(new_n569), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n901), .A2(G155gat), .A3(new_n451), .A4(new_n789), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT121), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n931), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n789), .B(new_n890), .C1(new_n896), .C2(new_n897), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n933), .B(new_n934), .C1(new_n935), .C2(new_n929), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n936), .ZN(G1346gat));
  AND2_X1   g736(.A1(new_n898), .A2(new_n692), .ZN(new_n938));
  INV_X1    g737(.A(G162gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n882), .A2(new_n939), .ZN(new_n940));
  OAI22_X1  g739(.A1(new_n938), .A2(new_n939), .B1(new_n901), .B2(new_n940), .ZN(G1347gat));
  NAND2_X1  g740(.A1(new_n917), .A2(new_n859), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n867), .A2(new_n451), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n463), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n534), .A2(new_n205), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n944), .A2(KEYINPUT122), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT122), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n451), .A2(new_n463), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT123), .Z(new_n950));
  NAND2_X1  g749(.A1(new_n862), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n535), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n948), .A2(KEYINPUT124), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1348gat));
  OAI21_X1  g756(.A(G176gat), .B1(new_n951), .B2(new_n648), .ZN(new_n958));
  INV_X1    g757(.A(new_n944), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n206), .A3(new_n649), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1349gat));
  OAI21_X1  g760(.A(G183gat), .B1(new_n951), .B2(new_n789), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n235), .A3(new_n569), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n951), .B2(new_n691), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT125), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n968), .B(G190gat), .C1(new_n951), .C2(new_n691), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n967), .A2(KEYINPUT61), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n236), .A3(new_n692), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n970), .B(new_n971), .C1(KEYINPUT61), .C2(new_n967), .ZN(G1351gat));
  AND4_X1   g771(.A1(new_n463), .A2(new_n942), .A3(new_n451), .A4(new_n900), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n534), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n672), .A2(new_n950), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n925), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n534), .A2(G197gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(G1352gat));
  XOR2_X1   g779(.A(KEYINPUT127), .B(G204gat), .Z(new_n981));
  NAND3_X1  g780(.A1(new_n973), .A2(new_n649), .A3(new_n981), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n977), .A2(new_n648), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n983), .B(new_n984), .C1(new_n985), .C2(new_n981), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n973), .A2(new_n371), .A3(new_n569), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n925), .A2(new_n569), .A3(new_n976), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  OAI21_X1  g790(.A(G218gat), .B1(new_n977), .B2(new_n691), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n973), .A2(new_n372), .A3(new_n692), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1355gat));
endmodule


