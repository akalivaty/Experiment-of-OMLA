//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  XOR2_X1   g000(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .A4(G128), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n201), .A2(G128), .B1(new_n195), .B2(new_n197), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n193), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT65), .A2(G137), .ZN(new_n207));
  AOI21_X1  g021(.A(G134), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n198), .B1(G143), .B2(new_n194), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n196), .A2(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n194), .A2(G143), .ZN(new_n215));
  OAI22_X1  g029(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT67), .A3(new_n199), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT11), .A2(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n206), .A2(new_n207), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT11), .A2(G134), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT11), .A2(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G137), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n203), .A2(new_n211), .A3(new_n217), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G116), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G119), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n227), .B(new_n229), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n229), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n195), .A2(new_n197), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n240), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n246), .A2(new_n195), .A3(new_n197), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n219), .A2(new_n222), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n219), .B2(new_n222), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n245), .B(new_n248), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n225), .A2(new_n238), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n253), .A2(KEYINPUT70), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT70), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n216), .A2(new_n199), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n211), .A3(new_n224), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n238), .B1(new_n252), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n253), .B1(new_n260), .B2(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n252), .A2(new_n259), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n262), .A2(KEYINPUT69), .A3(new_n237), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT28), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n192), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n225), .A2(new_n238), .A3(new_n252), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n238), .B1(new_n225), .B2(new_n252), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n257), .B1(new_n269), .B2(new_n254), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(KEYINPUT29), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G902), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n225), .A2(KEYINPUT30), .A3(new_n252), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n237), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n253), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(new_n192), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n272), .B1(new_n279), .B2(KEYINPUT29), .ZN(new_n280));
  OAI21_X1  g094(.A(G472), .B1(new_n271), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n253), .A3(new_n192), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n285));
  INV_X1    g099(.A(new_n192), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n265), .B2(new_n286), .ZN(new_n287));
  AOI211_X1 g101(.A(KEYINPUT71), .B(new_n192), .C1(new_n257), .C2(new_n264), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n281), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G475), .A2(G902), .ZN(new_n295));
  INV_X1    g109(.A(G237), .ZN(new_n296));
  INV_X1    g110(.A(G953), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G214), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G143), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT83), .B(G143), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n301), .B(new_n223), .C1(new_n298), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT84), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n301), .B1(new_n302), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G131), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n299), .A2(G143), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n196), .A2(KEYINPUT83), .ZN(new_n308));
  OAI211_X1 g122(.A(G214), .B(new_n188), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT84), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n223), .A4(new_n301), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT17), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n304), .A2(new_n306), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT72), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n314), .A2(KEYINPUT72), .A3(G125), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT16), .B1(new_n314), .B2(G125), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n194), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n194), .B1(new_n320), .B2(new_n322), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n305), .A2(KEYINPUT17), .A3(G131), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n313), .A2(new_n323), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT18), .A2(G131), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n305), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G146), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n314), .A2(KEYINPUT72), .A3(G125), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n330), .B2(KEYINPUT72), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n334), .A2(G146), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n329), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(G113), .B(G122), .Z(new_n337));
  XOR2_X1   g151(.A(KEYINPUT85), .B(G104), .Z(new_n338));
  XOR2_X1   g152(.A(new_n337), .B(new_n338), .Z(new_n339));
  AND3_X1   g153(.A1(new_n327), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n321), .B1(new_n334), .B2(KEYINPUT16), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT74), .B1(new_n341), .B2(new_n194), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n304), .A2(new_n306), .A3(new_n311), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n324), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT19), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n331), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n334), .B2(new_n346), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n194), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n339), .B1(new_n350), .B2(new_n336), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n295), .B1(new_n340), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT20), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT86), .B(new_n354), .C1(new_n340), .C2(new_n351), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n354), .B(new_n295), .C1(new_n340), .C2(new_n351), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(KEYINPUT86), .ZN(new_n358));
  INV_X1    g172(.A(new_n351), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n327), .A2(new_n339), .A3(new_n336), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n295), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n359), .B2(new_n360), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n339), .B1(new_n327), .B2(new_n336), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n272), .B1(new_n340), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n361), .A2(new_n363), .B1(new_n365), .B2(G475), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n297), .A2(G952), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT21), .B(G898), .Z(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(G902), .A3(G953), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT89), .Z(new_n373));
  INV_X1    g187(.A(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n228), .A2(G122), .ZN(new_n376));
  INV_X1    g190(.A(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n196), .A2(G128), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n196), .A2(G128), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n209), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n213), .A2(G143), .ZN(new_n383));
  OAI21_X1  g197(.A(G134), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n375), .B1(new_n376), .B2(KEYINPUT14), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT88), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n376), .A2(KEYINPUT88), .A3(KEYINPUT14), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n378), .B(new_n385), .C1(new_n391), .C2(new_n377), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n383), .A2(new_n379), .A3(G134), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n375), .A2(new_n376), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G107), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n395), .B2(new_n378), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT13), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n381), .B1(new_n379), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n383), .A2(KEYINPUT87), .A3(KEYINPUT13), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n381), .B2(new_n397), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G134), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n392), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT9), .B(G234), .ZN(new_n406));
  INV_X1    g220(.A(G217), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(G953), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n392), .A2(new_n404), .A3(new_n408), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G478), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n392), .A2(new_n404), .A3(new_n408), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n408), .B1(new_n392), .B2(new_n404), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n272), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n414), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n357), .A2(new_n366), .A3(new_n373), .A4(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n226), .A3(G116), .ZN(new_n426));
  OAI211_X1 g240(.A(G113), .B(new_n426), .C1(new_n234), .C2(new_n425), .ZN(new_n427));
  AND2_X1   g241(.A1(KEYINPUT78), .A2(G101), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT78), .A2(G101), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G104), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G107), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT3), .B1(new_n431), .B2(G107), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n377), .A3(G104), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n432), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n377), .A2(G104), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G101), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n427), .A2(new_n436), .A3(new_n233), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n433), .A2(new_n435), .A3(new_n432), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G101), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n442), .A2(KEYINPUT4), .A3(new_n436), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n444), .A3(G101), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n237), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n440), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G122), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n448), .B(new_n440), .C1(new_n443), .C2(new_n446), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n258), .A2(G125), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n316), .B1(new_n248), .B2(new_n245), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n297), .A2(G224), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n453), .B2(new_n454), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n447), .A2(new_n460), .A3(new_n449), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n452), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n452), .A2(KEYINPUT80), .A3(new_n459), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI22_X1  g280(.A1(new_n453), .A2(new_n454), .B1(KEYINPUT82), .B2(new_n456), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI221_X1 g284(.A(new_n468), .B1(KEYINPUT82), .B2(new_n456), .C1(new_n453), .C2(new_n454), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n451), .A3(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n448), .B(KEYINPUT8), .Z(new_n473));
  INV_X1    g287(.A(new_n440), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n427), .A2(new_n233), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n436), .A2(new_n439), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(KEYINPUT81), .B2(new_n477), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n477), .A2(KEYINPUT81), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n272), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n466), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G210), .B1(G237), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n466), .A2(new_n484), .A3(new_n482), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n406), .B2(G902), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT77), .Z(new_n490));
  INV_X1    g304(.A(G101), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n432), .B2(new_n437), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n433), .A2(new_n435), .A3(new_n432), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n493), .B2(new_n430), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n258), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n200), .A2(new_n202), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n476), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n250), .A2(new_n251), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT12), .ZN(new_n502));
  XNOR2_X1  g316(.A(G110), .B(G140), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n297), .A2(G227), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n203), .A2(new_n494), .A3(KEYINPUT10), .A4(new_n217), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n442), .A2(KEYINPUT4), .A3(new_n436), .ZN(new_n508));
  XNOR2_X1  g322(.A(G143), .B(G146), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n246), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n244), .A2(new_n241), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n247), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n512), .A3(new_n445), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT10), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n496), .B2(new_n476), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n507), .A2(new_n513), .A3(new_n515), .A4(new_n499), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n499), .B1(new_n495), .B2(new_n497), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT12), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n502), .A2(new_n506), .A3(new_n516), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n507), .A2(new_n513), .A3(new_n515), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n500), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n506), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n517), .B(KEYINPUT12), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(KEYINPUT79), .A3(new_n506), .A4(new_n516), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G469), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n272), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n502), .A2(new_n516), .A3(new_n519), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n505), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n522), .A2(new_n506), .A3(new_n516), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(G469), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(G469), .A2(G902), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n490), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G214), .B1(G237), .B2(G902), .ZN(new_n538));
  AND4_X1   g352(.A1(new_n424), .A2(new_n488), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n407), .B1(G234), .B2(new_n272), .ZN(new_n540));
  NOR2_X1   g354(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n226), .B2(G128), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .ZN(new_n545));
  INV_X1    g359(.A(G110), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n226), .A2(G128), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n213), .A2(G119), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n547), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT24), .B(G110), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n548), .A2(KEYINPUT73), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n332), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n342), .A2(new_n345), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT75), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n544), .A2(new_n547), .A3(new_n545), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G110), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n551), .B2(new_n552), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n320), .A2(new_n194), .A3(new_n322), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(new_n324), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n555), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT22), .B(G137), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n297), .A2(G221), .A3(G234), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n564), .B(new_n565), .Z(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n555), .A2(new_n562), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n563), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n571), .B2(new_n566), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n542), .B1(new_n572), .B2(new_n272), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n555), .A2(new_n556), .A3(new_n562), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n556), .B1(new_n555), .B2(new_n562), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n563), .A2(new_n567), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n272), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n541), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n540), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n540), .A2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n294), .A2(new_n539), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n430), .B(KEYINPUT90), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT91), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n585), .B(new_n587), .ZN(G3));
  XNOR2_X1  g402(.A(new_n282), .B(KEYINPUT31), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT69), .B1(new_n262), .B2(new_n237), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n267), .ZN(new_n591));
  INV_X1    g405(.A(new_n263), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n254), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n256), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n253), .A2(KEYINPUT70), .A3(new_n254), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n286), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT71), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n265), .A2(new_n285), .A3(new_n286), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n589), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n291), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n600), .B2(G902), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(KEYINPUT92), .ZN(new_n604));
  INV_X1    g418(.A(G472), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n289), .B2(new_n272), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n537), .A2(new_n580), .A3(new_n582), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n486), .A2(new_n611), .A3(new_n487), .ZN(new_n612));
  INV_X1    g426(.A(new_n538), .ZN(new_n613));
  AOI211_X1 g427(.A(new_n485), .B(new_n481), .C1(new_n464), .C2(new_n465), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(KEYINPUT93), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n357), .A2(new_n366), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT33), .B1(new_n417), .B2(new_n418), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n410), .A2(new_n619), .A3(new_n411), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n618), .A2(new_n620), .A3(G478), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n413), .A2(new_n272), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n419), .B2(G478), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT94), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n622), .B1(new_n412), .B2(new_n413), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n618), .A2(new_n620), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n626), .B(new_n627), .C1(new_n413), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n617), .A2(new_n373), .A3(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n610), .A2(new_n616), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n365), .A2(G475), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n635), .A2(new_n636), .B1(new_n353), .B2(new_n356), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n365), .A2(KEYINPUT95), .A3(G475), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n373), .B(KEYINPUT96), .Z(new_n639));
  NAND4_X1  g453(.A1(new_n637), .A2(new_n421), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n610), .A2(new_n616), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT35), .B(G107), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND3_X1  g457(.A1(new_n488), .A2(new_n537), .A3(new_n538), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n540), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n572), .A2(new_n272), .A3(new_n542), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n578), .A2(new_n541), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n569), .B(KEYINPUT97), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n653), .A2(new_n654), .A3(new_n581), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n423), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n604), .A2(new_n645), .A3(new_n608), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  OAI21_X1  g474(.A(new_n537), .B1(new_n649), .B2(new_n655), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n616), .ZN(new_n662));
  INV_X1    g476(.A(new_n369), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n371), .A2(G900), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n663), .B1(new_n665), .B2(KEYINPUT98), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(KEYINPUT98), .B2(new_n665), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT99), .Z(new_n668));
  AND4_X1   g482(.A1(new_n421), .A2(new_n637), .A3(new_n638), .A4(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n662), .A2(new_n294), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XNOR2_X1  g485(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n668), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n537), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT102), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT40), .ZN(new_n676));
  INV_X1    g490(.A(new_n656), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n277), .A2(new_n192), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n269), .A2(new_n286), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n272), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n292), .B2(new_n293), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(KEYINPUT100), .B(new_n682), .C1(new_n292), .C2(new_n293), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n488), .B(KEYINPUT38), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n357), .A2(new_n366), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n422), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n538), .A3(new_n691), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n676), .A2(new_n677), .A3(new_n688), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n196), .ZN(G45));
  AND3_X1   g508(.A1(new_n617), .A2(new_n630), .A3(new_n668), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n662), .A2(new_n294), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  NOR2_X1   g511(.A1(new_n616), .A2(new_n631), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n529), .B1(new_n528), .B2(new_n272), .ZN(new_n699));
  AOI211_X1 g513(.A(G469), .B(G902), .C1(new_n525), .C2(new_n527), .ZN(new_n700));
  INV_X1    g514(.A(new_n489), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n294), .A2(new_n698), .A3(new_n584), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  AOI21_X1  g519(.A(new_n484), .B1(new_n466), .B2(new_n482), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n706), .A2(new_n614), .A3(KEYINPUT93), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n538), .B1(new_n487), .B2(new_n611), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n640), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n294), .A2(new_n709), .A3(new_n584), .A4(new_n702), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  AND3_X1   g525(.A1(new_n702), .A2(new_n612), .A3(new_n615), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n294), .A2(new_n712), .A3(new_n657), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT103), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n294), .A2(new_n712), .A3(new_n715), .A4(new_n657), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  NAND2_X1  g532(.A1(new_n270), .A2(new_n286), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n601), .B1(new_n719), .B2(new_n284), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n606), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n617), .A2(new_n421), .A3(new_n639), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n712), .A2(new_n584), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  NOR3_X1   g538(.A1(new_n656), .A2(new_n606), .A3(new_n720), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n695), .A3(new_n712), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT104), .B(G125), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G27));
  XNOR2_X1  g542(.A(new_n535), .B(KEYINPUT105), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n534), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n489), .B1(new_n700), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n706), .A2(new_n614), .A3(new_n613), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n695), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n294), .A3(new_n584), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(new_n294), .A3(KEYINPUT42), .A4(new_n584), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  NAND3_X1  g554(.A1(new_n486), .A2(new_n538), .A3(new_n487), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n583), .A2(new_n741), .A3(new_n731), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n294), .A2(new_n742), .A3(new_n669), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  NAND2_X1  g558(.A1(new_n532), .A2(new_n533), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n529), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n746), .B2(new_n745), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT106), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT46), .B1(new_n748), .B2(new_n729), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n700), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n701), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n673), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n756), .A3(new_n673), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT43), .B1(new_n690), .B2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g573(.A(new_n630), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n617), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n759), .B(new_n761), .Z(new_n762));
  NAND2_X1  g576(.A1(new_n604), .A2(new_n608), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n677), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n758), .A2(new_n733), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  XNOR2_X1  g583(.A(new_n753), .B(KEYINPUT47), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  INV_X1    g585(.A(new_n294), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n772), .A2(new_n583), .A3(new_n695), .A4(new_n733), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n770), .B2(new_n773), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  NOR2_X1   g592(.A1(new_n699), .A2(new_n700), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT49), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n490), .A2(new_n613), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n584), .A3(new_n761), .A4(new_n781), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n687), .A2(new_n689), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n779), .A2(new_n490), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n770), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT116), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n762), .A2(new_n663), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n721), .A2(new_n584), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n741), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n785), .A2(KEYINPUT116), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n786), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n790), .ZN(new_n794));
  INV_X1    g608(.A(new_n702), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n689), .A2(new_n538), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT50), .Z(new_n798));
  NOR2_X1   g612(.A1(new_n795), .A2(new_n741), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n584), .A2(new_n688), .A3(new_n663), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n690), .A3(new_n760), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n787), .A2(new_n725), .A3(new_n799), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n793), .A2(new_n798), .A3(KEYINPUT51), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n772), .A2(new_n583), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n787), .A2(new_n805), .A3(new_n799), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n800), .A2(new_n617), .A3(new_n630), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n794), .A2(new_n712), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n367), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n798), .A2(new_n803), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n785), .B2(new_n791), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n804), .B(new_n810), .C1(new_n812), .C2(KEYINPUT51), .ZN(new_n813));
  INV_X1    g627(.A(new_n696), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n726), .A2(new_n670), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n691), .A2(new_n612), .A3(new_n615), .ZN(new_n818));
  INV_X1    g632(.A(new_n668), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n818), .A2(new_n819), .A3(new_n731), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n687), .A2(new_n656), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n726), .A2(new_n670), .A3(KEYINPUT112), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n817), .A2(KEYINPUT52), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n726), .A2(new_n670), .A3(new_n696), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n821), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n353), .A2(new_n356), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n636), .A2(new_n635), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n421), .A2(new_n819), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n829), .A2(new_n830), .A3(new_n638), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n537), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n656), .A3(new_n741), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n294), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n741), .A2(new_n731), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n721), .A2(new_n677), .A3(new_n695), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n743), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT110), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n743), .A2(new_n835), .A3(new_n840), .A4(new_n837), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n839), .A2(new_n739), .A3(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n538), .B(new_n639), .C1(new_n706), .C2(new_n614), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n630), .B1(new_n357), .B2(new_n366), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n357), .A2(new_n366), .A3(new_n422), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n604), .A2(new_n608), .A3(new_n846), .A4(new_n609), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n703), .A2(new_n710), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n658), .A2(new_n723), .A3(new_n585), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n848), .A2(new_n717), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT111), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n839), .A2(new_n739), .A3(new_n841), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n848), .A2(new_n849), .A3(new_n717), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n828), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n824), .A2(new_n821), .A3(KEYINPUT52), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(new_n824), .B2(new_n821), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n842), .A2(new_n850), .A3(KEYINPUT111), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n854), .B1(new_n852), .B2(new_n853), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n856), .B(KEYINPUT54), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n852), .A2(new_n853), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n823), .A2(new_n827), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n862), .B2(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT115), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n864), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n813), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n783), .B1(new_n876), .B2(new_n877), .ZN(G75));
  NOR2_X1   g692(.A1(new_n297), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n867), .A2(new_n868), .ZN(new_n881));
  INV_X1    g695(.A(new_n862), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n863), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n272), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(G210), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n452), .A2(new_n461), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n459), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n880), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n885), .B2(new_n889), .ZN(G51));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n883), .B2(new_n865), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n862), .A2(KEYINPUT53), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n893), .B(new_n866), .C1(new_n894), .C2(new_n881), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(new_n869), .C1(new_n862), .C2(KEYINPUT53), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n892), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n729), .B(KEYINPUT57), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n528), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n883), .A2(new_n272), .A3(new_n748), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n879), .B1(new_n903), .B2(new_n904), .ZN(G54));
  NAND3_X1  g719(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n340), .A2(new_n351), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n879), .ZN(G60));
  XNOR2_X1  g724(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n623), .B(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n872), .B2(new_n874), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n880), .B1(new_n913), .B2(new_n628), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n618), .B2(new_n620), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n900), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n900), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n917), .B2(new_n919), .ZN(G63));
  INV_X1    g734(.A(new_n883), .ZN(new_n921));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT121), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n572), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n921), .A2(new_n653), .A3(new_n654), .A4(new_n924), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n880), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n927), .A2(KEYINPUT61), .A3(new_n880), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(G66));
  NAND3_X1  g747(.A1(new_n370), .A2(G224), .A3(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n853), .B2(G953), .ZN(new_n935));
  INV_X1    g749(.A(G898), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n886), .B1(new_n936), .B2(G953), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  NAND2_X1  g752(.A1(new_n817), .A2(new_n822), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n693), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT62), .Z(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  INV_X1    g756(.A(new_n805), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n844), .A2(new_n845), .ZN(new_n944));
  OR4_X1    g758(.A1(new_n943), .A2(new_n675), .A3(new_n741), .A4(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n768), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n942), .B1(new_n768), .B2(new_n945), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n777), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n297), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n274), .A2(new_n275), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT122), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n348), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n739), .B(new_n743), .C1(new_n775), .C2(new_n776), .ZN(new_n956));
  INV_X1    g770(.A(new_n818), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n805), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n755), .B2(new_n757), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT125), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n939), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n768), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n768), .A2(KEYINPUT124), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n961), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n961), .B2(new_n967), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(G953), .ZN(new_n971));
  INV_X1    g785(.A(G900), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n953), .B1(new_n972), .B2(new_n297), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n955), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n297), .B1(G227), .B2(G900), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n977), .B(new_n955), .C1(new_n971), .C2(new_n973), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  OR2_X1    g795(.A1(new_n941), .A2(new_n949), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n853), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n879), .B1(new_n983), .B2(new_n679), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n969), .A2(new_n970), .A3(new_n853), .ZN(new_n985));
  INV_X1    g799(.A(new_n981), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n278), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n679), .A2(new_n278), .A3(new_n986), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n856), .B(new_n988), .C1(new_n862), .C2(new_n863), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT127), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n984), .A2(new_n987), .A3(new_n990), .ZN(G57));
endmodule


