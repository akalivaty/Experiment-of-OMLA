

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761;

  INV_X1 U375 ( .A(G953), .ZN(n750) );
  XOR2_X1 U376 ( .A(G143), .B(G140), .Z(n355) );
  AND2_X1 U377 ( .A1(n398), .A2(n362), .ZN(n356) );
  INV_X1 U378 ( .A(n636), .ZN(n375) );
  NOR2_X2 U379 ( .A1(n636), .A2(n677), .ZN(n729) );
  INV_X1 U380 ( .A(KEYINPUT48), .ZN(n441) );
  AND2_X1 U381 ( .A1(n425), .A2(n424), .ZN(n423) );
  XNOR2_X1 U382 ( .A(n418), .B(n552), .ZN(n417) );
  XNOR2_X1 U383 ( .A(n394), .B(KEYINPUT40), .ZN(n382) );
  AND2_X1 U384 ( .A1(n391), .A2(n468), .ZN(n569) );
  XNOR2_X1 U385 ( .A(n561), .B(KEYINPUT19), .ZN(n591) );
  NAND2_X1 U386 ( .A1(n568), .A2(n678), .ZN(n561) );
  AND2_X1 U387 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U388 ( .A1(n689), .A2(n688), .ZN(n582) );
  OR2_X1 U389 ( .A1(n565), .A2(n563), .ZN(n661) );
  XNOR2_X1 U390 ( .A(n404), .B(n363), .ZN(n547) );
  XNOR2_X1 U391 ( .A(n415), .B(n361), .ZN(n563) );
  XNOR2_X1 U392 ( .A(n477), .B(n476), .ZN(n731) );
  OR2_X1 U393 ( .A1(n726), .A2(G902), .ZN(n415) );
  XNOR2_X1 U394 ( .A(n748), .B(n472), .ZN(n477) );
  XNOR2_X1 U395 ( .A(n412), .B(n541), .ZN(n544) );
  XNOR2_X1 U396 ( .A(n515), .B(n457), .ZN(n495) );
  XNOR2_X1 U397 ( .A(n531), .B(n491), .ZN(n748) );
  XNOR2_X1 U398 ( .A(n511), .B(n469), .ZN(n531) );
  XNOR2_X1 U399 ( .A(n746), .B(n456), .ZN(n515) );
  XNOR2_X1 U400 ( .A(n393), .B(G125), .ZN(n511) );
  INV_X1 U401 ( .A(G146), .ZN(n393) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n523) );
  XNOR2_X1 U403 ( .A(n405), .B(KEYINPUT4), .ZN(n746) );
  INV_X1 U404 ( .A(n563), .ZN(n566) );
  NAND2_X1 U405 ( .A1(n591), .A2(n590), .ZN(n594) );
  XNOR2_X1 U406 ( .A(n498), .B(n497), .ZN(n560) );
  OR2_X1 U407 ( .A1(n721), .A2(G902), .ZN(n498) );
  XNOR2_X1 U408 ( .A(n508), .B(n357), .ZN(n379) );
  XNOR2_X1 U409 ( .A(n505), .B(n504), .ZN(n508) );
  XNOR2_X1 U410 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n504) );
  XOR2_X1 U411 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n527) );
  XNOR2_X1 U412 ( .A(G131), .B(KEYINPUT96), .ZN(n526) );
  OR2_X1 U413 ( .A1(n731), .A2(G902), .ZN(n404) );
  XNOR2_X1 U414 ( .A(n481), .B(n482), .ZN(n446) );
  INV_X1 U415 ( .A(n561), .ZN(n435) );
  NAND2_X1 U416 ( .A1(n381), .A2(n614), .ZN(n380) );
  INV_X1 U417 ( .A(n549), .ZN(n381) );
  INV_X1 U418 ( .A(n547), .ZN(n689) );
  XNOR2_X1 U419 ( .A(n392), .B(n360), .ZN(n533) );
  XNOR2_X1 U420 ( .A(n379), .B(n359), .ZN(n646) );
  XNOR2_X1 U421 ( .A(n421), .B(n420), .ZN(n711) );
  INV_X1 U422 ( .A(KEYINPUT41), .ZN(n420) );
  AND2_X1 U423 ( .A1(n679), .A2(n384), .ZN(n421) );
  NOR2_X1 U424 ( .A1(n681), .A2(n385), .ZN(n384) );
  XNOR2_X1 U425 ( .A(n522), .B(n366), .ZN(n546) );
  XNOR2_X1 U426 ( .A(n427), .B(KEYINPUT22), .ZN(n604) );
  AND2_X1 U427 ( .A1(n599), .A2(n688), .ZN(n428) );
  AND2_X1 U428 ( .A1(n403), .A2(n614), .ZN(n562) );
  BUF_X1 U429 ( .A(n689), .Z(n395) );
  INV_X1 U430 ( .A(G475), .ZN(n374) );
  NAND2_X1 U431 ( .A1(n376), .A2(n375), .ZN(n431) );
  NOR2_X1 U432 ( .A1(n677), .A2(n377), .ZN(n376) );
  NOR2_X1 U433 ( .A1(n660), .A2(n682), .ZN(n564) );
  XNOR2_X1 U434 ( .A(KEYINPUT83), .B(KEYINPUT46), .ZN(n552) );
  NAND2_X1 U435 ( .A1(G953), .A2(G902), .ZN(n586) );
  NOR2_X1 U436 ( .A1(G902), .A2(G237), .ZN(n459) );
  AND2_X1 U437 ( .A1(n609), .A2(n608), .ZN(n610) );
  INV_X1 U438 ( .A(KEYINPUT10), .ZN(n469) );
  XOR2_X1 U439 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n525) );
  XNOR2_X1 U440 ( .A(n528), .B(n529), .ZN(n392) );
  XNOR2_X1 U441 ( .A(n478), .B(G902), .ZN(n633) );
  XNOR2_X1 U442 ( .A(G134), .B(G131), .ZN(n744) );
  XOR2_X1 U443 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n510) );
  XNOR2_X1 U444 ( .A(KEYINPUT87), .B(KEYINPUT76), .ZN(n509) );
  INV_X1 U445 ( .A(G101), .ZN(n456) );
  INV_X1 U446 ( .A(KEYINPUT82), .ZN(n437) );
  NOR2_X1 U447 ( .A1(n548), .A2(n549), .ZN(n553) );
  XNOR2_X1 U448 ( .A(G119), .B(KEYINPUT3), .ZN(n454) );
  XNOR2_X1 U449 ( .A(G137), .B(G116), .ZN(n451) );
  INV_X1 U450 ( .A(KEYINPUT92), .ZN(n450) );
  XOR2_X1 U451 ( .A(G113), .B(KEYINPUT5), .Z(n449) );
  XNOR2_X1 U452 ( .A(G119), .B(G128), .ZN(n470) );
  XOR2_X1 U453 ( .A(KEYINPUT24), .B(G110), .Z(n471) );
  NAND2_X1 U454 ( .A1(G234), .A2(n750), .ZN(n473) );
  XOR2_X1 U455 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n539) );
  XNOR2_X1 U456 ( .A(G134), .B(G122), .ZN(n538) );
  XNOR2_X1 U457 ( .A(n413), .B(n501), .ZN(n412) );
  XNOR2_X1 U458 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n414) );
  XNOR2_X1 U459 ( .A(G107), .B(G104), .ZN(n487) );
  INV_X1 U460 ( .A(KEYINPUT72), .ZN(n488) );
  XNOR2_X1 U461 ( .A(G140), .B(G137), .ZN(n491) );
  NAND2_X1 U462 ( .A1(G234), .A2(G237), .ZN(n462) );
  NAND2_X1 U463 ( .A1(n561), .A2(n558), .ZN(n433) );
  INV_X1 U464 ( .A(KEYINPUT34), .ZN(n396) );
  NOR2_X1 U465 ( .A1(n380), .A2(n582), .ZN(n391) );
  INV_X1 U466 ( .A(G902), .ZN(n534) );
  INV_X1 U467 ( .A(KEYINPUT89), .ZN(n595) );
  BUF_X1 U468 ( .A(n625), .Z(n399) );
  XNOR2_X1 U469 ( .A(n419), .B(KEYINPUT42), .ZN(n551) );
  NAND2_X1 U470 ( .A1(n546), .A2(n666), .ZN(n641) );
  NAND2_X1 U471 ( .A1(n546), .A2(n545), .ZN(n394) );
  AND2_X1 U472 ( .A1(n602), .A2(n378), .ZN(n603) );
  AND2_X1 U473 ( .A1(n601), .A2(n547), .ZN(n378) );
  XNOR2_X1 U474 ( .A(n621), .B(n400), .ZN(n667) );
  XNOR2_X1 U475 ( .A(n401), .B(KEYINPUT31), .ZN(n400) );
  INV_X1 U476 ( .A(KEYINPUT94), .ZN(n401) );
  INV_X1 U477 ( .A(KEYINPUT60), .ZN(n387) );
  NAND2_X1 U478 ( .A1(n430), .A2(n429), .ZN(n389) );
  XNOR2_X1 U479 ( .A(n431), .B(n367), .ZN(n430) );
  XNOR2_X1 U480 ( .A(n551), .B(G137), .ZN(G39) );
  XNOR2_X1 U481 ( .A(n560), .B(n559), .ZN(n694) );
  XOR2_X1 U482 ( .A(n507), .B(n506), .Z(n357) );
  XOR2_X1 U483 ( .A(G472), .B(KEYINPUT93), .Z(n358) );
  XOR2_X1 U484 ( .A(n515), .B(n514), .Z(n359) );
  XOR2_X1 U485 ( .A(n525), .B(n524), .Z(n360) );
  XOR2_X1 U486 ( .A(n537), .B(KEYINPUT101), .Z(n361) );
  AND2_X1 U487 ( .A1(n694), .A2(n433), .ZN(n362) );
  XOR2_X1 U488 ( .A(n480), .B(n446), .Z(n363) );
  INV_X1 U489 ( .A(n694), .ZN(n408) );
  AND2_X1 U490 ( .A1(n435), .A2(n434), .ZN(n364) );
  AND2_X1 U491 ( .A1(n641), .A2(KEYINPUT2), .ZN(n365) );
  XOR2_X1 U492 ( .A(n521), .B(n520), .Z(n366) );
  XOR2_X1 U493 ( .A(n646), .B(n645), .Z(n367) );
  XOR2_X1 U494 ( .A(n638), .B(n637), .Z(n368) );
  XOR2_X1 U495 ( .A(n643), .B(n642), .Z(n369) );
  INV_X1 U496 ( .A(n733), .ZN(n429) );
  XNOR2_X1 U497 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n370) );
  NAND2_X1 U498 ( .A1(n371), .A2(n375), .ZN(n639) );
  NOR2_X1 U499 ( .A1(n677), .A2(n372), .ZN(n371) );
  INV_X1 U500 ( .A(G472), .ZN(n372) );
  NAND2_X1 U501 ( .A1(n373), .A2(n375), .ZN(n644) );
  NOR2_X1 U502 ( .A1(n677), .A2(n374), .ZN(n373) );
  INV_X1 U503 ( .A(G210), .ZN(n377) );
  XNOR2_X1 U504 ( .A(n495), .B(n458), .ZN(n638) );
  XNOR2_X1 U505 ( .A(n379), .B(G101), .ZN(n738) );
  NAND2_X1 U506 ( .A1(n382), .A2(n551), .ZN(n418) );
  XNOR2_X1 U507 ( .A(n382), .B(G131), .ZN(G33) );
  NOR2_X1 U508 ( .A1(n383), .A2(KEYINPUT65), .ZN(n606) );
  XNOR2_X1 U509 ( .A(n383), .B(KEYINPUT65), .ZN(n611) );
  XNOR2_X1 U510 ( .A(n383), .B(G122), .ZN(n757) );
  XNOR2_X2 U511 ( .A(n598), .B(KEYINPUT35), .ZN(n383) );
  NAND2_X1 U512 ( .A1(n679), .A2(n678), .ZN(n386) );
  INV_X1 U513 ( .A(n678), .ZN(n385) );
  NOR2_X1 U514 ( .A1(n682), .A2(n386), .ZN(n683) );
  OR2_X2 U515 ( .A1(n638), .A2(G902), .ZN(n406) );
  XNOR2_X1 U516 ( .A(n388), .B(n387), .ZN(G60) );
  NAND2_X1 U517 ( .A1(n390), .A2(n429), .ZN(n388) );
  XNOR2_X1 U518 ( .A(n613), .B(KEYINPUT6), .ZN(n625) );
  XNOR2_X1 U519 ( .A(n389), .B(n370), .ZN(G51) );
  XNOR2_X1 U520 ( .A(n644), .B(n369), .ZN(n390) );
  INV_X1 U521 ( .A(n669), .ZN(n439) );
  NAND2_X2 U522 ( .A1(n356), .A2(n432), .ZN(n436) );
  XNOR2_X1 U523 ( .A(n397), .B(n396), .ZN(n402) );
  NAND2_X1 U524 ( .A1(n612), .A2(n710), .ZN(n397) );
  NAND2_X1 U525 ( .A1(n562), .A2(n711), .ZN(n419) );
  AND2_X1 U526 ( .A1(n416), .A2(n575), .ZN(n411) );
  XNOR2_X1 U527 ( .A(n438), .B(n437), .ZN(n629) );
  NAND2_X1 U528 ( .A1(n409), .A2(n364), .ZN(n398) );
  NOR2_X1 U529 ( .A1(n623), .A2(n426), .ZN(n424) );
  NAND2_X1 U530 ( .A1(n611), .A2(n610), .ZN(n422) );
  NAND2_X1 U531 ( .A1(n402), .A2(n597), .ZN(n598) );
  XNOR2_X1 U532 ( .A(n445), .B(KEYINPUT81), .ZN(n444) );
  XNOR2_X1 U533 ( .A(n410), .B(n441), .ZN(n440) );
  NAND2_X1 U534 ( .A1(n440), .A2(n439), .ZN(n438) );
  NAND2_X1 U535 ( .A1(n530), .A2(n501), .ZN(n502) );
  XNOR2_X2 U536 ( .A(n499), .B(G122), .ZN(n530) );
  NAND2_X1 U537 ( .A1(n423), .A2(n422), .ZN(n627) );
  NAND2_X1 U538 ( .A1(n562), .A2(n591), .ZN(n660) );
  XNOR2_X1 U539 ( .A(n550), .B(KEYINPUT28), .ZN(n403) );
  XNOR2_X1 U540 ( .A(n405), .B(n414), .ZN(n413) );
  XNOR2_X2 U541 ( .A(G143), .B(G128), .ZN(n405) );
  NOR2_X1 U542 ( .A1(n625), .A2(n661), .ZN(n554) );
  XNOR2_X2 U543 ( .A(n406), .B(n358), .ZN(n613) );
  NAND2_X1 U544 ( .A1(n407), .A2(n558), .ZN(n432) );
  INV_X1 U545 ( .A(n409), .ZN(n407) );
  AND2_X1 U546 ( .A1(n409), .A2(n408), .ZN(n576) );
  XNOR2_X2 U547 ( .A(n555), .B(KEYINPUT106), .ZN(n409) );
  NAND2_X1 U548 ( .A1(n411), .A2(n417), .ZN(n410) );
  XNOR2_X1 U549 ( .A(n759), .B(KEYINPUT84), .ZN(n416) );
  NAND2_X1 U550 ( .A1(n607), .A2(KEYINPUT44), .ZN(n425) );
  INV_X1 U551 ( .A(n647), .ZN(n426) );
  NAND2_X1 U552 ( .A1(n618), .A2(n428), .ZN(n427) );
  XNOR2_X2 U553 ( .A(n594), .B(n593), .ZN(n618) );
  NAND2_X1 U554 ( .A1(n444), .A2(n670), .ZN(n628) );
  INV_X1 U555 ( .A(n558), .ZN(n434) );
  XNOR2_X2 U556 ( .A(n436), .B(KEYINPUT110), .ZN(n759) );
  XNOR2_X1 U557 ( .A(n442), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U558 ( .A1(n443), .A2(n429), .ZN(n442) );
  XNOR2_X1 U559 ( .A(n639), .B(n368), .ZN(n443) );
  NAND2_X1 U560 ( .A1(n629), .A2(n365), .ZN(n445) );
  XNOR2_X2 U561 ( .A(n628), .B(KEYINPUT73), .ZN(n677) );
  AND2_X1 U562 ( .A1(G224), .A2(n750), .ZN(n447) );
  XNOR2_X1 U563 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U564 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U565 ( .A(n511), .B(n447), .ZN(n512) );
  INV_X1 U566 ( .A(KEYINPUT64), .ZN(n592) );
  XNOR2_X1 U567 ( .A(n513), .B(n512), .ZN(n514) );
  INV_X1 U568 ( .A(KEYINPUT86), .ZN(n556) );
  XNOR2_X1 U569 ( .A(n592), .B(KEYINPUT0), .ZN(n593) );
  XNOR2_X1 U570 ( .A(n557), .B(n556), .ZN(n558) );
  INV_X1 U571 ( .A(KEYINPUT80), .ZN(n630) );
  NOR2_X1 U572 ( .A1(n408), .A2(n600), .ZN(n601) );
  XNOR2_X1 U573 ( .A(n618), .B(n595), .ZN(n612) );
  NAND2_X1 U574 ( .A1(n523), .A2(G210), .ZN(n448) );
  XNOR2_X1 U575 ( .A(n449), .B(n448), .ZN(n453) );
  XNOR2_X1 U576 ( .A(n454), .B(KEYINPUT67), .ZN(n507) );
  XNOR2_X1 U577 ( .A(n455), .B(n507), .ZN(n458) );
  XNOR2_X1 U578 ( .A(n744), .B(G146), .ZN(n457) );
  XNOR2_X1 U579 ( .A(n459), .B(KEYINPUT71), .ZN(n516) );
  NAND2_X1 U580 ( .A1(G214), .A2(n516), .ZN(n678) );
  NAND2_X1 U581 ( .A1(n613), .A2(n678), .ZN(n461) );
  INV_X1 U582 ( .A(KEYINPUT30), .ZN(n460) );
  XNOR2_X1 U583 ( .A(n461), .B(n460), .ZN(n468) );
  XOR2_X1 U584 ( .A(KEYINPUT14), .B(n462), .Z(n708) );
  NOR2_X1 U585 ( .A1(n708), .A2(n586), .ZN(n463) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(n463), .Z(n464) );
  NOR2_X1 U587 ( .A1(G900), .A2(n464), .ZN(n465) );
  XOR2_X1 U588 ( .A(KEYINPUT105), .B(n465), .Z(n467) );
  NAND2_X1 U589 ( .A1(n750), .A2(G952), .ZN(n585) );
  NOR2_X1 U590 ( .A1(n708), .A2(n585), .ZN(n466) );
  NOR2_X1 U591 ( .A1(n467), .A2(n466), .ZN(n549) );
  XNOR2_X1 U592 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(KEYINPUT78), .Z(n475) );
  XOR2_X1 U594 ( .A(KEYINPUT8), .B(n473), .Z(n542) );
  NAND2_X1 U595 ( .A1(G221), .A2(n542), .ZN(n474) );
  XNOR2_X1 U596 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U597 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n481) );
  XNOR2_X1 U598 ( .A(KEYINPUT88), .B(KEYINPUT15), .ZN(n478) );
  NAND2_X1 U599 ( .A1(n633), .A2(G234), .ZN(n479) );
  XNOR2_X1 U600 ( .A(KEYINPUT20), .B(n479), .ZN(n483) );
  NAND2_X1 U601 ( .A1(n483), .A2(G217), .ZN(n480) );
  INV_X1 U602 ( .A(KEYINPUT91), .ZN(n482) );
  NAND2_X1 U603 ( .A1(n483), .A2(G221), .ZN(n485) );
  INV_X1 U604 ( .A(KEYINPUT21), .ZN(n484) );
  XNOR2_X1 U605 ( .A(n485), .B(n484), .ZN(n688) );
  NAND2_X1 U606 ( .A1(n750), .A2(G227), .ZN(n486) );
  XNOR2_X1 U607 ( .A(n487), .B(n486), .ZN(n489) );
  XNOR2_X1 U608 ( .A(n488), .B(G110), .ZN(n506) );
  XNOR2_X1 U609 ( .A(n489), .B(n506), .ZN(n493) );
  XNOR2_X1 U610 ( .A(KEYINPUT75), .B(KEYINPUT90), .ZN(n490) );
  XNOR2_X1 U611 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U612 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U613 ( .A(n495), .B(n494), .ZN(n721) );
  INV_X1 U614 ( .A(KEYINPUT66), .ZN(n496) );
  XNOR2_X1 U615 ( .A(n496), .B(G469), .ZN(n497) );
  INV_X1 U616 ( .A(n560), .ZN(n614) );
  XOR2_X1 U617 ( .A(G116), .B(G107), .Z(n540) );
  XNOR2_X2 U618 ( .A(G113), .B(G104), .ZN(n499) );
  INV_X1 U619 ( .A(n530), .ZN(n500) );
  NAND2_X1 U620 ( .A1(n540), .A2(n500), .ZN(n503) );
  INV_X1 U621 ( .A(n540), .ZN(n501) );
  NAND2_X1 U622 ( .A1(n503), .A2(n502), .ZN(n505) );
  XNOR2_X1 U623 ( .A(n510), .B(n509), .ZN(n513) );
  NAND2_X1 U624 ( .A1(n646), .A2(n633), .ZN(n518) );
  AND2_X1 U625 ( .A1(G210), .A2(n516), .ZN(n517) );
  XNOR2_X2 U626 ( .A(n518), .B(n517), .ZN(n568) );
  INV_X1 U627 ( .A(KEYINPUT38), .ZN(n519) );
  XNOR2_X1 U628 ( .A(n568), .B(n519), .ZN(n679) );
  NAND2_X1 U629 ( .A1(n569), .A2(n679), .ZN(n522) );
  XNOR2_X1 U630 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n521) );
  INV_X1 U631 ( .A(KEYINPUT69), .ZN(n520) );
  NAND2_X1 U632 ( .A1(G214), .A2(n523), .ZN(n524) );
  XNOR2_X1 U633 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U634 ( .A(KEYINPUT97), .B(n355), .ZN(n529) );
  XNOR2_X1 U635 ( .A(n530), .B(n531), .ZN(n532) );
  XNOR2_X1 U636 ( .A(n533), .B(n532), .ZN(n643) );
  NAND2_X1 U637 ( .A1(n643), .A2(n534), .ZN(n536) );
  XNOR2_X1 U638 ( .A(KEYINPUT13), .B(G475), .ZN(n535) );
  XNOR2_X1 U639 ( .A(n536), .B(n535), .ZN(n565) );
  XNOR2_X1 U640 ( .A(G478), .B(KEYINPUT102), .ZN(n537) );
  XNOR2_X1 U641 ( .A(n539), .B(n538), .ZN(n541) );
  NAND2_X1 U642 ( .A1(G217), .A2(n542), .ZN(n543) );
  XNOR2_X1 U643 ( .A(n544), .B(n543), .ZN(n726) );
  INV_X1 U644 ( .A(n661), .ZN(n545) );
  NAND2_X1 U645 ( .A1(n565), .A2(n566), .ZN(n681) );
  NAND2_X1 U646 ( .A1(n547), .A2(n688), .ZN(n548) );
  AND2_X1 U647 ( .A1(n613), .A2(n553), .ZN(n550) );
  XNOR2_X1 U648 ( .A(KEYINPUT109), .B(KEYINPUT36), .ZN(n557) );
  INV_X1 U649 ( .A(KEYINPUT1), .ZN(n559) );
  AND2_X1 U650 ( .A1(n565), .A2(n563), .ZN(n666) );
  INV_X1 U651 ( .A(n666), .ZN(n657) );
  AND2_X1 U652 ( .A1(n661), .A2(n657), .ZN(n682) );
  XNOR2_X1 U653 ( .A(n564), .B(KEYINPUT47), .ZN(n574) );
  OR2_X1 U654 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U655 ( .A(KEYINPUT103), .B(n567), .Z(n596) );
  INV_X1 U656 ( .A(n568), .ZN(n580) );
  NOR2_X1 U657 ( .A1(n596), .A2(n580), .ZN(n570) );
  NAND2_X1 U658 ( .A1(n570), .A2(n569), .ZN(n572) );
  INV_X1 U659 ( .A(KEYINPUT108), .ZN(n571) );
  XNOR2_X1 U660 ( .A(n572), .B(n571), .ZN(n761) );
  INV_X1 U661 ( .A(n761), .ZN(n573) );
  AND2_X1 U662 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n678), .A2(n576), .ZN(n577) );
  XNOR2_X1 U664 ( .A(n577), .B(KEYINPUT43), .ZN(n579) );
  INV_X1 U665 ( .A(KEYINPUT107), .ZN(n578) );
  XNOR2_X1 U666 ( .A(n579), .B(n578), .ZN(n581) );
  AND2_X1 U667 ( .A1(n581), .A2(n580), .ZN(n669) );
  INV_X1 U668 ( .A(n582), .ZN(n695) );
  NAND2_X1 U669 ( .A1(n695), .A2(n694), .ZN(n619) );
  NOR2_X1 U670 ( .A1(n399), .A2(n619), .ZN(n584) );
  XNOR2_X1 U671 ( .A(KEYINPUT33), .B(KEYINPUT68), .ZN(n583) );
  XNOR2_X1 U672 ( .A(n584), .B(n583), .ZN(n686) );
  INV_X1 U673 ( .A(n686), .ZN(n710) );
  INV_X1 U674 ( .A(n585), .ZN(n588) );
  NOR2_X1 U675 ( .A1(G898), .A2(n586), .ZN(n587) );
  NOR2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U677 ( .A1(n708), .A2(n589), .ZN(n590) );
  XNOR2_X1 U678 ( .A(n596), .B(KEYINPUT77), .ZN(n597) );
  INV_X1 U679 ( .A(n681), .ZN(n599) );
  INV_X1 U680 ( .A(n604), .ZN(n602) );
  INV_X1 U681 ( .A(n399), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n603), .B(KEYINPUT32), .ZN(n758) );
  NOR2_X1 U683 ( .A1(n604), .A2(n694), .ZN(n624) );
  INV_X1 U684 ( .A(n613), .ZN(n691) );
  NAND2_X1 U685 ( .A1(n624), .A2(n691), .ZN(n605) );
  NOR2_X1 U686 ( .A1(n395), .A2(n605), .ZN(n655) );
  NOR2_X1 U687 ( .A1(n758), .A2(n655), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n606), .A2(n609), .ZN(n607) );
  INV_X1 U689 ( .A(KEYINPUT44), .ZN(n608) );
  INV_X1 U690 ( .A(n612), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n613), .A2(n582), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n652) );
  INV_X1 U694 ( .A(n618), .ZN(n620) );
  OR2_X1 U695 ( .A1(n691), .A2(n619), .ZN(n699) );
  NOR2_X1 U696 ( .A1(n620), .A2(n699), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n652), .A2(n667), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n682), .A2(n622), .ZN(n623) );
  AND2_X1 U699 ( .A1(n399), .A2(n624), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n626), .A2(n395), .ZN(n647) );
  XNOR2_X2 U701 ( .A(n627), .B(KEYINPUT45), .ZN(n670) );
  NAND2_X1 U702 ( .A1(n629), .A2(n641), .ZN(n631) );
  XNOR2_X2 U703 ( .A(n631), .B(n630), .ZN(n749) );
  NAND2_X1 U704 ( .A1(n670), .A2(n749), .ZN(n632) );
  INV_X1 U705 ( .A(KEYINPUT2), .ZN(n672) );
  NAND2_X1 U706 ( .A1(n632), .A2(n672), .ZN(n635) );
  INV_X1 U707 ( .A(n633), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U709 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n637) );
  INV_X1 U710 ( .A(G952), .ZN(n640) );
  AND2_X1 U711 ( .A1(n640), .A2(G953), .ZN(n733) );
  XNOR2_X1 U712 ( .A(n641), .B(G134), .ZN(G36) );
  XNOR2_X1 U713 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n642) );
  XNOR2_X1 U714 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n645) );
  XNOR2_X1 U715 ( .A(G101), .B(n647), .ZN(G3) );
  NAND2_X1 U716 ( .A1(n652), .A2(n545), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n648), .B(G104), .ZN(G6) );
  XOR2_X1 U718 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n650) );
  XNOR2_X1 U719 ( .A(G107), .B(KEYINPUT26), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT27), .B(n651), .Z(n654) );
  NAND2_X1 U722 ( .A1(n652), .A2(n666), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(G9) );
  XOR2_X1 U724 ( .A(G110), .B(n655), .Z(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT114), .B(n656), .ZN(G12) );
  NOR2_X1 U726 ( .A1(n657), .A2(n660), .ZN(n659) );
  XNOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(G30) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U730 ( .A(G146), .B(KEYINPUT115), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(G48) );
  NAND2_X1 U732 ( .A1(n667), .A2(n545), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(KEYINPUT116), .ZN(n665) );
  XNOR2_X1 U734 ( .A(G113), .B(n665), .ZN(G15) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n668), .B(G116), .ZN(G18) );
  XOR2_X1 U737 ( .A(G140), .B(n669), .Z(G42) );
  XOR2_X1 U738 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n718) );
  NOR2_X1 U739 ( .A1(n670), .A2(KEYINPUT2), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(KEYINPUT79), .ZN(n675) );
  INV_X1 U741 ( .A(n749), .ZN(n673) );
  NAND2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n715) );
  XNOR2_X1 U745 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n706) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U750 ( .A(KEYINPUT118), .B(n687), .Z(n704) );
  NOR2_X1 U751 ( .A1(n395), .A2(n688), .ZN(n690) );
  XNOR2_X1 U752 ( .A(n690), .B(KEYINPUT49), .ZN(n692) );
  NAND2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U754 ( .A(n693), .B(KEYINPUT117), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U756 ( .A(KEYINPUT50), .B(n696), .Z(n697) );
  NAND2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U759 ( .A(KEYINPUT51), .B(n701), .Z(n702) );
  NAND2_X1 U760 ( .A1(n711), .A2(n702), .ZN(n703) );
  NAND2_X1 U761 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U762 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U764 ( .A1(G952), .A2(n709), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n716), .A2(n750), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(G75) );
  NAND2_X1 U770 ( .A1(n729), .A2(G469), .ZN(n724) );
  XOR2_X1 U771 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n720) );
  XNOR2_X1 U772 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n722) );
  XOR2_X1 U774 ( .A(n722), .B(n721), .Z(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n733), .A2(n725), .ZN(G54) );
  NAND2_X1 U777 ( .A1(n729), .A2(G478), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n726), .B(n727), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n733), .A2(n728), .ZN(G63) );
  NAND2_X1 U780 ( .A1(n729), .A2(G217), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U782 ( .A1(n733), .A2(n732), .ZN(G66) );
  NAND2_X1 U783 ( .A1(n750), .A2(n670), .ZN(n737) );
  NAND2_X1 U784 ( .A1(G953), .A2(G224), .ZN(n734) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n734), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(G898), .ZN(n736) );
  NAND2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n742) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n738), .ZN(n740) );
  NOR2_X1 U789 ( .A1(G898), .A2(n750), .ZN(n739) );
  NOR2_X1 U790 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U791 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U792 ( .A(KEYINPUT126), .B(n743), .ZN(G69) );
  INV_X1 U793 ( .A(n744), .ZN(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n748), .B(n747), .ZN(n752) );
  XOR2_X1 U796 ( .A(n752), .B(n749), .Z(n751) );
  NAND2_X1 U797 ( .A1(n751), .A2(n750), .ZN(n756) );
  XNOR2_X1 U798 ( .A(G227), .B(n752), .ZN(n753) );
  NAND2_X1 U799 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n754), .A2(G953), .ZN(n755) );
  NAND2_X1 U801 ( .A1(n756), .A2(n755), .ZN(G72) );
  XNOR2_X1 U802 ( .A(n757), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U803 ( .A(G119), .B(n758), .Z(G21) );
  XOR2_X1 U804 ( .A(n759), .B(G125), .Z(n760) );
  XNOR2_X1 U805 ( .A(KEYINPUT37), .B(n760), .ZN(G27) );
  XOR2_X1 U806 ( .A(G143), .B(n761), .Z(G45) );
endmodule

