//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT27), .B(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT28), .B1(new_n205), .B2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  OR3_X1    g015(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT28), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n219), .A3(new_n208), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n206), .A2(new_n210), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n209), .A2(new_n227), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT25), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238));
  NOR4_X1   g037(.A1(new_n235), .A2(new_n229), .A3(new_n232), .A4(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n221), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G120gat), .ZN(new_n243));
  INV_X1    g042(.A(G120gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(G113gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G127gat), .B(G134gat), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n242), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(G113gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n244), .B2(G113gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n249), .B1(new_n254), .B2(KEYINPUT67), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n244), .A3(G113gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT66), .B1(new_n242), .B2(G120gat), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT67), .B(new_n256), .C1(new_n257), .C2(new_n243), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n241), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n248), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n203), .B1(new_n240), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n260), .ZN(new_n262));
  INV_X1    g061(.A(new_n259), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n256), .B1(new_n257), .B2(new_n243), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n247), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n263), .A2(new_n266), .B1(new_n246), .B2(new_n247), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n215), .A2(new_n228), .A3(new_n226), .A4(new_n224), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n238), .B1(new_n268), .B2(new_n235), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n233), .A2(new_n236), .A3(KEYINPUT25), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n267), .A2(new_n271), .A3(KEYINPUT68), .A4(new_n221), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n261), .A2(new_n262), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT34), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n274), .B(KEYINPUT64), .Z(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT34), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(new_n273), .B2(new_n277), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT33), .B1(new_n273), .B2(new_n277), .ZN(new_n283));
  XNOR2_X1  g082(.A(G15gat), .B(G43gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G71gat), .ZN(new_n285));
  INV_X1    g084(.A(G99gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n282), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  AOI221_X4 g088(.A(new_n281), .B1(KEYINPUT33), .B2(new_n287), .C1(new_n273), .C2(new_n277), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n280), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n277), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT33), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n282), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n273), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n278), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n298), .A2(new_n276), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n288), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n291), .A2(KEYINPUT70), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT36), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n304), .B(new_n280), .C1(new_n289), .C2(new_n290), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT36), .A3(new_n301), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n291), .A2(new_n301), .A3(KEYINPUT69), .A4(KEYINPUT36), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n240), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n271), .A2(KEYINPUT75), .A3(new_n221), .ZN(new_n314));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n315), .B(KEYINPUT74), .Z(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT29), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n271), .A2(new_n316), .A3(new_n221), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT71), .B(G204gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(G197gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n322), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n325), .B1(new_n329), .B2(new_n322), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n320), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n314), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n316), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n329), .ZN(new_n340));
  INV_X1    g139(.A(new_n325), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT73), .A3(new_n330), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n240), .A2(new_n317), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n337), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n346), .A3(new_n354), .A4(new_n350), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n316), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n313), .B2(new_n314), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n359));
  INV_X1    g158(.A(new_n345), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n333), .B1(new_n318), .B2(new_n319), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n349), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT76), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n335), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n366), .A3(new_n349), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n365), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n350), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n356), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G141gat), .B(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(G155gat), .B2(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT78), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT2), .ZN(new_n380));
  OR2_X1    g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(KEYINPUT78), .A3(new_n376), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n264), .A2(new_n265), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(new_n241), .A3(new_n249), .A4(new_n258), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n385), .A2(new_n387), .A3(new_n388), .A4(new_n248), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n389), .A2(KEYINPUT80), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n387), .A3(new_n248), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT4), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n394), .A3(KEYINPUT4), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n385), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n383), .A2(KEYINPUT78), .A3(new_n376), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n376), .B1(new_n383), .B2(KEYINPUT78), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n378), .A2(KEYINPUT79), .A3(new_n384), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n260), .B(new_n397), .C1(new_n403), .C2(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n393), .A2(new_n395), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n391), .B1(new_n403), .B2(new_n267), .ZN(new_n408));
  INV_X1    g207(.A(new_n405), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n410), .B2(KEYINPUT5), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  AOI211_X1 g211(.A(KEYINPUT81), .B(new_n412), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n406), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n392), .A2(new_n389), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n404), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n422), .A2(KEYINPUT5), .A3(new_n409), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n414), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n410), .A2(new_n407), .A3(KEYINPUT5), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n260), .A2(new_n402), .A3(new_n401), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n405), .B1(new_n431), .B2(new_n391), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT81), .B1(new_n432), .B2(new_n412), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n404), .A2(new_n395), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n409), .B1(new_n390), .B2(new_n392), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n430), .A2(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n419), .B1(new_n436), .B2(new_n423), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n425), .A2(KEYINPUT83), .A3(new_n426), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT6), .B(new_n419), .C1(new_n436), .C2(new_n423), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n371), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT29), .B1(new_n385), .B2(new_n396), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n342), .B2(new_n330), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(KEYINPUT3), .ZN(new_n446));
  OAI221_X1 g245(.A(new_n443), .B1(new_n359), .B2(new_n444), .C1(new_n403), .C2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n385), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n334), .A2(new_n444), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n442), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G22gat), .B(G50gat), .Z(new_n451));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n447), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n447), .B2(new_n450), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n311), .B1(new_n441), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n405), .B1(new_n421), .B2(new_n404), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(KEYINPUT39), .C1(new_n409), .C2(new_n408), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n464), .A2(KEYINPUT85), .A3(new_n420), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT85), .B1(new_n464), .B2(new_n420), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT40), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n371), .A2(new_n437), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n471), .A2(new_n458), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n440), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n414), .A2(new_n424), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n419), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n344), .B1(new_n337), .B2(new_n345), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n318), .A2(new_n333), .A3(new_n319), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT37), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n335), .A2(new_n346), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT38), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .A4(new_n349), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n484), .A2(new_n352), .A3(new_n355), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n437), .A2(new_n425), .A3(new_n426), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(KEYINPUT87), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n474), .A3(new_n476), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n352), .A3(new_n355), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n369), .A2(new_n481), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n482), .A2(new_n349), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n459), .B1(new_n472), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n458), .A2(new_n291), .A3(new_n301), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT89), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n458), .A2(new_n291), .A3(new_n499), .A4(new_n301), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n441), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n302), .A2(new_n305), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n371), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n505));
  AND3_X1   g304(.A1(new_n489), .A2(new_n458), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n501), .A2(KEYINPUT35), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n202), .B1(new_n496), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n459), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n495), .A2(new_n472), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n439), .A2(new_n440), .ZN(new_n512));
  INV_X1    g311(.A(new_n371), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n500), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT35), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n504), .A2(new_n506), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(KEYINPUT90), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(G1gat), .ZN(new_n522));
  AOI21_X1  g321(.A(G8gat), .B1(new_n522), .B2(KEYINPUT94), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n524), .B2(G1gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n523), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT21), .ZN(new_n528));
  XOR2_X1   g327(.A(G71gat), .B(G78gat), .Z(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT96), .ZN(new_n530));
  XOR2_X1   g329(.A(G57gat), .B(G64gat), .Z(new_n531));
  INV_X1    g330(.A(KEYINPUT9), .ZN(new_n532));
  INV_X1    g331(.A(G71gat), .ZN(new_n533));
  INV_X1    g332(.A(G78gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G71gat), .B(G78gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n530), .A2(new_n531), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(KEYINPUT9), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n529), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n527), .B1(new_n528), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(new_n207), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n539), .A2(new_n541), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n544), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT20), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n548), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G211gat), .ZN(new_n553));
  AND2_X1   g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n548), .A2(new_n550), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(new_n550), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  OR2_X1    g365(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(G85gat), .A3(G92gat), .A4(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G106gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT8), .B1(new_n286), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n565), .A2(new_n566), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G99gat), .B(G106gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT101), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G43gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(G50gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(G50gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT15), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT93), .B(G50gat), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n580), .B1(new_n584), .B2(new_n579), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n585), .B2(KEYINPUT15), .ZN(new_n586));
  NAND2_X1  g385(.A1(G29gat), .A2(G36gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT92), .Z(new_n588));
  OAI21_X1  g387(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g389(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT91), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n590), .B1(new_n591), .B2(KEYINPUT91), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(KEYINPUT15), .A3(new_n582), .A4(new_n581), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n593), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n578), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT99), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n593), .A2(new_n597), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n601), .B(new_n605), .C1(new_n606), .C2(new_n578), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n610));
  XOR2_X1   g409(.A(G134gat), .B(G162gat), .Z(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n576), .A2(new_n545), .A3(new_n577), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n572), .A2(new_n574), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n542), .B1(new_n619), .B2(new_n575), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n618), .A2(new_n620), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n576), .A2(new_n545), .A3(KEYINPUT10), .A4(new_n577), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI211_X1 g432(.A(KEYINPUT102), .B(new_n622), .C1(new_n629), .C2(new_n630), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n623), .B(new_n627), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n623), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n626), .B1(new_n636), .B2(new_n631), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n561), .A2(new_n617), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n527), .B1(new_n599), .B2(new_n600), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n606), .A2(new_n527), .ZN(new_n641));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT18), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n606), .B(new_n527), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n642), .B(KEYINPUT13), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT18), .A4(new_n642), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G113gat), .B(G141gat), .ZN(new_n651));
  INV_X1    g450(.A(G197gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT11), .B(G169gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n645), .A2(new_n656), .A3(new_n648), .A4(new_n649), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n520), .A2(new_n639), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n512), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g465(.A1(new_n664), .A2(new_n513), .ZN(new_n667));
  NAND2_X1  g466(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n668));
  INV_X1    g467(.A(G8gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n524), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n673), .B(new_n674), .C1(new_n669), .C2(new_n667), .ZN(G1325gat));
  INV_X1    g474(.A(G15gat), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n664), .A2(new_n676), .A3(new_n311), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n664), .A2(new_n503), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n676), .B2(new_n678), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n458), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(new_n638), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n520), .A2(new_n617), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n561), .ZN(new_n685));
  INV_X1    g484(.A(new_n663), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n684), .A2(G29gat), .A3(new_n512), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n658), .A2(new_n660), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT103), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n638), .B(KEYINPUT104), .Z(new_n693));
  NAND3_X1  g492(.A1(new_n561), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n508), .A2(new_n617), .A3(new_n519), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT105), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n698), .A3(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n495), .A2(new_n472), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n459), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT106), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n518), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n617), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n705), .A2(KEYINPUT107), .A3(new_n706), .A4(new_n617), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n694), .B1(new_n700), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n512), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n690), .A2(new_n714), .ZN(G1328gat));
  OAI21_X1  g514(.A(G36gat), .B1(new_n713), .B2(new_n513), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n684), .A2(G36gat), .A3(new_n513), .A4(new_n688), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  NOR4_X1   g519(.A1(new_n684), .A2(G43gat), .A3(new_n503), .A4(new_n688), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(KEYINPUT108), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n579), .B1(new_n712), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n725), .B2(new_n721), .ZN(new_n726));
  INV_X1    g525(.A(new_n721), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n697), .A2(new_n699), .B1(new_n709), .B2(new_n710), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(new_n311), .A3(new_n694), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n727), .B(new_n722), .C1(new_n729), .C2(new_n579), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  INV_X1    g531(.A(new_n584), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n458), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n728), .A2(new_n694), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n684), .A2(new_n688), .ZN(new_n737));
  INV_X1    g536(.A(new_n458), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n584), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT109), .B(new_n732), .C1(new_n736), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n712), .A2(new_n734), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n732), .A2(KEYINPUT109), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n732), .A2(KEYINPUT109), .ZN(new_n743));
  INV_X1    g542(.A(new_n739), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n740), .A2(new_n745), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n561), .A2(new_n617), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n705), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n692), .A2(new_n693), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n512), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n371), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n756));
  INV_X1    g555(.A(G64gat), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT110), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  OR4_X1    g558(.A1(KEYINPUT110), .A2(new_n750), .A3(new_n513), .A4(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1333gat));
  NAND3_X1  g563(.A1(new_n748), .A2(G71gat), .A3(new_n749), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n765), .A2(KEYINPUT111), .A3(new_n311), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT111), .B1(new_n765), .B2(new_n311), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n502), .B(KEYINPUT112), .Z(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n533), .B1(new_n750), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n768), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n768), .B2(new_n771), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1334gat));
  NOR2_X1   g574(.A1(new_n750), .A2(new_n458), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT114), .B(G78gat), .Z(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n685), .A2(new_n692), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n638), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n700), .B2(new_n711), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n512), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n705), .A2(new_n617), .A3(new_n779), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(new_n563), .A3(new_n752), .A4(new_n638), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(G1336gat));
  AOI21_X1  g587(.A(new_n564), .B1(new_n781), .B2(new_n371), .ZN(new_n789));
  INV_X1    g588(.A(new_n693), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n786), .A2(new_n564), .A3(new_n371), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT52), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n728), .A2(new_n513), .A3(new_n780), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n794), .B(new_n791), .C1(new_n795), .C2(new_n564), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n782), .B2(new_n311), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n786), .A2(new_n286), .A3(new_n638), .A4(new_n502), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1338gat));
  AOI21_X1  g599(.A(new_n570), .B1(new_n781), .B2(new_n738), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n790), .A2(new_n570), .A3(new_n738), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT115), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n728), .A2(new_n458), .A3(new_n780), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n807), .B(new_n804), .C1(new_n808), .C2(new_n570), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1339gat));
  NAND3_X1  g609(.A1(new_n629), .A2(new_n622), .A3(new_n630), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT54), .B(new_n811), .C1(new_n633), .C2(new_n634), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n627), .B1(new_n631), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n635), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT116), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n635), .B(new_n820), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n692), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n646), .A2(new_n647), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n642), .B1(new_n640), .B2(new_n641), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n655), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n638), .A2(new_n660), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n617), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n660), .A2(new_n825), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n616), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n819), .A3(new_n821), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n561), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n561), .A2(new_n617), .A3(new_n692), .A4(new_n638), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n515), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n512), .A2(new_n371), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n242), .A3(new_n692), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n832), .A2(new_n834), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(new_n752), .A3(new_n458), .A4(new_n504), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n686), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(G1340gat));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n244), .A3(new_n638), .ZN(new_n843));
  OAI21_X1  g642(.A(G120gat), .B1(new_n840), .B2(new_n693), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n837), .B2(new_n685), .ZN(new_n846));
  INV_X1    g645(.A(G127gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n840), .A2(new_n847), .A3(new_n561), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n848), .ZN(G1342gat));
  INV_X1    g648(.A(G134gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n837), .A2(new_n850), .A3(new_n617), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT56), .Z(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n840), .B2(new_n616), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1343gat));
  AOI21_X1  g653(.A(new_n458), .B1(new_n832), .B2(new_n834), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n836), .A2(new_n311), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(G141gat), .A3(new_n686), .ZN(new_n858));
  INV_X1    g657(.A(new_n856), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n818), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n635), .B(KEYINPUT117), .C1(new_n816), .C2(new_n817), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n663), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n826), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n616), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n830), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n617), .B1(new_n865), .B2(new_n826), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n867), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n561), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n458), .B1(new_n872), .B2(new_n834), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT119), .B(new_n861), .C1(new_n873), .C2(new_n860), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n870), .A2(new_n867), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n831), .B1(new_n870), .B2(new_n867), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n833), .B1(new_n878), .B2(new_n561), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT57), .B1(new_n879), .B2(new_n458), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT119), .B1(new_n880), .B2(new_n861), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n692), .B1(new_n875), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n858), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n663), .A3(new_n861), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT58), .B1(new_n885), .B2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  INV_X1    g686(.A(new_n858), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n883), .A2(new_n884), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(new_n857), .ZN(new_n892));
  INV_X1    g691(.A(G148gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n638), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n861), .B1(new_n873), .B2(new_n860), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n683), .B1(new_n897), .B2(new_n874), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(KEYINPUT59), .A3(new_n893), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n855), .A2(new_n860), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n818), .A2(new_n616), .A3(new_n828), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n561), .B1(new_n870), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n639), .A2(new_n686), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT57), .B(new_n458), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n856), .B(KEYINPUT121), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n683), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n893), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n894), .B1(new_n899), .B2(new_n913), .ZN(G1345gat));
  NOR3_X1   g713(.A1(new_n857), .A2(G155gat), .A3(new_n561), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n561), .B1(new_n897), .B2(new_n874), .ZN(new_n917));
  INV_X1    g716(.A(G155gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n916), .C1(new_n917), .C2(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1346gat));
  AOI21_X1  g722(.A(G162gat), .B1(new_n892), .B2(new_n617), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n616), .B1(new_n897), .B2(new_n874), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n752), .A2(new_n513), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n839), .A2(new_n458), .A3(new_n769), .A4(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n686), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n835), .A2(new_n927), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n222), .A3(new_n692), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1348gat));
  NOR3_X1   g733(.A1(new_n930), .A2(new_n223), .A3(new_n693), .ZN(new_n935));
  AOI21_X1  g734(.A(G176gat), .B1(new_n932), .B2(new_n638), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  OAI21_X1  g736(.A(G183gat), .B1(new_n930), .B2(new_n561), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n932), .A2(new_n685), .A3(new_n204), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(KEYINPUT125), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  OAI221_X1 g741(.A(G190gat), .B1(KEYINPUT126), .B2(new_n942), .C1(new_n930), .C2(new_n616), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n208), .A3(new_n617), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G1351gat));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n311), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT127), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n905), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n686), .ZN(new_n952));
  AOI211_X1 g751(.A(new_n458), .B(new_n949), .C1(new_n832), .C2(new_n834), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n652), .A3(new_n692), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1352gat));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n956), .A3(new_n638), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n951), .B2(new_n693), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n953), .A2(new_n327), .A3(new_n685), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n905), .A2(new_n685), .A3(new_n950), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  OAI21_X1  g765(.A(G218gat), .B1(new_n951), .B2(new_n616), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n953), .A2(new_n328), .A3(new_n617), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1355gat));
endmodule


