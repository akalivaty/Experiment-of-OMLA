//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(new_n459), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n473), .B2(new_n459), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n462), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT69), .Z(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n473), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G136), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n471), .B2(new_n472), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n487), .B(new_n490), .C1(new_n472), .C2(new_n471), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n471), .B2(new_n472), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n459), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n500), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n492), .A2(new_n499), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(G75), .A2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(G651), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(KEYINPUT73), .B(G651), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(new_n516), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(G651), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(G651), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n523), .A2(new_n529), .A3(G88), .A4(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n529), .A2(G50), .A3(G543), .A4(new_n530), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n521), .A2(new_n522), .A3(new_n531), .A4(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND4_X1  g109(.A1(new_n523), .A2(new_n529), .A3(G89), .A4(new_n530), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n539), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n523), .A2(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n529), .A2(G51), .A3(G543), .A4(new_n530), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(G168));
  NAND4_X1  g119(.A1(new_n523), .A2(new_n529), .A3(G90), .A4(new_n530), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n529), .A2(G52), .A3(G543), .A4(new_n530), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n527), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n514), .B2(new_n516), .ZN(new_n551));
  AND2_X1   g126(.A1(G68), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT74), .B(G81), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n523), .A2(new_n529), .A3(new_n530), .A4(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n529), .A2(G43), .A3(G543), .A4(new_n530), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND4_X1  g138(.A1(new_n529), .A2(G53), .A3(G543), .A4(new_n530), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n529), .A2(new_n530), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n566), .A2(KEYINPUT75), .A3(G91), .A4(new_n523), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n523), .A2(new_n529), .A3(G91), .A4(new_n530), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n523), .A2(G65), .ZN(new_n572));
  INV_X1    g147(.A(G78), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n513), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n565), .A2(new_n571), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n543), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n535), .A2(new_n541), .A3(new_n542), .A4(KEYINPUT76), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G286));
  NAND3_X1  g156(.A1(new_n566), .A2(G87), .A3(new_n523), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n529), .A2(G543), .A3(new_n530), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(G288));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n514), .B2(new_n516), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n523), .A2(new_n529), .A3(G86), .A4(new_n530), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n529), .A2(G48), .A3(G543), .A4(new_n530), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  NAND3_X1  g170(.A1(new_n566), .A2(G85), .A3(new_n523), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n583), .A2(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(new_n527), .C2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n566), .A2(KEYINPUT10), .A3(G92), .A4(new_n523), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n523), .A2(new_n529), .A3(G92), .A4(new_n530), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n514), .B2(new_n516), .ZN(new_n607));
  AND2_X1   g182(.A1(G79), .A2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT78), .B1(new_n607), .B2(new_n608), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n611), .A2(G651), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n583), .A2(G54), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n605), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G286), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G299), .B(KEYINPUT79), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G297));
  AOI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n557), .A2(new_n619), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n615), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n462), .A2(new_n460), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT13), .Z(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2100), .ZN(new_n635));
  INV_X1    g210(.A(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n459), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI22_X1  g213(.A1(new_n463), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(G123), .B2(new_n476), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n634), .A2(new_n635), .A3(new_n642), .A4(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n661), .B(KEYINPUT17), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n663), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n663), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n662), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g250(.A(KEYINPUT82), .B(new_n672), .C1(new_n668), .C2(new_n662), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n669), .C2(new_n670), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n666), .B(new_n671), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2096), .B(G2100), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1956), .B(G2474), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n691), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(new_n689), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT84), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n693), .B(KEYINPUT20), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G1981), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n700), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n700), .B2(new_n704), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n686), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n700), .A2(new_n704), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G1981), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n700), .A2(new_n704), .A3(new_n705), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(G1986), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT85), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n708), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n708), .B2(new_n712), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n685), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n706), .A2(new_n707), .A3(new_n686), .ZN(new_n719));
  AOI21_X1  g294(.A(G1986), .B1(new_n710), .B2(new_n711), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n708), .A2(new_n712), .A3(new_n715), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n721), .A2(new_n684), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n718), .A2(new_n723), .ZN(G229));
  NAND2_X1  g299(.A1(new_n616), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G4), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1348), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G19), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n558), .B2(new_n730), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1341), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G26), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G140), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n459), .A2(G116), .ZN(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n463), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G128), .B2(new_n476), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n737), .B1(new_n742), .B2(new_n735), .ZN(new_n743));
  INV_X1    g318(.A(G2067), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n728), .A2(new_n729), .A3(new_n733), .A4(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT90), .Z(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  INV_X1    g323(.A(G127), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n473), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n459), .B1(new_n750), .B2(KEYINPUT92), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(KEYINPUT92), .B2(new_n750), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G139), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n463), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n752), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2072), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n730), .A2(G20), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G299), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n735), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n735), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT29), .B(G2090), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n730), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n730), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(G1966), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n730), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n730), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n781), .B(new_n782), .C1(G1961), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n735), .A2(G32), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n476), .A2(G129), .ZN(new_n787));
  NAND3_X1  g362(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT26), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n460), .A2(G105), .ZN(new_n790));
  INV_X1    g365(.A(G141), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n789), .B(new_n790), .C1(new_n463), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n786), .B1(new_n793), .B2(new_n735), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n735), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n735), .ZN(new_n798));
  INV_X1    g373(.A(G2078), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(KEYINPUT24), .A2(G34), .ZN(new_n802));
  NOR2_X1   g377(.A1(KEYINPUT24), .A2(G34), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n735), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT94), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G160), .B2(G29), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G2084), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n784), .A2(G1961), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(G2084), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT95), .B(G28), .Z(new_n811));
  AOI21_X1  g386(.A(G29), .B1(new_n811), .B2(KEYINPUT30), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(KEYINPUT30), .B2(new_n811), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT31), .B(G11), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G29), .B2(new_n640), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n778), .A2(new_n785), .A3(new_n801), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n747), .A2(new_n774), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n730), .A2(G23), .ZN(new_n820));
  INV_X1    g395(.A(G288), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n730), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT33), .B(G1976), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n730), .A2(G22), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n730), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1971), .ZN(new_n827));
  MUX2_X1   g402(.A(G6), .B(G305), .S(G16), .Z(new_n828));
  XOR2_X1   g403(.A(KEYINPUT32), .B(G1981), .Z(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT86), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  OR3_X1    g406(.A1(new_n824), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n735), .A2(G25), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n476), .A2(G119), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n837));
  INV_X1    g412(.A(G107), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(G2105), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n482), .B2(G131), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n835), .B1(new_n841), .B2(new_n735), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n842), .B(new_n844), .ZN(new_n845));
  MUX2_X1   g420(.A(G24), .B(G290), .S(G16), .Z(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(G1986), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(G1986), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n833), .A2(new_n834), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT87), .B1(new_n850), .B2(KEYINPUT36), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(KEYINPUT87), .A3(KEYINPUT36), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n833), .A2(new_n855), .A3(new_n834), .A4(new_n849), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT88), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n819), .B1(new_n854), .B2(new_n858), .ZN(G311));
  INV_X1    g434(.A(new_n819), .ZN(new_n860));
  INV_X1    g435(.A(new_n853), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n851), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n856), .B(KEYINPUT88), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(G150));
  NAND2_X1  g439(.A1(new_n616), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  INV_X1    g441(.A(G67), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n514), .B2(new_n516), .ZN(new_n868));
  AND2_X1   g443(.A1(G80), .A2(G543), .ZN(new_n869));
  OAI21_X1  g444(.A(G651), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(KEYINPUT97), .B(G93), .Z(new_n871));
  NAND4_X1  g446(.A1(new_n523), .A2(new_n871), .A3(new_n529), .A4(new_n530), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n529), .A2(G55), .A3(G543), .A4(new_n530), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n557), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n557), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n866), .B(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n880), .A2(new_n881), .A3(G860), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n874), .A2(G860), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT37), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n882), .A2(new_n884), .ZN(G145));
  NOR2_X1   g460(.A1(new_n504), .A2(new_n507), .ZN(new_n886));
  INV_X1    g461(.A(new_n491), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n490), .B1(new_n462), .B2(new_n487), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n742), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n742), .A2(new_n889), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n793), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n793), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n764), .B(new_n763), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n761), .A3(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n836), .A2(new_n840), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n459), .A2(G118), .ZN(new_n899));
  OAI21_X1  g474(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n482), .A2(G142), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G130), .ZN(new_n903));
  INV_X1    g478(.A(new_n476), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n898), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n904), .B2(new_n903), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n841), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n632), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n907), .A3(new_n632), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n895), .A2(new_n897), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n640), .B(G160), .Z(new_n914));
  XNOR2_X1  g489(.A(new_n484), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n895), .A2(new_n912), .A3(new_n897), .ZN(new_n918));
  INV_X1    g493(.A(new_n911), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n895), .A2(new_n897), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT98), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n925));
  INV_X1    g500(.A(new_n910), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n908), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n895), .A2(new_n927), .A3(new_n897), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n915), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n897), .B2(new_n895), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n923), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(G395));
  NAND2_X1  g509(.A1(new_n874), .A2(new_n619), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(G288), .B(G305), .Z(new_n937));
  XNOR2_X1  g512(.A(G290), .B(G303), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n627), .A2(new_n877), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n876), .B(new_n875), .C1(new_n615), .C2(G559), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G299), .A2(new_n615), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n527), .B1(new_n609), .B2(new_n610), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n945), .A2(new_n612), .B1(G54), .B2(new_n583), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n567), .A2(new_n570), .B1(G651), .B2(new_n574), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n565), .A4(new_n605), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n944), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT41), .B1(new_n944), .B2(new_n948), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n953), .B1(new_n952), .B2(new_n956), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n940), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n959), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n939), .A3(new_n957), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n936), .B1(new_n963), .B2(G868), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT101), .ZN(G295));
  XNOR2_X1  g540(.A(new_n964), .B(KEYINPUT102), .ZN(G331));
  INV_X1    g541(.A(KEYINPUT41), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n949), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n944), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n969));
  AOI21_X1  g544(.A(G301), .B1(new_n578), .B2(new_n579), .ZN(new_n970));
  NOR2_X1   g545(.A1(G171), .A2(G168), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n876), .B(new_n875), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n877), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n968), .A2(new_n969), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n950), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT103), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n954), .A2(new_n955), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n974), .A2(new_n972), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n939), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n975), .A2(KEYINPUT103), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n949), .B1(new_n974), .B2(new_n972), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n980), .B2(new_n981), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n940), .B(new_n984), .C1(new_n986), .C2(KEYINPUT103), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n987), .A3(new_n924), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n975), .A2(new_n977), .ZN(new_n991));
  AOI21_X1  g566(.A(G37), .B1(new_n991), .B2(new_n939), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n987), .A2(KEYINPUT104), .A3(new_n992), .A4(new_n990), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n988), .A2(new_n990), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n987), .A2(KEYINPUT43), .A3(new_n992), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT44), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(KEYINPUT126), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n742), .B(new_n744), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n889), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n466), .A2(new_n467), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G2105), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n482), .A2(G137), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(G40), .A4(new_n461), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT105), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1005), .A2(KEYINPUT105), .A3(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n793), .B(new_n1017), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n1015), .B(new_n1016), .C1(new_n1014), .C2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n898), .A2(new_n844), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n742), .A2(new_n744), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(KEYINPUT125), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1014), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT125), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1004), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n793), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1014), .B1(new_n1005), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1014), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1029), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1028), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT47), .Z(new_n1034));
  NOR2_X1   g609(.A1(new_n841), .A2(new_n843), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1014), .B1(new_n1035), .B2(new_n1020), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1019), .A2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1029), .A2(G1986), .A3(G290), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1038), .B(KEYINPUT48), .Z(new_n1039));
  AOI21_X1  g614(.A(new_n1034), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1026), .A2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1024), .A2(new_n1004), .A3(new_n1025), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT107), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n496), .A2(new_n498), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n489), .B2(new_n491), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(G1384), .ZN(new_n1047));
  INV_X1    g622(.A(G40), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n465), .A2(new_n468), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n889), .A2(KEYINPUT107), .A3(new_n1006), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n582), .A2(new_n584), .A3(G1976), .A4(new_n585), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(G8), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n593), .A2(new_n594), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT5), .B1(new_n515), .B2(G543), .ZN(new_n1057));
  OAI21_X1  g632(.A(G61), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n589), .B(KEYINPUT77), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n527), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(G1981), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT110), .B(G1981), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(KEYINPUT49), .A3(new_n1063), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(G8), .A3(new_n1051), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1070), .A2(new_n1051), .A3(G8), .A4(new_n1052), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1054), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1054), .A2(new_n1068), .A3(KEYINPUT111), .A4(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT108), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G303), .A2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(G303), .A2(KEYINPUT108), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT106), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1384), .B1(new_n492), .B2(new_n886), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT106), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(KEYINPUT45), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n509), .A2(new_n1006), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1013), .B1(new_n1090), .B2(new_n1008), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1971), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1013), .B1(new_n1090), .B2(KEYINPUT50), .ZN(new_n1093));
  INV_X1    g668(.A(G2090), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1047), .A2(new_n1095), .A3(new_n1050), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1084), .B(G8), .C1(new_n1092), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT109), .ZN(new_n1099));
  INV_X1    g674(.A(G1971), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1087), .B1(new_n1086), .B2(KEYINPUT45), .ZN(new_n1101));
  NOR4_X1   g676(.A1(new_n1046), .A2(KEYINPUT106), .A3(new_n1008), .A4(G1384), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n489), .A2(new_n491), .B1(new_n1045), .B2(new_n500), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1384), .B1(new_n1104), .B2(new_n499), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1049), .B1(new_n1105), .B2(KEYINPUT45), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1100), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(G8), .A4(new_n1084), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1076), .A2(new_n1099), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1068), .A2(new_n1069), .A3(new_n821), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1063), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(G8), .A3(new_n1051), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1099), .A2(new_n1111), .ZN(new_n1117));
  OAI21_X1  g692(.A(G8), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT114), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1084), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1109), .A2(new_n1121), .A3(G8), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n580), .A2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(G1966), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT45), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1049), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT113), .B(G2084), .Z(new_n1130));
  NAND3_X1  g705(.A1(new_n1093), .A2(new_n1096), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1124), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1117), .A2(new_n1123), .A3(new_n1132), .A4(new_n1076), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1116), .B1(KEYINPUT63), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT112), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1072), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1054), .A2(new_n1068), .A3(KEYINPUT112), .A4(new_n1071), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1049), .B1(new_n1090), .B2(KEYINPUT50), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1095), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1139), .A2(new_n1140), .A3(G2090), .ZN(new_n1141));
  OAI21_X1  g716(.A(G8), .B1(new_n1141), .B2(new_n1092), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1120), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1117), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1089), .A2(new_n799), .A3(new_n1091), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1146));
  INV_X1    g721(.A(G1961), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1145), .A2(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n1150));
  OR3_X1    g725(.A1(new_n1126), .A2(new_n1128), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(G301), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1129), .A2(G168), .A3(new_n1131), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G8), .ZN(new_n1154));
  AOI21_X1  g729(.A(G168), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT51), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT51), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(new_n1157), .A3(G8), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT62), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1156), .A2(new_n1161), .A3(new_n1158), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1144), .A2(new_n1152), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1144), .A2(new_n1164), .A3(new_n1132), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1134), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT118), .B(KEYINPUT61), .Z(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT56), .B(G2072), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1089), .A2(KEYINPUT115), .A3(new_n1091), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n772), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(G299), .B(KEYINPUT57), .Z(new_n1172));
  NAND3_X1  g747(.A1(new_n1089), .A2(new_n1091), .A3(new_n1168), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT115), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1172), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1167), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1176), .B1(new_n1178), .B2(KEYINPUT120), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1171), .A2(new_n1182), .A3(new_n1172), .A4(new_n1175), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1181), .A2(new_n1183), .A3(KEYINPUT61), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1051), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1148), .A2(new_n727), .B1(new_n1185), .B2(new_n744), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1186), .A2(new_n1187), .A3(new_n616), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1189));
  XNOR2_X1  g764(.A(KEYINPUT116), .B(G1996), .ZN(new_n1190));
  XNOR2_X1  g765(.A(KEYINPUT58), .B(G1341), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1189), .A2(new_n1190), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT59), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n558), .A2(KEYINPUT117), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1188), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1186), .A2(new_n615), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1186), .A2(new_n615), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1187), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT119), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1202), .B(new_n1167), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1180), .A2(new_n1184), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1198), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1178), .B1(new_n1205), .B2(new_n1176), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(G301), .B(KEYINPUT54), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1148), .A2(new_n1147), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(KEYINPUT123), .B(G2078), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1089), .A2(KEYINPUT53), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1009), .A2(KEYINPUT122), .A3(new_n1049), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1086), .A2(KEYINPUT45), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1216), .B1(new_n1217), .B2(new_n1013), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1214), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1209), .B1(new_n1212), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1149), .A2(new_n1208), .A3(new_n1151), .ZN(new_n1221));
  AOI22_X1  g796(.A1(new_n1156), .A2(new_n1158), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g797(.A(KEYINPUT124), .B1(new_n1144), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1159), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1117), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n1227));
  NOR3_X1   g802(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n1223), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1166), .B1(new_n1207), .B2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g805(.A(G290), .B(new_n686), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1037), .B1(new_n1029), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1043), .B1(new_n1230), .B2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g808(.A(G319), .B1(new_n658), .B2(new_n659), .ZN(new_n1235));
  NOR2_X1   g809(.A1(G227), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g810(.A1(new_n718), .A2(new_n723), .A3(new_n1236), .ZN(new_n1237));
  NOR2_X1   g811(.A1(new_n1237), .A2(new_n932), .ZN(new_n1238));
  AND3_X1   g812(.A1(new_n997), .A2(new_n1238), .A3(KEYINPUT127), .ZN(new_n1239));
  AOI21_X1  g813(.A(KEYINPUT127), .B1(new_n997), .B2(new_n1238), .ZN(new_n1240));
  NOR2_X1   g814(.A1(new_n1239), .A2(new_n1240), .ZN(G308));
  NAND2_X1  g815(.A1(new_n997), .A2(new_n1238), .ZN(G225));
endmodule


