//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(G148gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT78), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT78), .B1(new_n221), .B2(new_n209), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n214), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT79), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n217), .B1(new_n215), .B2(new_n216), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(KEYINPUT78), .A3(new_n209), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n214), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n210), .B(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(G141gat), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n212), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(new_n209), .B2(new_n221), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n224), .A2(new_n229), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT84), .ZN(new_n238));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT1), .ZN(new_n241));
  XOR2_X1   g040(.A(G113gat), .B(G120gat), .Z(new_n242));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n237), .A2(new_n238), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n236), .A2(new_n231), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n227), .A2(new_n228), .A3(new_n214), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n228), .B1(new_n227), .B2(new_n214), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n246), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT84), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n247), .B(new_n252), .C1(new_n237), .C2(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n208), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT82), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n224), .A2(new_n229), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n258), .A4(new_n248), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n248), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n246), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n255), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT4), .B1(new_n247), .B2(new_n252), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n251), .A2(KEYINPUT4), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n251), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n267), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT85), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n267), .B(new_n276), .C1(new_n268), .C2(new_n273), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n257), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT4), .B1(new_n237), .B2(new_n246), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n247), .A2(new_n252), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(KEYINPUT4), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(new_n267), .A3(new_n208), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n207), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n277), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n251), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT83), .B1(new_n251), .B2(KEYINPUT4), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n238), .B1(new_n237), .B2(new_n246), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n251), .A2(KEYINPUT84), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n276), .B1(new_n293), .B2(new_n267), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n256), .B1(new_n285), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n206), .A3(new_n282), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n284), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT91), .ZN(new_n299));
  XOR2_X1   g098(.A(G8gat), .B(G36gat), .Z(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  AND2_X1   g102(.A1(G211gat), .A2(G218gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(KEYINPUT22), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G211gat), .A2(G218gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n305), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT26), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR3_X1   g113(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(KEYINPUT27), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G183gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n322), .A3(new_n317), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(KEYINPUT68), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n323), .B2(KEYINPUT68), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n319), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT64), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT65), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n311), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(new_n312), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g140(.A(KEYINPUT66), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT25), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n311), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n341), .B2(new_n342), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n334), .B1(G183gat), .B2(G190gat), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(new_n329), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n328), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n354), .B(KEYINPUT75), .Z(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n329), .B(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n343), .B1(new_n358), .B2(new_n335), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n359), .A2(new_n360), .B1(new_n351), .B2(new_n349), .ZN(new_n361));
  INV_X1    g160(.A(new_n327), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n318), .B1(new_n362), .B2(new_n325), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(KEYINPUT29), .ZN(new_n365));
  INV_X1    g164(.A(new_n354), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n310), .B(new_n356), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n310), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n355), .B1(new_n353), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n364), .A2(new_n354), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT37), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT93), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n302), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n367), .A2(new_n372), .A3(KEYINPUT93), .A4(new_n373), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n367), .A2(new_n372), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT76), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n367), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n373), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT38), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(KEYINPUT6), .B(new_n207), .C1(new_n278), .C2(new_n283), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n372), .A3(new_n302), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n353), .A2(new_n366), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n310), .C1(new_n365), .C2(new_n355), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT92), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n370), .A2(new_n371), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n310), .ZN(new_n394));
  INV_X1    g193(.A(new_n365), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(new_n354), .B1(new_n355), .B2(new_n353), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n391), .B(new_n394), .C1(new_n310), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT37), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT38), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n388), .B1(new_n400), .B2(new_n378), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT38), .B1(new_n397), .B2(KEYINPUT37), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(KEYINPUT94), .A3(new_n377), .A4(new_n376), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n284), .A2(new_n296), .A3(new_n405), .A4(new_n297), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n299), .A2(new_n387), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT40), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n264), .A2(new_n266), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n254), .B1(new_n281), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT39), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n207), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT90), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT90), .B(KEYINPUT39), .C1(new_n253), .C2(new_n255), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n408), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n386), .A2(KEYINPUT77), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT30), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n386), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n380), .A2(new_n382), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n419), .B(new_n421), .C1(new_n422), .C2(new_n302), .ZN(new_n423));
  OAI221_X1 g222(.A(KEYINPUT40), .B1(new_n410), .B2(new_n415), .C1(new_n412), .C2(new_n413), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n417), .A2(new_n423), .A3(new_n284), .A4(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  INV_X1    g225(.A(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n264), .A2(new_n369), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n368), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n260), .B2(new_n263), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT89), .B1(new_n435), .B2(new_n310), .ZN(new_n436));
  INV_X1    g235(.A(G228gat), .ZN(new_n437));
  INV_X1    g236(.A(G233gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n258), .B1(new_n309), .B2(KEYINPUT29), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n265), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n435), .A2(new_n310), .ZN(new_n442));
  INV_X1    g241(.A(new_n307), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT29), .B1(new_n305), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n443), .B2(new_n305), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT3), .B1(new_n445), .B2(new_n446), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n237), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n442), .A2(new_n449), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n441), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n441), .B2(new_n450), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n431), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n441), .A2(new_n450), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G22gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n452), .A3(new_n430), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n425), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n407), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g262(.A(new_n246), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n361), .B2(new_n363), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n328), .B(new_n246), .C1(new_n344), .C2(new_n352), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G227gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n438), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n463), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  AOI211_X1 g270(.A(KEYINPUT70), .B(new_n471), .C1(new_n465), .C2(new_n466), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT32), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT33), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n470), .B2(new_n472), .ZN(new_n475));
  XOR2_X1   g274(.A(G15gat), .B(G43gat), .Z(new_n476));
  XNOR2_X1  g275(.A(G71gat), .B(G99gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  OAI221_X1 g279(.A(KEYINPUT32), .B1(new_n474), .B2(new_n480), .C1(new_n470), .C2(new_n472), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n471), .A3(new_n466), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n483), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT71), .B1(new_n483), .B2(KEYINPUT34), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n483), .A2(KEYINPUT34), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n481), .A3(new_n487), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT36), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT72), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n482), .B2(new_n492), .ZN(new_n493));
  AOI211_X1 g292(.A(KEYINPUT72), .B(new_n487), .C1(new_n479), .C2(new_n481), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(KEYINPUT36), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n298), .A2(new_n385), .ZN(new_n497));
  INV_X1    g296(.A(new_n423), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n499), .B2(new_n459), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n497), .A2(new_n460), .A3(new_n498), .A4(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n299), .A2(new_n385), .A3(new_n406), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n455), .A2(new_n458), .A3(new_n489), .A4(new_n490), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n504), .A2(KEYINPUT35), .A3(new_n423), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n462), .A2(new_n500), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G43gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n427), .A2(G43gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT15), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT97), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT15), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n513), .B(new_n514), .C1(KEYINPUT97), .C2(new_n510), .ZN(new_n515));
  INV_X1    g314(.A(G36gat), .ZN(new_n516));
  AND2_X1   g315(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n512), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n512), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT17), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT17), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(G1gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  INV_X1    g330(.A(G1gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT16), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n531), .B1(new_n530), .B2(new_n534), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n526), .A2(new_n527), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n523), .A2(new_n525), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT18), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n540), .B(new_n541), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n539), .B(KEYINPUT13), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n545), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n538), .A2(new_n539), .A3(new_n542), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n553));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT95), .B(KEYINPUT11), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G169gat), .B(G197gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT12), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n552), .A2(new_n553), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n552), .B2(new_n553), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT101), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G155gat), .ZN(new_n566));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT99), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g371(.A1(KEYINPUT99), .A2(G71gat), .A3(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G57gat), .B(G64gat), .Z(new_n577));
  INV_X1    g376(.A(new_n570), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(KEYINPUT9), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n579), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G127gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n540), .B1(new_n583), .B2(KEYINPUT21), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(G127gat), .B1(new_n586), .B2(new_n587), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n592), .B1(new_n590), .B2(new_n593), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n569), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n593), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n591), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n594), .A3(new_n568), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n526), .A2(new_n527), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT105), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT104), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n609), .A2(KEYINPUT8), .ZN(new_n610));
  NOR2_X1   g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G85gat), .ZN(new_n613));
  INV_X1    g412(.A(G92gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT103), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n607), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G99gat), .B(G106gat), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n618), .B(new_n607), .C1(new_n616), .C2(new_n612), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n604), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n604), .B1(new_n617), .B2(new_n619), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n603), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n605), .B(new_n606), .Z(new_n626));
  NOR3_X1   g425(.A1(new_n610), .A2(new_n608), .A3(new_n611), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n615), .A2(KEYINPUT103), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n618), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n617), .A2(new_n619), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT104), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n632), .A2(KEYINPUT105), .A3(new_n623), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n602), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT105), .B1(new_n632), .B2(new_n623), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n603), .A3(new_n624), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n541), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n634), .A2(new_n636), .A3(new_n637), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT106), .ZN(new_n642));
  XNOR2_X1  g441(.A(G134gat), .B(G162gat), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT107), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n634), .A2(new_n637), .A3(new_n640), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n635), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n641), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n642), .A2(new_n652), .A3(new_n645), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n647), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n642), .B2(new_n645), .ZN(new_n655));
  INV_X1    g454(.A(new_n645), .ZN(new_n656));
  AOI211_X1 g455(.A(KEYINPUT107), .B(new_n656), .C1(new_n641), .C2(KEYINPUT106), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n650), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT10), .A4(new_n583), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n620), .A2(new_n621), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n583), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n630), .A2(new_n631), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n623), .B1(new_n665), .B2(new_n604), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n663), .B(new_n664), .C1(new_n666), .C2(new_n583), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n660), .B1(new_n661), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n663), .B1(new_n666), .B2(new_n583), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(new_n660), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT108), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n674), .B(new_n668), .C1(new_n669), .C2(new_n660), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n601), .A2(new_n654), .A3(new_n658), .A4(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n507), .A2(new_n563), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n497), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n423), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT109), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT16), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G8gat), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n680), .A2(new_n531), .A3(new_n423), .A4(new_n687), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n684), .A2(new_n685), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(G1325gat));
  INV_X1    g491(.A(new_n680), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n482), .A2(new_n492), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n487), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n482), .A2(new_n492), .A3(new_n488), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(KEYINPUT36), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT36), .ZN(new_n698));
  INV_X1    g497(.A(new_n490), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n487), .B1(new_n479), .B2(new_n481), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n693), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(G15gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n680), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(G1326gat));
  NAND2_X1  g506(.A1(new_n680), .A2(new_n459), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  AND2_X1   g509(.A1(new_n654), .A2(new_n658), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n462), .A2(new_n500), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n502), .A2(new_n506), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n678), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n601), .A3(new_n563), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n520), .A3(new_n681), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n507), .B2(new_n711), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n654), .A2(new_n658), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n423), .B1(new_n298), .B2(new_n385), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n702), .B1(new_n724), .B2(new_n460), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n407), .B2(new_n461), .ZN(new_n726));
  AOI22_X1  g525(.A1(KEYINPUT35), .A2(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT44), .B(new_n723), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n681), .A3(new_n716), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G29gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n720), .A2(new_n731), .ZN(G1328gat));
  NAND4_X1  g531(.A1(new_n722), .A2(new_n423), .A3(new_n728), .A4(new_n716), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G36gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  AOI21_X1  g534(.A(G36gat), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n423), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n717), .A2(new_n738), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n735), .A2(KEYINPUT46), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n718), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n734), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n734), .A2(new_n741), .A3(KEYINPUT111), .A4(new_n739), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1329gat));
  NAND4_X1  g545(.A1(new_n722), .A2(new_n496), .A3(new_n728), .A4(new_n716), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G43gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n718), .A2(new_n508), .A3(new_n705), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(KEYINPUT47), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1330gat));
  NAND4_X1  g553(.A1(new_n722), .A2(new_n459), .A3(new_n728), .A4(new_n716), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G50gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT112), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n718), .A2(new_n427), .A3(new_n459), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n756), .B(new_n758), .C1(KEYINPUT112), .C2(KEYINPUT48), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n712), .A2(new_n713), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765));
  INV_X1    g564(.A(new_n601), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n723), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n678), .A2(new_n562), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n764), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT113), .B1(new_n507), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n681), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g574(.A(KEYINPUT49), .B(G64gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n423), .A3(new_n776), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n772), .A2(new_n498), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1333gat));
  OAI21_X1  g578(.A(G71gat), .B1(new_n772), .B2(new_n702), .ZN(new_n780));
  INV_X1    g579(.A(G71gat), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n769), .A2(new_n771), .A3(new_n781), .A4(new_n705), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n780), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n773), .A2(new_n459), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT115), .B(G78gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n601), .A2(new_n562), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n790), .B(new_n723), .C1(new_n726), .C2(new_n727), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n714), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(KEYINPUT116), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n681), .A2(new_n613), .A3(new_n715), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n601), .A2(new_n562), .A3(new_n678), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n729), .A2(new_n681), .A3(new_n801), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n799), .A2(new_n800), .B1(new_n613), .B2(new_n802), .ZN(G1336gat));
  NAND3_X1  g602(.A1(new_n715), .A2(new_n423), .A3(new_n614), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n797), .B2(new_n798), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n722), .A2(new_n423), .A3(new_n728), .A4(new_n801), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G92gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n804), .B(KEYINPUT117), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n795), .A2(new_n810), .B1(new_n806), .B2(G92gat), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n805), .A2(new_n809), .B1(new_n808), .B2(new_n811), .ZN(G1337gat));
  INV_X1    g611(.A(G99gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n715), .A2(new_n705), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n729), .A2(new_n496), .A3(new_n801), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n799), .A2(new_n814), .B1(new_n813), .B2(new_n815), .ZN(G1338gat));
  NOR3_X1   g615(.A1(new_n460), .A2(G106gat), .A3(new_n678), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n797), .B2(new_n798), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n722), .A2(new_n459), .A3(new_n728), .A4(new_n801), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n795), .A2(new_n817), .B1(new_n820), .B2(G106gat), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n819), .A2(new_n823), .B1(new_n822), .B2(new_n824), .ZN(G1339gat));
  NOR2_X1   g624(.A1(new_n679), .A2(new_n562), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n661), .A2(new_n667), .A3(new_n660), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n828), .A2(new_n668), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n661), .A2(new_n667), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n829), .A3(new_n659), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n674), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n670), .A2(new_n675), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n659), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n661), .A2(new_n667), .A3(new_n660), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n675), .B1(new_n668), .B2(new_n829), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n834), .A2(new_n562), .A3(new_n835), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n539), .B1(new_n538), .B2(new_n542), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT118), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(KEYINPUT118), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n843), .B(new_n844), .C1(new_n547), .C2(new_n548), .ZN(new_n845));
  INV_X1    g644(.A(new_n552), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n845), .A2(new_n558), .B1(new_n846), .B2(new_n559), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n676), .B2(new_n677), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n711), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n834), .A2(new_n835), .A3(new_n840), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n723), .A2(new_n851), .A3(new_n847), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n826), .B1(new_n853), .B2(new_n766), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n497), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n460), .A3(new_n498), .A4(new_n705), .ZN(new_n856));
  INV_X1    g655(.A(G113gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n856), .A2(new_n857), .A3(new_n563), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n459), .A2(new_n493), .A3(new_n494), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n601), .B1(new_n850), .B2(new_n852), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n681), .B(new_n859), .C1(new_n860), .C2(new_n826), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n423), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n562), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n858), .A2(new_n863), .ZN(G1340gat));
  INV_X1    g663(.A(G120gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n856), .A2(new_n865), .A3(new_n678), .ZN(new_n866));
  AOI21_X1  g665(.A(G120gat), .B1(new_n862), .B2(new_n715), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(G1341gat));
  NOR3_X1   g667(.A1(new_n861), .A2(new_n423), .A3(new_n766), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n589), .B1(new_n869), .B2(KEYINPUT119), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n601), .A2(G127gat), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n870), .A2(new_n871), .B1(new_n856), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT120), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  OAI221_X1 g674(.A(new_n875), .B1(new_n856), .B2(new_n872), .C1(new_n870), .C2(new_n871), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1342gat));
  OAI21_X1  g676(.A(G134gat), .B1(new_n856), .B2(new_n711), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n711), .A2(G134gat), .A3(new_n423), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n861), .A2(KEYINPUT56), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT56), .B1(new_n861), .B2(new_n879), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  OAI21_X1  g681(.A(KEYINPUT57), .B1(new_n854), .B2(new_n460), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(new_n459), .C1(new_n860), .C2(new_n826), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n496), .A2(new_n497), .A3(new_n423), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(G141gat), .A3(new_n562), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n496), .A2(new_n460), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n855), .A2(new_n498), .A3(new_n562), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n211), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(G1344gat));
  AND3_X1   g693(.A1(new_n715), .A2(new_n232), .A3(new_n233), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n855), .A2(new_n498), .A3(new_n889), .A4(new_n895), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT121), .Z(new_n897));
  NAND4_X1  g696(.A1(new_n883), .A2(new_n715), .A3(new_n885), .A4(new_n887), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT59), .B1(new_n232), .B2(new_n233), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(KEYINPUT122), .A3(new_n899), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n898), .B2(G148gat), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n904), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(G1345gat));
  NAND2_X1  g708(.A1(new_n855), .A2(new_n889), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(new_n219), .A3(new_n498), .A4(new_n601), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n886), .A2(new_n601), .A3(new_n887), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n219), .ZN(G1346gat));
  NAND4_X1  g713(.A1(new_n911), .A2(new_n220), .A3(new_n498), .A4(new_n723), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n886), .A2(new_n723), .A3(new_n887), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G162gat), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n854), .A2(new_n681), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n504), .A2(new_n498), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(G169gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(new_n563), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n859), .A2(new_n423), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n562), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n925), .B2(new_n930), .ZN(G1348gat));
  INV_X1    g730(.A(G176gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n924), .A2(new_n932), .A3(new_n678), .ZN(new_n933));
  AOI21_X1  g732(.A(G176gat), .B1(new_n929), .B2(new_n715), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1349gat));
  OAI21_X1  g736(.A(G183gat), .B1(new_n924), .B2(new_n766), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n601), .A2(new_n320), .A3(new_n322), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n928), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n929), .A2(new_n317), .A3(new_n723), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n922), .A2(new_n723), .A3(new_n923), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n945), .A3(G190gat), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n945), .B1(new_n944), .B2(G190gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  XNOR2_X1  g748(.A(KEYINPUT127), .B(G197gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n496), .A2(new_n681), .A3(new_n498), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n886), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n563), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n922), .A2(new_n423), .A3(new_n889), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n563), .A2(new_n950), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(G1352gat));
  OAI21_X1  g755(.A(G204gat), .B1(new_n952), .B2(new_n678), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n678), .A2(G204gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT62), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n954), .A2(KEYINPUT62), .A3(new_n959), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  OR3_X1    g761(.A1(new_n954), .A2(G211gat), .A3(new_n766), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n886), .A2(new_n601), .A3(new_n951), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  OAI21_X1  g766(.A(G218gat), .B1(new_n952), .B2(new_n711), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n711), .A2(G218gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n954), .B2(new_n969), .ZN(G1355gat));
endmodule


