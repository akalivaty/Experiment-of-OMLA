//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(new_n454), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n470), .A2(new_n471), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n463), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND2_X1  g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n470), .B2(new_n471), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n463), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n470), .B2(new_n471), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n466), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n511), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(new_n505), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n508), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n503), .A2(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n512), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n521), .B(new_n523), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n507), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  OR3_X1    g114(.A1(new_n538), .A2(new_n539), .A3(new_n507), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n538), .B2(new_n507), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n522), .A2(G81), .B1(new_n512), .B2(G43), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  AND2_X1   g125(.A1(KEYINPUT5), .A2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(KEYINPUT5), .A2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(KEYINPUT73), .A3(G651), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n558), .A2(new_n559), .B1(G91), .B2(new_n522), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n512), .A2(G53), .ZN(new_n561));
  NAND2_X1  g136(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n512), .A2(G53), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n565), .A2(KEYINPUT72), .A3(new_n566), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n560), .A2(new_n569), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n507), .B1(new_n553), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(G49), .B2(new_n512), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n522), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G288));
  AND2_X1   g153(.A1(G48), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n511), .ZN(new_n580));
  NOR2_X1   g155(.A1(KEYINPUT6), .A2(G651), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n514), .A2(KEYINPUT75), .A3(new_n579), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(new_n585), .B1(new_n522), .B2(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(G61), .B1(new_n551), .B2(new_n552), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT74), .B1(new_n589), .B2(G651), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n591));
  AOI211_X1 g166(.A(new_n591), .B(new_n507), .C1(new_n587), .C2(new_n588), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n586), .B1(new_n590), .B2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n507), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n512), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n515), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n522), .A2(G92), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT10), .Z(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n553), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n543), .A2(new_n612), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n608), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n466), .A2(new_n474), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n479), .A2(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n481), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n463), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT79), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G1341), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n642), .A2(G1341), .ZN(new_n645));
  OAI21_X1  g220(.A(G1348), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT78), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2451), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2454), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n649), .B(new_n651), .Z(new_n652));
  OR2_X1    g227(.A1(new_n642), .A2(G1341), .ZN(new_n653));
  INV_X1    g228(.A(G1348), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(new_n643), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n646), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n646), .A2(new_n655), .ZN(new_n658));
  INV_X1    g233(.A(new_n652), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  INV_X1    g244(.A(new_n662), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n669), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(KEYINPUT82), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(KEYINPUT82), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n683), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n687));
  MUX2_X1   g262(.A(new_n686), .B(new_n683), .S(new_n687), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(KEYINPUT83), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n685), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n693), .B1(new_n690), .B2(new_n692), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n675), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(new_n675), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n697), .A2(new_n700), .A3(new_n702), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G32), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G141), .ZN(new_n713));
  INV_X1    g288(.A(new_n481), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n474), .A2(G105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT90), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n479), .A2(G129), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n709), .B1(new_n721), .B2(new_n708), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT92), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT27), .B(G1996), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n708), .A2(G26), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT28), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n481), .A2(G140), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G104), .A2(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT88), .Z(new_n732));
  INV_X1    g307(.A(G116), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n473), .B1(new_n733), .B2(G2105), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n732), .A2(new_n734), .B1(new_n479), .B2(G128), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n727), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2067), .ZN(new_n738));
  INV_X1    g313(.A(G2090), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n708), .A2(G35), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G162), .B2(new_n708), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT29), .Z(new_n742));
  OAI211_X1 g317(.A(new_n725), .B(new_n738), .C1(new_n739), .C2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G20), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT94), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  INV_X1    g322(.A(G299), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n744), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT95), .B(G1956), .Z(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G19), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n544), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT86), .B(G1341), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n749), .A2(new_n750), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n751), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n744), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n744), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(G1966), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  OR2_X1    g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  NAND2_X1  g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n762), .A2(new_n708), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n633), .B2(new_n708), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n744), .A2(G5), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G171), .B2(new_n744), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n766), .B1(new_n768), .B2(G1961), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n760), .A2(new_n761), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G34), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G29), .B2(G160), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G2084), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  INV_X1    g353(.A(G139), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n714), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(new_n463), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G29), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G29), .B2(G33), .ZN(new_n786));
  INV_X1    g361(.A(G2072), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n776), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G2084), .B2(new_n775), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n768), .A2(G1961), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n708), .A2(G27), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G164), .B2(new_n708), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2078), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n790), .B(new_n793), .C1(new_n786), .C2(new_n787), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n744), .A2(G4), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n609), .B2(new_n744), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(new_n654), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n742), .A2(new_n739), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n789), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n743), .A2(new_n757), .A3(new_n771), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n708), .A2(G25), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n481), .A2(G131), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT84), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n804));
  INV_X1    g379(.A(G107), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(G2105), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n479), .B2(G119), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n801), .B1(new_n809), .B2(new_n708), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  XOR2_X1   g386(.A(new_n810), .B(new_n811), .Z(new_n812));
  INV_X1    g387(.A(KEYINPUT85), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n744), .A2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n599), .B2(new_n744), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1986), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n744), .A2(G22), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G166), .B2(new_n744), .ZN(new_n820));
  INV_X1    g395(.A(G1971), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(G6), .A2(G16), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G305), .B2(new_n744), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT32), .B(G1981), .Z(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n744), .A2(G23), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n576), .A2(new_n577), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n744), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT33), .B(G1976), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n822), .A2(new_n826), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n812), .A2(new_n813), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n818), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT36), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n800), .A2(new_n838), .ZN(G150));
  INV_X1    g414(.A(G150), .ZN(G311));
  AOI22_X1  g415(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n507), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n512), .A2(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n515), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n842), .A2(new_n845), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT96), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n543), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n544), .A2(new_n852), .A3(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n608), .A2(new_n616), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT97), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n847), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n850), .B1(new_n863), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n808), .B(new_n624), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n481), .A2(G142), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT100), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n870));
  INV_X1    g445(.A(G118), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(G2105), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n870), .B2(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n479), .A2(G130), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n866), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT102), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n499), .A2(new_n501), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n489), .A2(new_n494), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n487), .B1(new_n464), .B2(new_n465), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n463), .A2(G114), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT99), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n878), .A2(new_n880), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n736), .B(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(new_n784), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n784), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n721), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n892), .A2(new_n720), .A3(new_n888), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n877), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n633), .B(G160), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n485), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n720), .B1(new_n892), .B2(new_n888), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n889), .A2(new_n721), .A3(new_n890), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT102), .A4(new_n876), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n876), .B1(new_n891), .B2(new_n893), .ZN(new_n902));
  INV_X1    g477(.A(new_n876), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n898), .A3(new_n899), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n904), .A3(new_n896), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g483(.A1(G290), .A2(G288), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n829), .A2(new_n599), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT105), .ZN(new_n911));
  XNOR2_X1  g486(.A(G303), .B(G305), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT105), .B1(new_n909), .B2(new_n910), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n913), .A2(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT42), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(KEYINPUT106), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n858), .B(new_n619), .Z(new_n920));
  NOR2_X1   g495(.A1(G299), .A2(new_n608), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(G299), .A2(new_n608), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  INV_X1    g500(.A(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n919), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n922), .A2(KEYINPUT103), .A3(new_n923), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT103), .B1(new_n922), .B2(new_n923), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n920), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT104), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n918), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(KEYINPUT104), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n933), .B2(new_n920), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n919), .B(new_n929), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n918), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n851), .A2(new_n612), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(G331));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g522(.A1(G286), .A2(G301), .ZN(new_n948));
  NAND2_X1  g523(.A1(G168), .A2(G171), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n856), .A2(new_n948), .A3(new_n857), .A4(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n856), .A2(new_n857), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n927), .B(new_n924), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n916), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(new_n949), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n858), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n956), .A2(new_n923), .A3(new_n922), .A4(new_n950), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n906), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n954), .B1(new_n953), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n947), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n956), .B(new_n950), .C1(new_n931), .C2(new_n932), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n953), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n916), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n906), .A4(new_n958), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT44), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n959), .B2(new_n960), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n964), .A2(new_n947), .A3(new_n906), .A4(new_n958), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n961), .B2(new_n965), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT44), .B1(new_n968), .B2(new_n969), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT107), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n886), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G125), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n468), .B1(new_n478), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G2105), .ZN(new_n984));
  INV_X1    g559(.A(new_n476), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(G40), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT115), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n469), .A2(new_n989), .A3(new_n476), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n499), .A2(new_n501), .B1(new_n495), .B2(KEYINPUT99), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n880), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n988), .B(new_n990), .C1(new_n992), .C2(new_n979), .ZN(new_n993));
  INV_X1    g568(.A(new_n495), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n878), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n979), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n987), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1956), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT57), .B1(new_n565), .B2(new_n566), .ZN(new_n1000));
  AOI22_X1  g575(.A1(G299), .A2(KEYINPUT57), .B1(new_n560), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT112), .B(new_n1004), .C1(G164), .C2(G1384), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n886), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1003), .A2(new_n990), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT56), .B(G2072), .Z(new_n1008));
  OR2_X1    g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n999), .A2(new_n1001), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n998), .B2(new_n997), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1013), .B2(new_n1001), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1001), .ZN(new_n1015));
  INV_X1    g590(.A(new_n996), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n981), .A2(new_n986), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n988), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1956), .B1(new_n1018), .B2(new_n987), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT117), .B(new_n1015), .C1(new_n1019), .C2(new_n1012), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n886), .A2(new_n979), .A3(new_n980), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n990), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n886), .A2(new_n980), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(new_n986), .ZN(new_n1026));
  INV_X1    g601(.A(G2067), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1024), .A2(new_n654), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n608), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1010), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT61), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n999), .A2(new_n1001), .A3(new_n1009), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1001), .B1(new_n999), .B2(new_n1009), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n544), .A2(KEYINPUT119), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n986), .A2(G1996), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1003), .A2(new_n1005), .A3(new_n1036), .A4(new_n1006), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n990), .A2(new_n980), .A3(new_n886), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT58), .B(G1341), .Z(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT59), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n1035), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1028), .A2(KEYINPUT60), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1024), .A2(new_n654), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT60), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT121), .B1(new_n1052), .B2(new_n608), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n609), .C1(new_n1028), .C2(KEYINPUT60), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1049), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1053), .A2(new_n1049), .A3(new_n1055), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1034), .B(new_n1048), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1010), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n999), .A2(KEYINPUT120), .A3(new_n1001), .A4(new_n1009), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT61), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1021), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1030), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1007), .B2(G2078), .ZN(new_n1066));
  INV_X1    g641(.A(G1961), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1024), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1025), .A2(new_n1004), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1065), .A2(G2078), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n995), .A2(KEYINPUT45), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n990), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1068), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1075));
  OAI211_X1 g650(.A(G301), .B(new_n1066), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT54), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1025), .A2(KEYINPUT108), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n1025), .B2(KEYINPUT108), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G2078), .ZN(new_n1082));
  AND4_X1   g657(.A1(KEYINPUT53), .A2(new_n1006), .A3(new_n1082), .A4(new_n990), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1081), .A2(new_n1083), .B1(new_n1067), .B2(new_n1024), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1066), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1085), .B2(G171), .ZN(new_n1086));
  AOI211_X1 g661(.A(KEYINPUT123), .B(G301), .C1(new_n1084), .C2(new_n1066), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1077), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1966), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1071), .A2(new_n990), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT45), .B1(new_n886), .B2(new_n980), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2084), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1022), .A2(new_n1023), .A3(new_n1093), .A4(new_n990), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(G168), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT51), .B1(new_n1095), .B2(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G168), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1092), .A2(G286), .A3(new_n1094), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1007), .A2(new_n821), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n997), .B2(G2090), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G8), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G303), .A2(G8), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1024), .A2(G2090), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1103), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n1108), .A3(G8), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n1114));
  INV_X1    g689(.A(G1981), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n586), .B(new_n1115), .C1(new_n590), .C2(new_n592), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n588), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n505), .B2(G61), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n591), .B1(new_n1119), .B2(new_n507), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n589), .A2(KEYINPUT74), .A3(G651), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1115), .B1(new_n1122), .B2(new_n586), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1114), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G305), .A2(G1981), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT49), .A3(new_n1116), .ZN(new_n1126));
  INV_X1    g701(.A(G8), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n992), .B2(new_n990), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT114), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1124), .A2(new_n1131), .A3(new_n1128), .A4(new_n1126), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n576), .A2(G1976), .A3(new_n577), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1039), .A2(G8), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OR3_X1    g711(.A1(new_n829), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1130), .A2(new_n1132), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1102), .A2(new_n1110), .A3(new_n1113), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(G171), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1084), .A2(G301), .A3(new_n1066), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT54), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1088), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1064), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1102), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1143), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1113), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1108), .B1(new_n1104), .B2(G8), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1102), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1151), .A2(new_n1152), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1097), .A2(G8), .A3(G168), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1110), .A2(new_n1140), .A3(new_n1113), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1155), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1108), .B1(new_n1112), .B2(G8), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1165), .A2(new_n1163), .A3(new_n1160), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1162), .A2(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(G288), .A2(G1976), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1153), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1116), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1128), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1113), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1140), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT116), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1155), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1177), .B2(KEYINPUT63), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1170), .A2(new_n1128), .B1(new_n1172), .B2(new_n1140), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1147), .A2(new_n1159), .A3(new_n1175), .A4(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1079), .A2(new_n990), .A3(new_n1080), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(G1996), .A3(new_n720), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT110), .Z(new_n1186));
  OR2_X1    g761(.A1(new_n1183), .A2(G1996), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1187), .A2(new_n720), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n736), .A2(G2067), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n730), .A2(new_n1027), .A3(new_n735), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1184), .A2(new_n1191), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1192), .A2(KEYINPUT111), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(KEYINPUT111), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1188), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n809), .A2(new_n811), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n809), .A2(new_n811), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1184), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1186), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(G1986), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n599), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT109), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1204), .B1(new_n1201), .B2(new_n599), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1200), .B1(new_n1184), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1182), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1186), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1190), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1208), .B1(new_n1210), .B2(new_n1184), .ZN(new_n1211));
  AOI211_X1 g786(.A(KEYINPUT125), .B(new_n1183), .C1(new_n1209), .C2(new_n1190), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1184), .B1(new_n720), .B2(new_n1191), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT126), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT47), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1187), .B(KEYINPUT46), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1215), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1204), .A2(new_n1183), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT48), .ZN(new_n1221));
  OAI22_X1  g796(.A1(new_n1218), .A2(new_n1219), .B1(new_n1200), .B2(new_n1221), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1211), .A2(new_n1212), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1207), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g799(.A(new_n907), .B1(new_n968), .B2(new_n969), .ZN(new_n1226));
  OR2_X1    g800(.A1(G227), .A2(new_n461), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n657), .B2(new_n660), .ZN(new_n1228));
  AND3_X1   g802(.A1(new_n706), .A2(new_n1228), .A3(KEYINPUT127), .ZN(new_n1229));
  AOI21_X1  g803(.A(KEYINPUT127), .B1(new_n706), .B2(new_n1228), .ZN(new_n1230));
  OAI21_X1  g804(.A(new_n1226), .B1(new_n1229), .B2(new_n1230), .ZN(G225));
  INV_X1    g805(.A(G225), .ZN(G308));
endmodule


