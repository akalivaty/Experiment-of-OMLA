//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n643, new_n645, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G567), .B1(new_n456), .B2(G2106), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n461), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT70), .B1(new_n461), .B2(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT71), .A3(G101), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G137), .A4(new_n461), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n462), .A2(new_n463), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n465), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n480), .B1(new_n468), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n468), .A2(KEYINPUT72), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n471), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n461), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G136), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(new_n488), .B2(new_n490), .ZN(new_n494));
  OAI221_X1 g069(.A(new_n487), .B1(new_n491), .B2(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n461), .A2(G138), .ZN(new_n498));
  OAI211_X1 g073(.A(KEYINPUT73), .B(new_n497), .C1(new_n468), .C2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n471), .A2(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n498), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n497), .A2(KEYINPUT73), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n497), .A2(KEYINPUT73), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n471), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n499), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n517), .A2(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n515), .A2(new_n525), .ZN(G166));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT74), .B1(new_n512), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(KEYINPUT74), .B(new_n534), .C1(new_n520), .C2(new_n519), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n528), .B(new_n533), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n512), .A2(new_n516), .A3(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n542), .B1(new_n539), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n534), .B1(new_n520), .B2(new_n519), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(new_n536), .B1(G51), .B2(new_n532), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n528), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n527), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n539), .A2(new_n541), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n555), .A2(new_n557), .A3(KEYINPUT77), .A4(new_n538), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n551), .A2(new_n558), .ZN(G168));
  NAND2_X1  g134(.A1(G77), .A2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n520), .A2(new_n519), .ZN(new_n561));
  INV_X1    g136(.A(G64), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n514), .B1(new_n563), .B2(KEYINPUT78), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n564), .B1(KEYINPUT78), .B2(new_n563), .ZN(new_n565));
  INV_X1    g140(.A(new_n523), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G90), .B1(G52), .B2(new_n532), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G301));
  INV_X1    g143(.A(G301), .ZN(G171));
  AOI22_X1  g144(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n514), .ZN(new_n571));
  INV_X1    g146(.A(G43), .ZN(new_n572));
  INV_X1    g147(.A(G81), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n517), .A2(new_n572), .B1(new_n523), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  AND2_X1   g155(.A1(KEYINPUT79), .A2(G53), .ZN(new_n581));
  OAI211_X1 g156(.A(G543), .B(new_n581), .C1(new_n521), .C2(new_n522), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT9), .Z(new_n583));
  AOI22_X1  g158(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G91), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n584), .A2(new_n514), .B1(new_n585), .B2(new_n523), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT80), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G78), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G65), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n561), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(G651), .A2(new_n590), .B1(new_n566), .B2(G91), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n582), .B(KEYINPUT9), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G299));
  INV_X1    g171(.A(G168), .ZN(G286));
  OR2_X1    g172(.A1(new_n515), .A2(new_n525), .ZN(G303));
  INV_X1    g173(.A(G74), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n514), .B1(new_n561), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(G49), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n516), .A2(KEYINPUT82), .A3(G49), .A4(G543), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n606));
  INV_X1    g181(.A(G87), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n523), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT81), .A4(G87), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(G288));
  NAND2_X1  g186(.A1(new_n512), .A2(G61), .ZN(new_n612));
  NAND2_X1  g187(.A1(G73), .A2(G543), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n514), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n566), .A2(G86), .B1(G48), .B2(new_n532), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(G305));
  AOI22_X1  g192(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(new_n514), .ZN(new_n619));
  INV_X1    g194(.A(G47), .ZN(new_n620));
  INV_X1    g195(.A(G85), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n517), .A2(new_n620), .B1(new_n523), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(G290));
  NAND2_X1  g199(.A1(G301), .A2(G868), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT83), .B1(new_n523), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n512), .A2(new_n516), .A3(new_n628), .A4(G92), .ZN(new_n629));
  AOI21_X1  g204(.A(KEYINPUT10), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n532), .A2(G54), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(new_n514), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n629), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n625), .B1(new_n637), .B2(G868), .ZN(G321));
  XOR2_X1   g213(.A(G321), .B(KEYINPUT84), .Z(G284));
  NOR2_X1   g214(.A1(G299), .A2(G868), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g216(.A(new_n640), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g217(.A(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n637), .B1(new_n643), .B2(G860), .ZN(G148));
  OAI21_X1  g219(.A(KEYINPUT85), .B1(new_n575), .B2(G868), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n637), .A2(new_n643), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G868), .ZN(new_n647));
  MUX2_X1   g222(.A(KEYINPUT85), .B(new_n645), .S(new_n647), .Z(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n464), .A2(new_n471), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  INV_X1    g228(.A(new_n491), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G135), .ZN(new_n655));
  INV_X1    g230(.A(new_n494), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G123), .ZN(new_n657));
  OR2_X1    g232(.A1(G99), .A2(G2105), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n658), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2096), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n653), .A2(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT87), .Z(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n665), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2427), .B(G2438), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2430), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT15), .B(G2435), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  AND3_X1   g251(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT14), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G14), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n671), .A2(new_n677), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(G401));
  XOR2_X1   g256(.A(G2067), .B(G2678), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT90), .Z(new_n684));
  NOR2_X1   g259(.A1(G2072), .A2(G2078), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n442), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2084), .B(G2090), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n686), .B(KEYINPUT91), .Z(new_n691));
  OAI211_X1 g266(.A(new_n689), .B(new_n690), .C1(new_n684), .C2(new_n691), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n683), .A2(new_n686), .A3(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT18), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n684), .A2(new_n690), .A3(new_n688), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G2096), .B(G2100), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G227));
  XOR2_X1   g273(.A(G1971), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  XOR2_X1   g275(.A(G1956), .B(G2474), .Z(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT20), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n700), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n700), .B2(new_n706), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(G1991), .B(G1996), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(G229));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G35), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT103), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n495), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G2090), .ZN(new_n724));
  INV_X1    g299(.A(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n718), .A2(G32), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT26), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n464), .A2(G105), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G141), .ZN(new_n732));
  INV_X1    g307(.A(G129), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n731), .B1(new_n491), .B2(new_n732), .C1(new_n733), .C2(new_n494), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n726), .B1(new_n735), .B2(new_n718), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(KEYINPUT27), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(KEYINPUT27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n725), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n736), .A2(KEYINPUT27), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(KEYINPUT27), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n740), .A2(G1996), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n721), .B(KEYINPUT29), .ZN(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND4_X1   g320(.A1(new_n724), .A2(new_n739), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT98), .B(KEYINPUT28), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n718), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n461), .A2(G116), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n656), .A2(G128), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n654), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(G29), .ZN(new_n757));
  AOI211_X1 g332(.A(KEYINPUT97), .B(new_n718), .C1(new_n754), .C2(new_n755), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n749), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G4), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n637), .B2(new_n762), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT96), .B(G1348), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n764), .B(new_n765), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n595), .B2(new_n762), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT104), .B(G1956), .Z(new_n770));
  XOR2_X1   g345(.A(new_n769), .B(new_n770), .Z(new_n771));
  NOR2_X1   g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n484), .A2(G29), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n762), .A2(G5), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G301), .B2(G16), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n778), .A2(G2084), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n773), .A2(new_n783), .A3(new_n777), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n782), .B(new_n784), .C1(new_n779), .C2(new_n781), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  AOI22_X1  g362(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  INV_X1    g363(.A(G139), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(new_n461), .B2(new_n788), .C1(new_n491), .C2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G2072), .ZN(new_n792));
  INV_X1    g367(.A(G28), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT30), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n793), .B2(KEYINPUT30), .ZN(new_n795));
  OR2_X1    g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  NAND2_X1  g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G2078), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n718), .A2(G27), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT102), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n510), .B2(G29), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n792), .B(new_n798), .C1(new_n799), .C2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n660), .A2(new_n804), .A3(new_n718), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n660), .B2(new_n718), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n805), .B(new_n806), .C1(G2072), .C2(new_n791), .ZN(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G19), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n575), .B2(G16), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n809), .A2(G1341), .B1(new_n799), .B2(new_n802), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G1341), .B2(new_n809), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n785), .A2(new_n803), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n746), .A2(new_n761), .A3(new_n772), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n762), .A2(G21), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G168), .B2(new_n762), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(G1966), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT101), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(G1966), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT99), .Z(new_n819));
  NOR3_X1   g394(.A1(new_n813), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT105), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  OR2_X1    g397(.A1(G6), .A2(G16), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G305), .B2(new_n762), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT32), .B(G1981), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G23), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT94), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G288), .B2(new_n762), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT33), .B(G1976), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n762), .A2(G22), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G166), .B2(new_n762), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT95), .B(G1971), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n829), .A2(new_n831), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n822), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n826), .A2(new_n832), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n841), .A2(KEYINPUT34), .A3(new_n838), .A4(new_n837), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n762), .A2(G24), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n623), .B2(new_n762), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(G1986), .Z(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n654), .A2(G131), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n656), .A2(G119), .ZN(new_n849));
  OR2_X1    g424(.A1(G95), .A2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G29), .ZN(new_n854));
  OR2_X1    g429(.A1(G25), .A2(G29), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT35), .B(G1991), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT93), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n860), .A3(new_n855), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n847), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n843), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT36), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n820), .A2(new_n821), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n821), .B1(new_n820), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(G311));
  NAND2_X1  g442(.A1(new_n820), .A2(new_n864), .ZN(G150));
  NAND2_X1  g443(.A1(new_n637), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n514), .ZN(new_n872));
  INV_X1    g447(.A(G55), .ZN(new_n873));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n517), .A2(new_n873), .B1(new_n523), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n575), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n870), .B(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  INV_X1    g455(.A(G860), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n876), .A2(new_n881), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G145));
  XNOR2_X1  g461(.A(G160), .B(new_n660), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G162), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n890));
  INV_X1    g465(.A(G142), .ZN(new_n891));
  INV_X1    g466(.A(G130), .ZN(new_n892));
  OAI221_X1 g467(.A(new_n890), .B1(new_n491), .B2(new_n891), .C1(new_n892), .C2(new_n494), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(new_n651), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n651), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n853), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n756), .A2(new_n510), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n754), .A2(G164), .A3(new_n755), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n735), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n790), .A2(KEYINPUT106), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n734), .A3(new_n901), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(KEYINPUT106), .A3(new_n790), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n896), .A2(new_n897), .A3(new_n852), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n790), .A2(KEYINPUT106), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n903), .A2(new_n909), .A3(new_n904), .A4(new_n905), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n899), .A2(new_n907), .A3(new_n908), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n899), .A2(new_n908), .B1(new_n907), .B2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n888), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n899), .A2(new_n908), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n907), .A2(new_n910), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n888), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n911), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g497(.A(new_n646), .B(new_n877), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n595), .A2(new_n636), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n587), .A2(new_n634), .A3(new_n594), .A4(new_n635), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(KEYINPUT41), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  INV_X1    g502(.A(new_n925), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n587), .A2(new_n594), .B1(new_n634), .B2(new_n635), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n925), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  OR3_X1    g508(.A1(new_n931), .A2(new_n933), .A3(KEYINPUT110), .ZN(new_n934));
  AND2_X1   g509(.A1(G166), .A2(KEYINPUT109), .ZN(new_n935));
  NOR2_X1   g510(.A1(G166), .A2(KEYINPUT109), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(G290), .A2(KEYINPUT108), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n623), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n938), .B(new_n940), .C1(new_n935), .C2(new_n936), .ZN(new_n943));
  XNOR2_X1  g518(.A(G288), .B(G305), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n942), .B2(new_n943), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT42), .Z(new_n948));
  AND2_X1   g523(.A1(new_n934), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT110), .B1(new_n931), .B2(new_n933), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n934), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(G868), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(G868), .B2(new_n876), .ZN(G295));
  OAI21_X1  g528(.A(new_n952), .B1(G868), .B2(new_n876), .ZN(G331));
  NAND2_X1  g529(.A1(new_n930), .A2(new_n926), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n551), .A2(new_n558), .A3(G301), .ZN(new_n956));
  AOI21_X1  g531(.A(G301), .B1(new_n551), .B2(new_n558), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n956), .A2(new_n957), .A3(new_n877), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n553), .A2(new_n554), .B1(new_n549), .B2(new_n528), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT77), .B1(new_n959), .B2(new_n557), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n545), .A2(new_n527), .A3(new_n550), .ZN(new_n961));
  OAI21_X1  g536(.A(G171), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n551), .A2(new_n558), .A3(G301), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n878), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n958), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n877), .B1(new_n956), .B2(new_n957), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n878), .A3(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n932), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n947), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n965), .A2(new_n947), .A3(KEYINPUT112), .A4(new_n968), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT43), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n947), .B1(new_n965), .B2(new_n968), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(G37), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n972), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n974), .B2(G37), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n966), .A2(new_n967), .A3(new_n932), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n966), .A2(new_n967), .B1(new_n930), .B2(new_n926), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(KEYINPUT111), .B(new_n915), .C1(new_n981), .C2(new_n947), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n976), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  AOI221_X4 g558(.A(KEYINPUT44), .B1(new_n973), .B2(new_n975), .C1(new_n983), .C2(KEYINPUT43), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n976), .A2(new_n975), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n973), .A2(new_n978), .A3(new_n982), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n984), .A2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n510), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n482), .B2(G2105), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n996), .A2(new_n465), .A3(new_n474), .A4(new_n478), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n852), .B(new_n860), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT115), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n756), .B(new_n760), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n734), .B(new_n725), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n998), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G290), .A2(G1986), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n1007));
  OR3_X1    g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(G290), .A2(new_n1007), .A3(G1986), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n998), .A3(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT114), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n615), .B2(new_n616), .ZN(new_n1015));
  INV_X1    g590(.A(G48), .ZN(new_n1016));
  INV_X1    g591(.A(G86), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n517), .A2(new_n1016), .B1(new_n523), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1018), .A2(new_n614), .A3(G1981), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1013), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n615), .A2(new_n616), .A3(new_n1014), .ZN(new_n1021));
  OAI21_X1  g596(.A(G1981), .B1(new_n1018), .B2(new_n614), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(G8), .B1(new_n997), .B2(new_n992), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n605), .A2(new_n610), .A3(G1976), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(G8), .C1(new_n997), .C2(new_n992), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n605), .A2(new_n610), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(G1976), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1024), .A2(new_n1025), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1027), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n1028), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1027), .A2(KEYINPUT120), .A3(KEYINPUT52), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G303), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT118), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n1040));
  NAND4_X1  g615(.A1(G303), .A2(new_n1040), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT119), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1044), .A3(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n474), .A2(new_n996), .A3(new_n465), .A4(new_n478), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n993), .A2(G1384), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n510), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n994), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT116), .ZN(new_n1053));
  INV_X1    g628(.A(G1971), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n992), .A2(new_n993), .B1(new_n510), .B2(new_n1050), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n1049), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n510), .A2(new_n1060), .A3(new_n991), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1049), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(G2090), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1048), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1036), .B1(new_n1047), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1058), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1053), .A2(KEYINPUT117), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1048), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1066), .B1(new_n1047), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1055), .A2(new_n1049), .A3(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n583), .A2(KEYINPUT57), .A3(new_n586), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n591), .B2(new_n593), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n510), .A2(new_n1060), .A3(new_n991), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1060), .B1(new_n510), .B2(new_n991), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n997), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT122), .B(G1956), .Z(new_n1083));
  OAI211_X1 g658(.A(new_n1075), .B(new_n1079), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1083), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1062), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1079), .B1(new_n1086), .B2(new_n1075), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1062), .A2(new_n1088), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n997), .A2(new_n992), .A3(G2067), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n636), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1073), .B(new_n1084), .C1(new_n1087), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1081), .A2(new_n997), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1083), .B1(new_n1095), .B2(new_n1061), .ZN(new_n1096));
  AND4_X1   g671(.A1(new_n1049), .A2(new_n994), .A3(new_n1051), .A4(new_n1074), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1096), .A2(new_n1097), .B1(new_n1078), .B2(new_n1076), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1348), .B1(new_n1095), .B2(new_n1061), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n637), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1073), .B1(new_n1101), .B2(new_n1084), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1084), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1087), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT124), .B(new_n1104), .C1(new_n1105), .C2(new_n1087), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n1091), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n636), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n637), .A4(new_n1091), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1098), .A2(KEYINPUT61), .A3(new_n1084), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  INV_X1    g693(.A(new_n992), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1049), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(G1996), .B2(new_n1052), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1118), .B1(new_n1123), .B2(new_n575), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1123), .A2(new_n1118), .A3(new_n575), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1116), .B(new_n1117), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1103), .B1(new_n1110), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1057), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1056), .B1(new_n1055), .B2(new_n1049), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n799), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1131), .A2(G2078), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1082), .A2(G1961), .B1(new_n1052), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(G301), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(G171), .B(new_n1135), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT54), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(G2078), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1140), .B2(KEYINPUT53), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1132), .A2(G301), .A3(new_n1136), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1082), .A2(new_n783), .ZN(new_n1147));
  INV_X1    g722(.A(G1966), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1052), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1048), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n1152));
  OAI22_X1  g727(.A1(G168), .A2(new_n1048), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR4_X1   g728(.A1(new_n1150), .A2(new_n1153), .A3(KEYINPUT126), .A4(KEYINPUT51), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(G8), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1153), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1156), .A2(new_n1157), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1150), .A2(KEYINPUT125), .A3(G286), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT125), .B1(new_n1150), .B2(G286), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n1154), .A2(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1127), .A2(new_n1146), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(KEYINPUT62), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  OAI221_X1 g739(.A(new_n1164), .B1(new_n1159), .B2(new_n1160), .C1(new_n1154), .C2(new_n1158), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1165), .A3(new_n1137), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1072), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1156), .A2(G286), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n1071), .B2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1070), .A2(new_n1047), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1070), .A2(new_n1047), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(KEYINPUT63), .A3(new_n1036), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1070), .A2(new_n1047), .A3(new_n1036), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1175), .A2(G1976), .A3(G288), .ZN(new_n1176));
  OAI211_X1 g751(.A(G8), .B(new_n1120), .C1(new_n1176), .C2(new_n1019), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1174), .A2(KEYINPUT121), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT121), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1169), .A2(new_n1173), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1012), .B1(new_n1167), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n998), .A2(new_n725), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT46), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1001), .A2(new_n735), .ZN(new_n1184));
  INV_X1    g759(.A(new_n998), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT47), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n1187), .A2(KEYINPUT127), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(KEYINPUT127), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1001), .A2(new_n860), .A3(new_n853), .A4(new_n1002), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n754), .A2(new_n760), .A3(new_n755), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1185), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n998), .A2(new_n1006), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT48), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1192), .B1(new_n1004), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1188), .A2(new_n1189), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1181), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g772(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n975), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g775(.A(G319), .B1(new_n679), .B2(new_n680), .ZN(new_n1202));
  NOR2_X1   g776(.A1(G227), .A2(new_n1202), .ZN(new_n1203));
  AND2_X1   g777(.A1(new_n716), .A2(new_n1203), .ZN(new_n1204));
  AND3_X1   g778(.A1(new_n1201), .A2(new_n921), .A3(new_n1204), .ZN(G308));
  NAND3_X1  g779(.A1(new_n1201), .A2(new_n921), .A3(new_n1204), .ZN(G225));
endmodule


