//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT64), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n461), .A2(new_n462), .B1(G113), .B2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n463), .B1(new_n462), .B2(new_n461), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT65), .B(G2105), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g042(.A(KEYINPUT67), .B(G2104), .Z(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT69), .Z(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(new_n477), .A3(KEYINPUT3), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G137), .A3(new_n465), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n479), .A2(new_n466), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n479), .A2(new_n490), .A3(new_n466), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n492), .B2(G124), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT71), .Z(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND3_X1  g070(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(new_n484), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n479), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n465), .A2(new_n460), .A3(G138), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT72), .A2(G114), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT72), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(G2105), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n500), .A2(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT74), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n516), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G543), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n523), .A2(new_n514), .A3(new_n524), .ZN(new_n527));
  AOI22_X1  g102(.A1(G50), .A2(new_n526), .B1(new_n527), .B2(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n518), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n526), .A2(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n527), .A2(G89), .ZN(new_n532));
  AND2_X1   g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n516), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n536), .A2(G63), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n531), .A2(new_n532), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(new_n526), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n516), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n527), .A2(G90), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n516), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n523), .A2(G43), .A3(G543), .A4(new_n524), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n523), .A2(G81), .A3(new_n514), .A4(new_n524), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n553), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n533), .B2(new_n534), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n512), .A2(new_n567), .A3(new_n513), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(G78), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n527), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n564), .A2(new_n571), .A3(new_n572), .ZN(G299));
  OAI21_X1  g148(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT78), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(G49), .B2(new_n526), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n527), .A2(G87), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n535), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT79), .ZN(new_n585));
  AOI22_X1  g160(.A1(G48), .A2(new_n526), .B1(new_n527), .B2(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n535), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT80), .B(new_n588), .C1(new_n535), .C2(new_n589), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n592), .A2(G651), .A3(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(KEYINPUT81), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(KEYINPUT81), .ZN(new_n596));
  AOI22_X1  g171(.A1(G47), .A2(new_n526), .B1(new_n527), .B2(G85), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n523), .A2(G92), .A3(new_n514), .A4(new_n524), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT10), .ZN(new_n601));
  NOR3_X1   g176(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT76), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n567), .B1(new_n512), .B2(new_n513), .ZN(new_n603));
  OAI21_X1  g178(.A(G66), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n516), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n523), .A2(G54), .A3(G543), .A4(new_n524), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT82), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n566), .B2(new_n568), .ZN(new_n611));
  INV_X1    g186(.A(new_n605), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n613), .A2(new_n614), .A3(new_n607), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n601), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n599), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n599), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(new_n601), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n613), .A2(new_n614), .A3(new_n607), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n614), .B1(new_n613), .B2(new_n607), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G860), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n626), .B1(G559), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT83), .Z(G148));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n556), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n626), .A2(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(new_n630), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n466), .B2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n485), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G135), .ZN(new_n639));
  INV_X1    g214(.A(new_n492), .ZN(new_n640));
  INV_X1    g215(.A(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n469), .A2(new_n460), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT13), .B(G2100), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n644), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(G14), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT86), .ZN(G401));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2096), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n683), .A2(new_n685), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n681), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n689), .A2(new_n686), .A3(new_n681), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n687), .B1(new_n686), .B2(new_n681), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(G6), .ZN(new_n707));
  INV_X1    g282(.A(G305), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n702), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n702), .A2(G23), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G288), .B2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT33), .B(G1976), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT91), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT92), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n706), .B(new_n711), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  OAI221_X1 g298(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n465), .C2(G107), .ZN(new_n724));
  INV_X1    g299(.A(G131), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n485), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n492), .B2(G119), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n723), .B1(new_n727), .B2(new_n722), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT90), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT35), .B(G1991), .Z(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n731), .ZN(new_n733));
  MUX2_X1   g308(.A(G24), .B(G290), .S(G16), .Z(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1986), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n721), .A2(new_n732), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT29), .B(G2090), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n492), .A2(G129), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT26), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n469), .A2(G105), .ZN(new_n746));
  INV_X1    g321(.A(G141), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n745), .B(new_n746), .C1(new_n485), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(new_n722), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n722), .B2(G32), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT93), .B(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n616), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G4), .B2(G16), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n751), .A2(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n753), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n756), .B(new_n757), .C1(new_n751), .C2(new_n752), .ZN(new_n758));
  NOR2_X1   g333(.A1(G171), .A2(new_n702), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G5), .B2(new_n702), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT99), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n557), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G16), .B2(G19), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(G1341), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n702), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1956), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G1341), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n765), .ZN(new_n774));
  INV_X1    g349(.A(new_n642), .ZN(new_n775));
  INV_X1    g350(.A(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(G29), .A2(G33), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n638), .A2(G139), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT96), .B(KEYINPUT25), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n460), .A2(G127), .ZN(new_n783));
  INV_X1    g358(.A(G115), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n472), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n782), .B1(new_n466), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n778), .B1(new_n787), .B2(new_n722), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n775), .A2(G29), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G34), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(KEYINPUT24), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(KEYINPUT24), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(KEYINPUT97), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(KEYINPUT97), .B2(new_n792), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n481), .B2(new_n722), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2084), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n789), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(G164), .A2(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G27), .B2(G29), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  INV_X1    g375(.A(G1966), .ZN(new_n801));
  NAND2_X1  g376(.A1(G168), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G16), .B2(G21), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n801), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n804), .B(new_n805), .C1(new_n800), .C2(new_n799), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT98), .B(G28), .Z(new_n807));
  AOI21_X1  g382(.A(G29), .B1(new_n807), .B2(KEYINPUT30), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(KEYINPUT30), .B2(new_n807), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n760), .B2(new_n761), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n776), .B2(new_n788), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n797), .A2(new_n806), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n767), .A2(new_n774), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n722), .A2(G26), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT28), .Z(new_n817));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(G116), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n466), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n638), .B2(G140), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G128), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n489), .B2(new_n491), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n818), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(KEYINPUT94), .B(new_n822), .C1(new_n640), .C2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n817), .B1(new_n828), .B2(G29), .ZN(new_n829));
  INV_X1    g404(.A(G2067), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR4_X1   g406(.A1(new_n742), .A2(new_n758), .A3(new_n815), .A4(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n738), .A2(new_n833), .ZN(G311));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n737), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n832), .ZN(G150));
  NAND2_X1  g412(.A1(new_n526), .A2(G55), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n516), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n527), .A2(G93), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  AND3_X1   g419(.A1(new_n556), .A2(KEYINPUT101), .A3(new_n842), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n556), .A2(KEYINPUT101), .ZN(new_n847));
  INV_X1    g422(.A(new_n842), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(new_n550), .C1(new_n554), .C2(new_n555), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n616), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n855));
  XOR2_X1   g430(.A(new_n854), .B(new_n855), .Z(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n627), .B1(new_n857), .B2(KEYINPUT39), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n844), .B1(new_n858), .B2(new_n859), .ZN(G145));
  INV_X1    g435(.A(new_n749), .ZN(new_n861));
  AOI21_X1  g436(.A(G164), .B1(new_n826), .B2(new_n827), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n826), .A2(new_n827), .A3(G164), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n787), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  INV_X1    g441(.A(new_n787), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n866), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n861), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n492), .A2(G130), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n638), .A2(G142), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n465), .A2(new_n872), .A3(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n465), .B2(G118), .ZN(new_n874));
  OR2_X1    g449(.A1(G106), .A2(G2105), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(G2104), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n870), .B(new_n871), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(new_n727), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n727), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n647), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n647), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n863), .A2(new_n787), .A3(new_n864), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n867), .B1(new_n866), .B2(new_n862), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n749), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n869), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n869), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(KEYINPUT103), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n869), .A2(new_n891), .A3(new_n884), .A4(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G162), .A2(new_n775), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n494), .A2(new_n642), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n894), .A2(G160), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(G160), .B1(new_n894), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n888), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n889), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT40), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n898), .B1(new_n890), .B2(new_n892), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n906), .A2(new_n907), .A3(new_n903), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n905), .A2(new_n908), .ZN(G395));
  NAND2_X1  g484(.A1(new_n842), .A2(new_n630), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT104), .B1(new_n616), .B2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n616), .A2(G299), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n626), .A2(new_n913), .A3(new_n620), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT41), .A4(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n852), .B(new_n632), .ZN(new_n920));
  MUX2_X1   g495(.A(new_n915), .B(new_n919), .S(new_n920), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n596), .A2(new_n597), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(new_n579), .A3(new_n576), .A4(new_n595), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n923), .A2(new_n595), .B1(new_n576), .B2(new_n579), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT105), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G303), .B(G305), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n931), .A2(new_n928), .A3(new_n929), .A4(new_n924), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n922), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n910), .B1(new_n936), .B2(new_n630), .ZN(G295));
  OAI21_X1  g512(.A(new_n910), .B1(new_n936), .B2(new_n630), .ZN(G331));
  NAND2_X1  g513(.A1(G171), .A2(G168), .ZN(new_n939));
  NAND2_X1  g514(.A1(G301), .A2(G286), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n850), .A2(new_n848), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n551), .A2(new_n552), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT75), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n849), .B1(new_n946), .B2(new_n550), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n948), .B2(new_n845), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n846), .A2(new_n851), .A3(new_n940), .A4(new_n939), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n919), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n915), .A2(new_n949), .A3(new_n950), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n917), .A2(new_n918), .B1(new_n950), .B2(new_n949), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT106), .B1(new_n957), .B2(new_n954), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n933), .A2(new_n934), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n901), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n954), .B1(new_n919), .B2(new_n951), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n935), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n961), .B1(new_n960), .B2(new_n901), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(KEYINPUT43), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n917), .A2(new_n970), .A3(new_n918), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n951), .B1(new_n917), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n955), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n959), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n963), .B2(new_n935), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n967), .A2(new_n968), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n965), .B2(new_n966), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(new_n975), .A3(new_n969), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT109), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n974), .A2(new_n975), .A3(new_n982), .A4(new_n969), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n978), .B1(new_n985), .B2(new_n968), .ZN(new_n986));
  AOI211_X1 g561(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n979), .C2(new_n984), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n977), .B1(new_n986), .B2(new_n987), .ZN(G397));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n471), .A2(new_n989), .A3(G40), .A4(new_n480), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n480), .A2(G40), .A3(new_n467), .A4(new_n470), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT111), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n499), .B2(new_n507), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(KEYINPUT112), .A3(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(KEYINPUT114), .A3(new_n999), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n828), .A2(G2067), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n826), .A2(new_n827), .A3(new_n830), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n749), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n998), .A2(new_n1008), .A3(new_n999), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1004), .A2(new_n1007), .B1(KEYINPUT46), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT127), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1011), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1010), .A2(new_n749), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1005), .B(new_n1006), .C1(new_n1008), .C2(new_n749), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1002), .A2(new_n1020), .A3(new_n1003), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1004), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n727), .B(new_n731), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1019), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1000), .A2(G1986), .A3(G290), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT48), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1017), .A2(new_n1018), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1021), .A2(new_n1019), .A3(new_n730), .A4(new_n727), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT126), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n1006), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1028), .B2(new_n1006), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1022), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n508), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT50), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n994), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1037), .A2(new_n990), .A3(new_n992), .A4(new_n1039), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1040), .A2(G2090), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(new_n990), .A3(new_n992), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n705), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1034), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT55), .Z(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(new_n1054));
  INV_X1    g629(.A(G288), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G1976), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(KEYINPUT116), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(KEYINPUT116), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n1059), .A3(KEYINPUT52), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  OR2_X1    g636(.A1(G305), .A2(G1981), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n586), .A2(new_n584), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G1981), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1065), .B2(KEYINPUT117), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(KEYINPUT49), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1054), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1057), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1069), .A2(new_n1071), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1053), .A2(new_n1060), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1044), .A2(new_n990), .A3(new_n992), .A4(new_n1045), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n801), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(G2084), .B2(new_n1040), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(G8), .A3(G168), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1076), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1050), .A2(KEYINPUT119), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1050), .A2(KEYINPUT119), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n1052), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(new_n1053), .A3(new_n1060), .A4(new_n1075), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1082), .A2(KEYINPUT63), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G168), .A2(new_n1034), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1966), .B1(new_n1092), .B2(new_n993), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1040), .A2(G2084), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(KEYINPUT51), .B(new_n1091), .C1(new_n1095), .C2(new_n1034), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(G8), .C1(new_n1080), .C2(G286), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1080), .A2(new_n1099), .A3(new_n1090), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1099), .B1(new_n1080), .B2(new_n1090), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1096), .B(new_n1098), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1040), .A2(new_n761), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(G2078), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1092), .A2(new_n993), .A3(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1046), .A2(new_n1048), .A3(G2078), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1105), .B(new_n1108), .C1(new_n1109), .C2(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1076), .A2(new_n1111), .A3(new_n1077), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1102), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1100), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1104), .A2(new_n1112), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1073), .A3(new_n1055), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1062), .B(KEYINPUT118), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1070), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1053), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1060), .A2(new_n1075), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1089), .A2(new_n1117), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(G299), .B(KEYINPUT57), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1040), .A2(new_n771), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1054), .A2(G2067), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n753), .B2(new_n1040), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(new_n626), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1129), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1135), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1131), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1131), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1126), .A2(new_n1008), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(new_n773), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1142), .A2(new_n1143), .B1(new_n1054), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1126), .A2(KEYINPUT120), .A3(new_n1008), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n556), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1140), .B(new_n1141), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1133), .A2(KEYINPUT60), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1133), .A2(KEYINPUT60), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT122), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n616), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(KEYINPUT122), .A3(new_n626), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1154), .A2(KEYINPUT122), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1136), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n991), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1162), .A2(KEYINPUT124), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(KEYINPUT124), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1092), .A2(new_n1107), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1105), .C1(new_n1109), .C2(KEYINPUT53), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(G171), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(KEYINPUT54), .C1(G171), .C2(new_n1110), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT125), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1166), .A2(G171), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(G171), .B2(new_n1110), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1170), .B(new_n1103), .C1(new_n1172), .C2(KEYINPUT54), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1125), .B1(new_n1161), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT113), .B1(G290), .B2(G1986), .ZN(new_n1176));
  NAND2_X1  g751(.A1(G290), .A2(G1986), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1176), .B(new_n1177), .Z(new_n1178));
  NOR2_X1   g753(.A1(new_n1000), .A2(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1024), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1033), .B1(new_n1175), .B2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g756(.A1(new_n906), .A2(new_n903), .ZN(new_n1183));
  INV_X1    g757(.A(new_n985), .ZN(new_n1184));
  OR4_X1    g758(.A1(new_n458), .A2(G401), .A3(G227), .A4(G229), .ZN(new_n1185));
  NOR3_X1   g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(G308));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n900), .B2(new_n904), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1187), .A2(new_n985), .ZN(G225));
endmodule


