//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  NOR2_X1   g000(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(KEYINPUT78), .A3(G125), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(KEYINPUT16), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n188), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AOI211_X1 g016(.A(new_n201), .B(new_n188), .C1(new_n196), .C2(new_n198), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n190), .A2(new_n192), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n188), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT77), .A3(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT77), .B1(new_n207), .B2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT24), .B(G110), .Z(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n207), .A2(G128), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(KEYINPUT23), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n213), .A2(new_n214), .B1(new_n218), .B2(G110), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n202), .A2(new_n204), .A3(new_n206), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(new_n214), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(G110), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n196), .A2(new_n188), .A3(new_n198), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n200), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT70), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G953), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n220), .A2(new_n226), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n234), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n199), .A2(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n219), .A2(new_n206), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n237), .A2(new_n238), .A3(new_n203), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n236), .B1(new_n239), .B2(new_n225), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n187), .B1(new_n241), .B2(G902), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  INV_X1    g057(.A(new_n187), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n235), .A2(new_n240), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n242), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G217), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(G234), .B2(new_n243), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(G902), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT81), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n240), .A2(new_n235), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G128), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT65), .B(G143), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n258), .B(new_n260), .C1(new_n261), .C2(G146), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(G128), .B1(new_n258), .B2(new_n259), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G143), .ZN(new_n267));
  AOI21_X1  g081(.A(G146), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT66), .B1(new_n188), .B2(G143), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n257), .A3(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT68), .B(new_n264), .C1(new_n268), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n269), .B(new_n271), .C1(new_n261), .C2(G146), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT68), .B1(new_n275), .B2(new_n264), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n263), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT67), .B(G137), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G134), .ZN(new_n279));
  INV_X1    g093(.A(G134), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G137), .ZN(new_n281));
  OAI21_X1  g095(.A(G131), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(KEYINPUT11), .A3(G134), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  INV_X1    g098(.A(G137), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT11), .B1(new_n285), .B2(G134), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n280), .B2(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n277), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT2), .B(G113), .Z(new_n292));
  XNOR2_X1  g106(.A(G116), .B(G119), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT0), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT64), .B1(new_n296), .B2(new_n209), .ZN(new_n297));
  OR3_X1    g111(.A1(new_n296), .A2(new_n209), .A3(KEYINPUT64), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n209), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n275), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n258), .B1(new_n261), .B2(G146), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT0), .A3(G128), .ZN(new_n302));
  INV_X1    g116(.A(new_n288), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n284), .B1(new_n283), .B2(new_n287), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n300), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n291), .A2(new_n295), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n264), .B1(new_n268), .B2(new_n272), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n262), .B1(new_n310), .B2(new_n273), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n305), .B(KEYINPUT30), .C1(new_n311), .C2(new_n289), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n277), .A2(KEYINPUT69), .A3(new_n290), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n311), .B2(new_n289), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n305), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n307), .B1(new_n319), .B2(new_n294), .ZN(new_n320));
  INV_X1    g134(.A(G237), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n231), .A2(G210), .A3(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G101), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n324), .B(new_n325), .Z(new_n326));
  OAI21_X1  g140(.A(new_n256), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n317), .A2(new_n318), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n294), .A3(new_n312), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n306), .ZN(new_n330));
  INV_X1    g144(.A(new_n326), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(KEYINPUT74), .A3(new_n331), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n317), .A2(new_n336), .A3(new_n294), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n306), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n317), .B2(new_n294), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT28), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n307), .A2(KEYINPUT28), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n326), .B(KEYINPUT72), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n333), .A2(new_n334), .A3(new_n335), .A4(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n335), .A3(new_n327), .A4(new_n332), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n291), .A2(new_n305), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n294), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n306), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(KEYINPUT76), .A3(new_n294), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT28), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT29), .A3(new_n341), .A4(new_n326), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n243), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n345), .A2(new_n347), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G472), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n340), .A2(new_n341), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n329), .A2(new_n306), .A3(new_n326), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT31), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n320), .A2(KEYINPUT31), .A3(new_n326), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n359), .A2(new_n342), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G472), .A2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT32), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n362), .A2(new_n363), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n343), .B1(new_n340), .B2(new_n341), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n368), .B(new_n365), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n255), .B1(new_n358), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G110), .B(G122), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n376), .A2(new_n379), .A3(new_n383), .A4(new_n380), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n386), .A3(G101), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n294), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n389));
  INV_X1    g203(.A(G116), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n390), .A2(KEYINPUT5), .A3(G119), .ZN(new_n391));
  INV_X1    g205(.A(G113), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n389), .A2(new_n393), .B1(new_n292), .B2(new_n293), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n378), .A2(G104), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n375), .A2(G107), .ZN(new_n396));
  OAI21_X1  g210(.A(G101), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n384), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n388), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n374), .B1(new_n400), .B2(KEYINPUT88), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n402), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT89), .A2(KEYINPUT6), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n403), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n399), .A4(new_n374), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI211_X1 g223(.A(G125), .B(new_n262), .C1(new_n310), .C2(new_n273), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n191), .B1(new_n300), .B2(new_n302), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT90), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n311), .A2(new_n191), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  INV_X1    g228(.A(new_n411), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n227), .A2(G224), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n412), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n412), .B2(new_n416), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n409), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT7), .ZN(new_n423));
  OAI22_X1  g237(.A1(new_n410), .A2(new_n411), .B1(new_n423), .B2(new_n418), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n374), .B(KEYINPUT8), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n394), .A2(new_n398), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n394), .A2(new_n398), .A3(KEYINPUT91), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT91), .B1(new_n394), .B2(new_n398), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n418), .A2(new_n423), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n413), .A2(new_n415), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n388), .A2(new_n399), .A3(new_n374), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n424), .A2(new_n430), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n243), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n422), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n422), .A2(new_n438), .A3(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n231), .A2(G227), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G140), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n301), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(KEYINPUT1), .C1(new_n261), .C2(G146), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n265), .A2(new_n267), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n188), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n454), .B2(KEYINPUT1), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n449), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n263), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT10), .B1(new_n457), .B2(new_n398), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n300), .A2(new_n385), .A3(new_n302), .A4(new_n387), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n398), .A2(KEYINPUT10), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n311), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT87), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n303), .A2(new_n304), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT10), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT85), .B1(new_n268), .B2(new_n259), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(G128), .A3(new_n451), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n262), .B1(new_n467), .B2(new_n449), .ZN(new_n468));
  INV_X1    g282(.A(new_n398), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  INV_X1    g285(.A(new_n460), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n277), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n470), .A2(new_n471), .A3(new_n459), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n462), .A2(new_n464), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n470), .A2(new_n463), .A3(new_n459), .A4(new_n473), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n448), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n448), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n310), .A2(new_n273), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n263), .A3(new_n469), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n469), .B2(new_n468), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT12), .B1(new_n481), .B2(new_n464), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n468), .A2(new_n469), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n262), .B(new_n398), .C1(new_n310), .C2(new_n273), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT12), .B(new_n464), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n478), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n445), .B(new_n243), .C1(new_n477), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n478), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n476), .A2(KEYINPUT86), .A3(new_n448), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n475), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n486), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n476), .B1(new_n493), .B2(new_n482), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n448), .B(KEYINPUT84), .Z(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n496), .A3(G469), .ZN(new_n497));
  NAND2_X1  g311(.A1(G469), .A2(G902), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n488), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT9), .B(G234), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT82), .ZN(new_n501));
  OAI21_X1  g315(.A(G221), .B1(new_n501), .B2(G902), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT83), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT97), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n265), .A2(new_n267), .A3(G128), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n257), .A2(G128), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n506), .A2(new_n280), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n511));
  INV_X1    g325(.A(G122), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(G116), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n390), .A2(KEYINPUT94), .A3(G122), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(G116), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n378), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n378), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n510), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g334(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n506), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT96), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n506), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n508), .B1(new_n521), .B2(new_n506), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n520), .B1(new_n529), .B2(G134), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n515), .A2(KEYINPUT14), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n515), .A2(KEYINPUT14), .B1(G116), .B2(new_n512), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n378), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n280), .B1(new_n506), .B2(new_n508), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n517), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n501), .A2(new_n248), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n530), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n536), .ZN(new_n540));
  INV_X1    g354(.A(new_n519), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n509), .B1(new_n541), .B2(new_n517), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n527), .B1(new_n523), .B2(new_n525), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n280), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n537), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n243), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n538), .B1(new_n530), .B2(new_n536), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n540), .A2(new_n544), .A3(new_n537), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n548), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n505), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n548), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n553), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT97), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G475), .A2(G902), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n231), .A2(G143), .A3(G214), .A4(new_n321), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n228), .A2(new_n230), .A3(G214), .A4(new_n321), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n261), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G131), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n284), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n224), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(new_n199), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(KEYINPUT17), .A3(G131), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(G113), .B(G122), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(new_n375), .ZN(new_n574));
  AND2_X1   g388(.A1(KEYINPUT18), .A2(G131), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n561), .A2(new_n575), .A3(new_n563), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n561), .B2(new_n563), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n578), .A2(new_n206), .A3(KEYINPUT92), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT92), .B1(new_n578), .B2(new_n206), .ZN(new_n580));
  OAI22_X1  g394(.A1(new_n576), .A2(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n572), .A2(new_n574), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n194), .A2(new_n195), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(KEYINPUT19), .B2(new_n205), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n565), .A2(new_n567), .B1(new_n586), .B2(new_n188), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n237), .A2(new_n203), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n574), .B1(new_n589), .B2(new_n581), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n560), .B1(new_n583), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT20), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n576), .A2(new_n577), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n579), .A2(new_n580), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n588), .A2(new_n587), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n582), .B1(new_n595), .B2(new_n574), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT20), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n560), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n572), .A2(new_n581), .ZN(new_n599));
  INV_X1    g413(.A(new_n574), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT93), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n582), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n574), .B1(new_n572), .B2(new_n581), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n243), .B(new_n601), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n592), .A2(new_n598), .B1(new_n605), .B2(G475), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n227), .A2(G952), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(G234), .B2(G237), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n243), .B(new_n231), .C1(G234), .C2(G237), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT21), .B(G898), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT98), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n559), .A2(new_n606), .A3(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n444), .A2(new_n504), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n373), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  OAI21_X1  g430(.A(G472), .B1(new_n364), .B2(G902), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n499), .A2(new_n503), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n359), .A2(new_n342), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n362), .A2(new_n363), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n365), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n617), .A2(new_n618), .A3(new_n622), .A4(new_n254), .ZN(new_n623));
  INV_X1    g437(.A(new_n443), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n440), .B2(new_n441), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n546), .A2(new_n626), .A3(new_n547), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT100), .B1(new_n552), .B2(G478), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n630), .B(new_n631), .C1(new_n539), .C2(new_n545), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT99), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n547), .A2(G902), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n627), .A2(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n606), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n625), .A2(new_n612), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n623), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT34), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NAND3_X1  g455(.A1(new_n442), .A2(new_n443), .A3(new_n612), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n597), .B1(new_n596), .B2(new_n560), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n643), .A2(KEYINPUT101), .B1(new_n605), .B2(G475), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n592), .A2(new_n598), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n644), .A2(new_n646), .A3(new_n558), .A4(new_n555), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n623), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n378), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  INV_X1    g465(.A(new_n613), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT103), .B1(new_n239), .B2(new_n225), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n654));
  OR3_X1    g468(.A1(new_n239), .A2(KEYINPUT103), .A3(new_n225), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n653), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n252), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n250), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n618), .A2(new_n625), .A3(new_n652), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n617), .A2(new_n622), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT37), .B(G110), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  AOI22_X1  g480(.A1(new_n357), .A2(G472), .B1(new_n367), .B2(new_n371), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n438), .B1(new_n422), .B2(new_n436), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n439), .B(new_n435), .C1(new_n409), .C2(new_n421), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n659), .B(new_n443), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n609), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n608), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n647), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n671), .A2(new_n618), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT106), .B1(new_n667), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n676), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n367), .A2(new_n371), .ZN(new_n680));
  INV_X1    g494(.A(G472), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n355), .B1(new_n346), .B2(KEYINPUT75), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n681), .B1(new_n682), .B2(new_n345), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n674), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n618), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n668), .A2(new_n669), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n659), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n559), .A2(new_n606), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n443), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n342), .A2(new_n352), .A3(new_n351), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n360), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n681), .B1(new_n698), .B2(new_n243), .ZN(new_n699));
  AOI211_X1 g513(.A(KEYINPUT108), .B(new_n699), .C1(new_n367), .C2(new_n371), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n701));
  INV_X1    g515(.A(new_n699), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n701), .B1(new_n372), .B2(new_n702), .ZN(new_n703));
  OAI221_X1 g517(.A(new_n696), .B1(KEYINPUT40), .B2(new_n688), .C1(new_n700), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n453), .ZN(G45));
  NAND2_X1  g519(.A1(new_n358), .A2(new_n372), .ZN(new_n706));
  INV_X1    g520(.A(new_n636), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n592), .A2(new_n598), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n605), .A2(G475), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n674), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n670), .A2(new_n504), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  OAI21_X1  g529(.A(new_n243), .B1(new_n477), .B2(new_n487), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n503), .A3(new_n488), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n638), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n254), .B(new_n719), .C1(new_n680), .C2(new_n683), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NOR3_X1   g536(.A1(new_n642), .A2(new_n718), .A3(new_n647), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n254), .B(new_n723), .C1(new_n680), .C2(new_n683), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR3_X1   g539(.A1(new_n670), .A2(new_n718), .A3(new_n613), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n680), .B2(new_n683), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n729));
  AOI21_X1  g543(.A(G902), .B1(new_n619), .B2(new_n620), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n729), .B1(new_n730), .B2(new_n681), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT109), .B(G472), .C1(new_n364), .C2(G902), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n625), .A2(new_n694), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n717), .A2(new_n503), .A3(new_n488), .A4(new_n612), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n353), .A2(new_n341), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n342), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n366), .B1(new_n620), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n733), .A2(new_n254), .A3(new_n736), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n739), .B1(new_n731), .B2(new_n732), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT110), .A3(new_n254), .A4(new_n736), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NOR3_X1   g561(.A1(new_n670), .A2(new_n718), .A3(new_n712), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n621), .A2(new_n243), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT109), .B1(new_n749), .B2(G472), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n730), .A2(new_n729), .A3(new_n681), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n740), .B(new_n748), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  NAND4_X1  g567(.A1(new_n690), .A2(new_n637), .A3(new_n443), .A4(new_n711), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n498), .B(KEYINPUT111), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n488), .A2(new_n497), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n503), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n759), .A3(new_n503), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n754), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(new_n254), .C1(new_n680), .C2(new_n683), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n706), .A2(KEYINPUT42), .A3(new_n254), .A4(new_n761), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND3_X1  g581(.A1(new_n440), .A2(new_n443), .A3(new_n441), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n758), .A2(new_n760), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n373), .A2(new_n675), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT113), .B(G134), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G36));
  AOI211_X1 g587(.A(KEYINPUT43), .B(new_n710), .C1(KEYINPUT114), .C2(new_n707), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(KEYINPUT114), .B2(new_n707), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n636), .B1(new_n710), .B2(KEYINPUT115), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(KEYINPUT115), .B2(new_n710), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT43), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n661), .A3(new_n659), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n768), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n492), .A2(new_n496), .A3(KEYINPUT45), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT45), .B1(new_n492), .B2(new_n496), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n445), .ZN(new_n785));
  INV_X1    g599(.A(new_n755), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n488), .B1(new_n787), .B2(KEYINPUT46), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n503), .B(new_n687), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n782), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n285), .ZN(G39));
  NOR3_X1   g606(.A1(new_n706), .A2(new_n254), .A3(new_n754), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n503), .B1(new_n788), .B2(new_n789), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n793), .A2(new_n794), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  AND3_X1   g615(.A1(new_n775), .A2(new_n608), .A3(new_n778), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n718), .A2(new_n768), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n373), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n607), .B(KEYINPUT121), .Z(new_n808));
  NAND2_X1  g622(.A1(new_n733), .A2(new_n740), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n255), .ZN(new_n810));
  INV_X1    g624(.A(new_n718), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n802), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n707), .A2(new_n710), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n703), .A2(new_n700), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n254), .A3(new_n608), .A4(new_n803), .ZN(new_n815));
  OAI221_X1 g629(.A(new_n808), .B1(new_n812), .B2(new_n444), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n807), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n692), .A2(new_n624), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n812), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n818), .B1(new_n812), .B2(new_n819), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n815), .A2(new_n710), .A3(new_n707), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n804), .A2(new_n693), .A3(new_n809), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n810), .A2(new_n802), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n717), .A2(new_n488), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n503), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n769), .B(new_n827), .C1(new_n798), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT51), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n817), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n822), .A2(new_n825), .A3(KEYINPUT120), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n830), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n677), .A2(new_n684), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n693), .A2(new_n711), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n734), .A2(new_n841), .A3(new_n757), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n703), .B2(new_n700), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n714), .A3(new_n752), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n839), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n372), .A2(new_n702), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT108), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n372), .A2(new_n701), .A3(new_n702), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n713), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n752), .B1(new_n667), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n685), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n720), .A2(new_n724), .A3(new_n727), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n766), .A2(new_n857), .A3(new_n746), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n744), .A2(new_n761), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n549), .A2(new_n554), .A3(new_n674), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n644), .A2(new_n646), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n768), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n644), .A2(new_n646), .A3(new_n861), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n690), .A3(KEYINPUT117), .A4(new_n443), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n865), .A3(new_n618), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n358), .B2(new_n372), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n659), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n606), .B1(new_n554), .B2(new_n549), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n813), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n625), .A3(new_n612), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n623), .A2(new_n871), .B1(new_n660), .B2(new_n661), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n373), .B2(new_n614), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n868), .A2(new_n873), .A3(new_n771), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n858), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT53), .B1(new_n856), .B2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n840), .A2(new_n844), .A3(new_n839), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT52), .B1(new_n853), .B2(new_n685), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT118), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n845), .A2(new_n854), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(KEYINPUT54), .B(new_n877), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT53), .B1(new_n855), .B2(new_n875), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n880), .A2(new_n882), .ZN(new_n888));
  AND4_X1   g702(.A1(KEYINPUT53), .A2(new_n766), .A3(new_n857), .A4(new_n746), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n868), .A2(new_n873), .A3(KEYINPUT119), .A4(new_n771), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n874), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n887), .B1(new_n888), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n838), .A2(new_n886), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n254), .A2(new_n503), .A3(new_n443), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n777), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n828), .B(KEYINPUT49), .Z(new_n902));
  NAND4_X1  g716(.A1(new_n814), .A2(new_n692), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(G75));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n895), .B2(new_n243), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n893), .B1(new_n882), .B2(new_n880), .ZN(new_n907));
  OAI211_X1 g721(.A(KEYINPUT123), .B(G902), .C1(new_n907), .C2(new_n887), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n439), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n409), .B(new_n421), .ZN(new_n910));
  XOR2_X1   g724(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT124), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n231), .A2(G952), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT125), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(G210), .B(G902), .C1(new_n907), .C2(new_n887), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n921), .B2(new_n912), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n915), .A2(new_n922), .ZN(G51));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n907), .B2(new_n887), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n897), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n755), .B(KEYINPUT57), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n477), .A2(new_n487), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n906), .A2(new_n785), .A3(new_n908), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n918), .B1(new_n929), .B2(new_n930), .ZN(G54));
  AND3_X1   g745(.A1(new_n596), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n906), .A2(new_n908), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n917), .ZN(new_n934));
  INV_X1    g748(.A(new_n596), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n906), .A2(new_n908), .A3(KEYINPUT58), .A4(G475), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(G60));
  NAND2_X1  g751(.A1(new_n897), .A2(new_n886), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n634), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n634), .A2(new_n941), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n897), .B2(new_n924), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n942), .A2(new_n918), .A3(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI221_X1 g762(.A(new_n948), .B1(new_n656), .B2(new_n657), .C1(new_n907), .C2(new_n887), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n241), .B1(new_n895), .B2(new_n947), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n950), .A3(new_n917), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G66));
  INV_X1    g767(.A(new_n610), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n227), .B1(new_n954), .B2(G224), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n857), .A2(new_n746), .A3(new_n873), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n231), .ZN(new_n957));
  INV_X1    g771(.A(new_n409), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(G898), .B2(new_n231), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT126), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n957), .B(new_n960), .ZN(G69));
  AOI21_X1  g775(.A(new_n231), .B1(G227), .B2(G900), .ZN(new_n962));
  INV_X1    g776(.A(new_n791), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n800), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n840), .A2(new_n852), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n704), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n769), .A2(new_n870), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n805), .A2(new_n688), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT127), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n964), .A2(new_n967), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n972), .A2(new_n231), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n319), .B(new_n586), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n771), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n805), .A2(new_n790), .A3(new_n734), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n791), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(new_n766), .A3(new_n800), .A4(new_n965), .ZN(new_n979));
  INV_X1    g793(.A(new_n231), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(G900), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n974), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n962), .B1(new_n975), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n962), .ZN(new_n986));
  OAI221_X1 g800(.A(new_n986), .B1(new_n981), .B2(new_n983), .C1(new_n973), .C2(new_n974), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G72));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n972), .B2(new_n956), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n326), .A3(new_n330), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n333), .A2(new_n360), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n993), .A2(new_n990), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n877), .B(new_n994), .C1(new_n883), .C2(new_n885), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n990), .B1(new_n979), .B2(new_n956), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n330), .A2(new_n326), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n918), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n992), .A2(new_n995), .A3(new_n998), .ZN(G57));
endmodule


