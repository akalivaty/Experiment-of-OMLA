//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G137), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n460), .B2(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n467), .B1(new_n470), .B2(new_n461), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n468), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n471), .B2(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n461), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n461), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n472), .A2(new_n473), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n460), .A2(KEYINPUT68), .A3(new_n461), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n484), .B1(new_n489), .B2(G136), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(KEYINPUT71), .C1(new_n473), .C2(new_n472), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(KEYINPUT70), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n461), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n480), .A2(G126), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n461), .A2(G138), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n502), .B1(new_n478), .B2(new_n479), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n503), .B2(KEYINPUT71), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n493), .B(new_n501), .C1(new_n473), .C2(new_n472), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n496), .B(new_n500), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n520), .A2(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n516), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NOR2_X1   g105(.A1(new_n523), .A2(new_n522), .ZN(new_n531));
  OAI21_X1  g106(.A(G89), .B1(new_n524), .B2(new_n525), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n537), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g114(.A(G51), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n534), .A2(new_n541), .ZN(G168));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n543));
  OAI211_X1 g118(.A(G52), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n526), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(G64), .B1(new_n523), .B2(new_n522), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n515), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n543), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n511), .B2(new_n512), .ZN(new_n552));
  INV_X1    g127(.A(new_n548), .ZN(new_n553));
  OAI21_X1  g128(.A(G651), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n519), .A2(new_n513), .A3(G90), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n554), .A2(KEYINPUT72), .A3(new_n544), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n550), .A2(new_n556), .ZN(G171));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  INV_X1    g133(.A(G68), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n531), .A2(new_n558), .B1(new_n559), .B2(new_n510), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI221_X1 g137(.A(KEYINPUT73), .B1(new_n559), .B2(new_n510), .C1(new_n531), .C2(new_n558), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(G651), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n526), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(G81), .B1(G43), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  XOR2_X1   g149(.A(KEYINPUT74), .B(KEYINPUT9), .Z(new_n575));
  NAND3_X1  g150(.A1(new_n566), .A2(new_n575), .A3(G53), .ZN(new_n576));
  INV_X1    g151(.A(G91), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n576), .A2(KEYINPUT75), .B1(new_n577), .B2(new_n526), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n511), .A2(new_n579), .A3(new_n512), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n579), .B1(new_n511), .B2(new_n512), .ZN(new_n582));
  OAI21_X1  g157(.A(G65), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n578), .B1(new_n585), .B2(G651), .ZN(new_n586));
  INV_X1    g161(.A(G53), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT9), .B1(new_n520), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(KEYINPUT75), .A3(new_n576), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(G299));
  INV_X1    g165(.A(G171), .ZN(G301));
  INV_X1    g166(.A(G168), .ZN(G286));
  OAI21_X1  g167(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  INV_X1    g169(.A(G49), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n526), .B2(new_n594), .C1(new_n595), .C2(new_n520), .ZN(G288));
  AOI22_X1  g171(.A1(new_n565), .A2(G86), .B1(G48), .B2(new_n566), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n513), .A2(G61), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n515), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(KEYINPUT77), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  AOI211_X1 g177(.A(new_n602), .B(new_n515), .C1(new_n598), .C2(new_n599), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n597), .B1(new_n601), .B2(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n515), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT78), .B(G47), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n520), .A2(new_n607), .B1(new_n526), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G290));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(G301), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n513), .A2(KEYINPUT76), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n580), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT79), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(G66), .B1(new_n581), .B2(new_n582), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(new_n621), .A3(new_n617), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n619), .A2(new_n622), .A3(G651), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n565), .A2(KEYINPUT10), .A3(G92), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n526), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n624), .A2(new_n627), .B1(G54), .B2(new_n566), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n613), .B1(new_n632), .B2(new_n612), .ZN(G284));
  AOI21_X1  g208(.A(new_n613), .B1(new_n632), .B2(new_n612), .ZN(G321));
  NAND2_X1  g209(.A1(G299), .A2(new_n612), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g211(.A(new_n635), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n632), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n568), .A2(new_n612), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n631), .A2(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n480), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n461), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n489), .B2(G135), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT82), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n460), .A2(new_n464), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT13), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n658), .B(new_n660), .Z(new_n661));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n661), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT84), .ZN(new_n674));
  NOR2_X1   g249(.A1(G2072), .A2(G2078), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n442), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n676), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(KEYINPUT17), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n678), .C1(new_n674), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n674), .A2(new_n682), .A3(new_n677), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT85), .ZN(new_n691));
  XOR2_X1   g266(.A(G1971), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(KEYINPUT85), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n688), .A2(new_n689), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(new_n690), .ZN(new_n698));
  MUX2_X1   g273(.A(new_n698), .B(new_n697), .S(new_n693), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT86), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G32), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n489), .A2(G141), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n464), .A2(G105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT89), .Z(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n480), .A2(G129), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n710), .B1(new_n718), .B2(new_n709), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT27), .B(G1996), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n719), .A2(new_n721), .B1(new_n649), .B2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT31), .B(G11), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT90), .ZN(new_n725));
  INV_X1    g300(.A(G28), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n726), .B2(KEYINPUT30), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(KEYINPUT30), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G21), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G168), .B2(new_n730), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n729), .B1(new_n732), .B2(G1966), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G1966), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n709), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  AOI22_X1  g312(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n487), .A2(new_n488), .ZN(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n737), .B1(new_n461), .B2(new_n738), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n735), .B1(new_n742), .B2(new_n709), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2072), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n723), .A2(new_n734), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n709), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n709), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT29), .ZN(new_n748));
  INV_X1    g323(.A(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(KEYINPUT29), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G5), .A2(G16), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G171), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n709), .A2(G27), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT91), .Z(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n507), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2078), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n745), .A2(new_n751), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n730), .A2(G19), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n569), .B2(new_n730), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT88), .ZN(new_n764));
  INV_X1    g339(.A(G1341), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n709), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n480), .A2(G128), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n461), .A2(G116), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G140), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n769), .B1(new_n770), .B2(new_n771), .C1(new_n739), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n777));
  INV_X1    g352(.A(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G160), .B2(new_n709), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(G2084), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(G2084), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n776), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n764), .A2(new_n765), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n730), .A2(G20), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT23), .Z(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1956), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n766), .A2(new_n784), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n761), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n730), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n632), .B2(new_n730), .ZN(new_n795));
  INV_X1    g370(.A(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n792), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n793), .B1(new_n792), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n730), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n730), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G6), .B(G305), .S(G16), .Z(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT32), .B(G1981), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n730), .A2(G23), .ZN(new_n809));
  INV_X1    g384(.A(G288), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n730), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT33), .B(G1976), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n804), .A2(new_n807), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n489), .A2(G131), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n818));
  INV_X1    g393(.A(G107), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G2105), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G119), .B2(new_n480), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G29), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G25), .B2(G29), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  AND2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n730), .A2(G24), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n610), .B2(new_n730), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(G1986), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n829), .A2(G1986), .ZN(new_n831));
  NOR4_X1   g406(.A1(new_n826), .A2(new_n827), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n815), .A2(new_n816), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT87), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT87), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n815), .A2(new_n835), .A3(new_n816), .A4(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(KEYINPUT36), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n800), .A2(new_n841), .ZN(G311));
  OR2_X1    g417(.A1(new_n800), .A2(new_n841), .ZN(G150));
  NAND2_X1  g418(.A1(new_n632), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n515), .ZN(new_n847));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n520), .A2(new_n848), .B1(new_n526), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n568), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n564), .A3(new_n567), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n845), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  NAND2_X1  g437(.A1(new_n489), .A2(G142), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  INV_X1    g439(.A(G118), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(G2105), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G130), .B2(new_n480), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n653), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n817), .A2(new_n821), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT93), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(KEYINPUT93), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n653), .A3(new_n871), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n868), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n876), .A3(new_n868), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n879), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n874), .A2(new_n876), .A3(new_n868), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n877), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n773), .A2(new_n507), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n773), .A2(new_n507), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(new_n741), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n741), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n718), .ZN(new_n891));
  OR3_X1    g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n885), .A2(new_n886), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G162), .B(G160), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n649), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n895), .B1(new_n885), .B2(new_n886), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n898), .B1(new_n885), .B2(new_n894), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n881), .A3(new_n884), .ZN(new_n903));
  AOI21_X1  g478(.A(G37), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT40), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT40), .B1(new_n901), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(G395));
  NAND2_X1  g482(.A1(new_n629), .A2(G299), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n623), .A2(new_n586), .A3(new_n589), .A4(new_n628), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT41), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n855), .B(KEYINPUT97), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n641), .B(new_n915), .ZN(new_n916));
  MUX2_X1   g491(.A(new_n911), .B(new_n914), .S(new_n916), .Z(new_n917));
  XNOR2_X1  g492(.A(G305), .B(G303), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n810), .B(new_n610), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n919), .A2(KEYINPUT98), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(KEYINPUT98), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n918), .B2(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(KEYINPUT42), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n925), .B(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n917), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n917), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(G868), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n852), .A2(new_n612), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(G295));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n932), .ZN(G331));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n550), .A2(G168), .A3(new_n556), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(KEYINPUT101), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n550), .A2(new_n556), .A3(new_n938), .A4(G168), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(G171), .B2(G286), .ZN(new_n942));
  AOI211_X1 g517(.A(KEYINPUT102), .B(G168), .C1(new_n550), .C2(new_n556), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n937), .A2(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n855), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n936), .A2(KEYINPUT101), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n939), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n855), .B(new_n949), .C1(new_n942), .C2(new_n943), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n944), .A2(KEYINPUT103), .A3(new_n945), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n910), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(KEYINPUT104), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n944), .A2(new_n955), .A3(new_n945), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n950), .A3(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n953), .A2(KEYINPUT106), .B1(new_n957), .B2(new_n914), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n951), .A2(new_n952), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n910), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n923), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n951), .A2(new_n914), .A3(new_n952), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n954), .A2(new_n911), .A3(new_n950), .A4(new_n956), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n923), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n964), .ZN(new_n969));
  INV_X1    g544(.A(new_n923), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n966), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n923), .B1(new_n963), .B2(new_n964), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT105), .B1(new_n974), .B2(G37), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n975), .A3(new_n976), .A4(new_n965), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n935), .B1(new_n968), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n965), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n969), .B2(new_n970), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n980), .B2(new_n972), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n976), .B1(new_n981), .B2(new_n975), .ZN(new_n982));
  INV_X1    g557(.A(new_n976), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n962), .A2(new_n983), .A3(new_n967), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n978), .B1(new_n985), .B2(new_n935), .ZN(G397));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT45), .B1(new_n507), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n989), .B(new_n466), .C1(new_n471), .C2(new_n476), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n891), .A2(G1996), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n773), .B(new_n775), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n991), .A2(G1996), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n718), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n991), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n822), .A2(new_n825), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n822), .A2(new_n825), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n610), .B(G1986), .Z(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n597), .ZN(new_n1007));
  OAI21_X1  g582(.A(G1981), .B1(new_n1007), .B2(new_n600), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(G305), .B2(G1981), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(KEYINPUT110), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n1012));
  OAI221_X1 g587(.A(new_n1008), .B1(new_n1012), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n507), .A2(new_n987), .ZN(new_n1014));
  INV_X1    g589(.A(new_n466), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT67), .B1(new_n475), .B2(G2105), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n467), .B(new_n461), .C1(new_n474), .C2(new_n468), .ZN(new_n1017));
  OAI211_X1 g592(.A(G40), .B(new_n1015), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT109), .B(G8), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1011), .A2(new_n1013), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n810), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(G1981), .B2(G305), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n1021), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n810), .A2(G1976), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1021), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1029), .A2(new_n1022), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT55), .Z(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(new_n990), .C1(new_n988), .C2(KEYINPUT108), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n1038), .B(KEYINPUT45), .C1(new_n507), .C2(new_n987), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n803), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n507), .A2(new_n1041), .A3(new_n987), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n507), .B2(new_n987), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1018), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n749), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1035), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1032), .A2(new_n1034), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1026), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT63), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1034), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1043), .A2(new_n1018), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1042), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT111), .B1(new_n1043), .B2(new_n1018), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n749), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1020), .B1(new_n1055), .B2(new_n1040), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1032), .B(new_n1050), .C1(new_n1056), .C2(new_n1034), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n507), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n987), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n500), .A2(new_n496), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(KEYINPUT4), .A3(new_n505), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1059), .B(new_n990), .C1(new_n1063), .C2(KEYINPUT45), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1036), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1058), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT113), .B(G2084), .Z(new_n1068));
  NAND2_X1  g643(.A1(new_n1044), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1020), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(G168), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1049), .B1(new_n1057), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1049), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1046), .A2(new_n1034), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1050), .A4(new_n1032), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1048), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT45), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1014), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1038), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1018), .B1(new_n1063), .B2(KEYINPUT45), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n988), .A2(KEYINPUT108), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n758), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1042), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1051), .A2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT122), .B(G1961), .Z(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n988), .A2(new_n1018), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1036), .A2(new_n1065), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1084), .A2(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1059), .A4(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1085), .A2(G301), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT54), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n475), .A2(G2105), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1015), .A2(new_n1097), .A3(G40), .A4(new_n1093), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n988), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1083), .A2(new_n1084), .B1(new_n1036), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1044), .B2(new_n1088), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1087), .A2(KEYINPUT123), .A3(new_n1089), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(G301), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1096), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n1057), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1100), .A2(new_n1104), .A3(G301), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1110), .B2(new_n1085), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G168), .A2(new_n1020), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1092), .A2(new_n1079), .A3(new_n1059), .A4(new_n990), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1058), .A2(new_n1115), .B1(new_n1044), .B2(new_n1068), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1116), .B2(new_n1035), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1070), .A2(G286), .A3(new_n1071), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(KEYINPUT51), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1116), .B2(new_n1020), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1119), .A2(KEYINPUT121), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT121), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1107), .B(new_n1112), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1037), .A2(new_n1039), .A3(G1996), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n1126), .C1(new_n1014), .C2(new_n1018), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n569), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT120), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n569), .B(new_n1134), .C1(new_n1125), .C2(new_n1131), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1087), .A2(new_n796), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1019), .A2(new_n775), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n629), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1138), .A3(new_n1139), .A4(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1136), .A2(new_n1137), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(G299), .B(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT114), .B(G1956), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT56), .B(G2072), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT116), .Z(new_n1154));
  NAND4_X1  g729(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1150), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n990), .B(new_n1052), .C1(new_n1063), .C2(new_n1041), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(new_n1054), .A3(new_n1086), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1151), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT61), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1157), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1146), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1149), .B1(new_n1161), .B2(new_n1155), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n629), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1162), .B(KEYINPUT117), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1167), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1077), .B1(new_n1124), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1035), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT51), .B1(new_n1178), .B2(new_n1113), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1116), .A2(G168), .A3(new_n1020), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1121), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1119), .A2(KEYINPUT121), .A3(new_n1121), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1110), .A2(new_n1085), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1057), .A2(G301), .A3(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1177), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1006), .B1(new_n1176), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1004), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n991), .A2(G1986), .A3(G290), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1192), .B(KEYINPUT48), .Z(new_n1193));
  NAND2_X1  g768(.A1(new_n995), .A2(KEYINPUT46), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT125), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n991), .B1(new_n993), .B2(new_n718), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n995), .A2(KEYINPUT46), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1195), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1203));
  AOI22_X1  g778(.A1(new_n1191), .A2(new_n1193), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n999), .A2(new_n1001), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n773), .A2(G2067), .ZN(new_n1206));
  OAI211_X1 g781(.A(KEYINPUT124), .B(new_n1000), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1206), .B1(new_n999), .B2(new_n1001), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1208), .B1(new_n1209), .B2(new_n991), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1204), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(KEYINPUT127), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1204), .A2(new_n1207), .A3(new_n1213), .A4(new_n1210), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1190), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g791(.A(G319), .ZN(new_n1218));
  NOR3_X1   g792(.A1(G401), .A2(new_n1218), .A3(G227), .ZN(new_n1219));
  INV_X1    g793(.A(new_n904), .ZN(new_n1220));
  NOR2_X1   g794(.A1(new_n899), .A2(new_n900), .ZN(new_n1221));
  OAI211_X1 g795(.A(new_n707), .B(new_n1219), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g796(.A1(new_n985), .A2(new_n1222), .ZN(G308));
  AND2_X1   g797(.A1(new_n707), .A2(new_n1219), .ZN(new_n1224));
  OAI221_X1 g798(.A(new_n1224), .B1(new_n1220), .B2(new_n1221), .C1(new_n982), .C2(new_n984), .ZN(G225));
endmodule


