//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1167, new_n1168, new_n1169, new_n1171,
    new_n1172, new_n1173, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n203), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n207), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n202), .A2(new_n203), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n210), .B1(new_n222), .B2(KEYINPUT1), .C1(new_n226), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT66), .B(G50), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n223), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G50), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n224), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(G20), .B2(new_n204), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n254), .A2(new_n223), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n258), .B1(G50), .B2(new_n252), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G222), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G223), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n275), .B1(new_n217), .B2(new_n273), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n223), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n285), .A3(G274), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n279), .A2(new_n285), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(G226), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G200), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n268), .B(new_n291), .C1(new_n292), .C2(new_n290), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n291), .B2(KEYINPUT69), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n293), .B(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n290), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n267), .B1(new_n297), .B2(G169), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n290), .A2(G179), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  XOR2_X1   g0101(.A(KEYINPUT15), .B(G87), .Z(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n260), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n259), .A2(new_n263), .B1(new_n224), .B2(new_n217), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n255), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n256), .A2(G77), .A3(new_n257), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n306), .B(new_n307), .C1(G77), .C2(new_n252), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n273), .A2(G232), .A3(new_n274), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n309), .B1(new_n219), .B2(new_n273), .C1(new_n276), .C2(new_n212), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n279), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n287), .B1(G244), .B2(new_n288), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT68), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n308), .B1(new_n315), .B2(G200), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n292), .B2(new_n315), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n308), .C1(G179), .C2(new_n315), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n296), .A2(new_n301), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n263), .A2(new_n201), .B1(new_n224), .B2(G68), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n260), .A2(new_n217), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n255), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT11), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT70), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(KEYINPUT70), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n328));
  OR3_X1    g0128(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n203), .B1(new_n251), .B2(G20), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n328), .A2(new_n329), .B1(new_n256), .B2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n326), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n283), .A2(new_n284), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n273), .A2(G232), .A3(G1698), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n273), .A2(G226), .A3(new_n274), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n286), .B1(new_n212), .B2(new_n334), .C1(new_n338), .C2(new_n283), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT13), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n341), .A2(KEYINPUT14), .B1(new_n344), .B2(new_n340), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n333), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n340), .A2(new_n292), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n340), .A2(G200), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n332), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(G58), .B(G68), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(G20), .B1(G159), .B2(new_n262), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT71), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G33), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n355), .A3(new_n269), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n357));
  AOI21_X1  g0157(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n271), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n356), .A2(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n352), .B1(new_n361), .B2(new_n203), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n266), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT71), .B(G33), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n224), .B(new_n271), .C1(new_n365), .C2(new_n269), .ZN(new_n366));
  OR2_X1    g0166(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n369));
  NOR2_X1   g0169(.A1(KEYINPUT3), .A2(G33), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n353), .A2(new_n355), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(KEYINPUT3), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n369), .B1(new_n372), .B2(new_n224), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT16), .B(new_n352), .C1(new_n368), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n259), .A2(new_n253), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT8), .B(G58), .Z(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n257), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n266), .A2(new_n252), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT73), .B(new_n376), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G274), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n281), .B2(new_n282), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n288), .A2(G232), .B1(new_n387), .B2(new_n285), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n270), .A2(new_n213), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n271), .B1(new_n365), .B2(new_n269), .ZN(new_n390));
  NOR2_X1   g0190(.A1(G223), .A2(G1698), .ZN(new_n391));
  INV_X1    g0191(.A(G226), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n388), .B1(new_n394), .B2(new_n283), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G169), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n286), .B1(new_n334), .B2(new_n234), .ZN(new_n397));
  INV_X1    g0197(.A(new_n389), .ZN(new_n398));
  INV_X1    g0198(.A(new_n393), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n372), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n400), .B2(new_n279), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G179), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n375), .A2(new_n385), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT18), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n388), .B(new_n292), .C1(new_n394), .C2(new_n283), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n401), .B2(G200), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n375), .A2(new_n406), .A3(new_n385), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n321), .A2(new_n350), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n390), .A2(G250), .A3(new_n274), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n371), .A2(G294), .ZN(new_n413));
  AND2_X1   g0213(.A1(G257), .A2(G1698), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n390), .A2(KEYINPUT77), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT77), .B1(new_n390), .B2(new_n414), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n412), .B(new_n413), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n283), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n412), .A2(new_n413), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(KEYINPUT78), .C1(new_n417), .C2(new_n416), .ZN(new_n422));
  INV_X1    g0222(.A(G45), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G1), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT5), .B(G41), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n279), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n420), .A2(new_n422), .B1(G264), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n387), .A2(new_n424), .A3(new_n425), .ZN(new_n428));
  AOI21_X1  g0228(.A(G169), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(new_n419), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n279), .A3(new_n422), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(G264), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n344), .A2(new_n431), .A3(new_n428), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n371), .A2(G116), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT23), .B1(new_n219), .B2(G20), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT23), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n437), .A2(new_n224), .A3(G107), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n435), .A2(G20), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n390), .A2(new_n224), .A3(G87), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n390), .A2(KEYINPUT76), .A3(new_n224), .A4(G87), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT22), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n273), .ZN(new_n445));
  OR4_X1    g0245(.A1(KEYINPUT22), .A2(new_n445), .A3(G20), .A4(new_n213), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n439), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT24), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(KEYINPUT24), .B(new_n439), .C1(new_n444), .C2(new_n446), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n255), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n253), .A2(new_n219), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT25), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n251), .A2(G33), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n266), .A2(new_n252), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT74), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT74), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n256), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n453), .B1(new_n460), .B2(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n451), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n434), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n224), .C1(G33), .C2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n255), .C1(new_n224), .C2(G116), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT20), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n253), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n455), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(G257), .A2(G1698), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n220), .B2(G1698), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n390), .A2(new_n475), .B1(G303), .B2(new_n445), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n283), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n426), .A2(G270), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n428), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n473), .B1(new_n481), .B2(G200), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n292), .B2(new_n481), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n480), .A2(new_n472), .A3(new_n318), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n484), .A2(KEYINPUT21), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT75), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(G179), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT21), .B(G169), .C1(new_n477), .C2(new_n479), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n489), .B2(new_n473), .ZN(new_n490));
  AOI211_X1 g0290(.A(KEYINPUT75), .B(new_n472), .C1(new_n487), .C2(new_n488), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n483), .B(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n431), .A2(new_n428), .A3(new_n432), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n431), .A2(G190), .A3(new_n428), .A4(new_n432), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n451), .A3(new_n461), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n390), .A2(new_n224), .A3(G68), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n224), .B1(new_n337), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(G97), .A2(G107), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n213), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n224), .A2(G33), .A3(G97), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n500), .A2(new_n502), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n266), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n302), .A2(new_n252), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n460), .A2(new_n302), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n390), .A2(G238), .A3(new_n274), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n390), .A2(G244), .A3(G1698), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n435), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n279), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n387), .A2(new_n424), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n424), .A2(new_n214), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n283), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n344), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n517), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n512), .B2(new_n279), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n509), .B(new_n518), .C1(G169), .C2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(G190), .A3(new_n517), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n456), .A2(new_n458), .A3(G87), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n523), .A2(new_n505), .A3(new_n506), .ZN(new_n524));
  INV_X1    g0324(.A(G200), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n522), .B(new_n524), .C1(new_n525), .C2(new_n520), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n428), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(G257), .B2(new_n426), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n218), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n273), .A2(new_n274), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n272), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(G1698), .C1(new_n534), .C2(new_n370), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n535), .A3(new_n464), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n390), .A2(G244), .A3(new_n274), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n531), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n530), .B1(new_n538), .B2(new_n283), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G169), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n530), .B(G179), .C1(new_n538), .C2(new_n283), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n358), .A2(KEYINPUT7), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n365), .B2(new_n269), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT7), .B1(new_n271), .B2(new_n358), .ZN(new_n545));
  OAI21_X1  g0345(.A(G107), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n219), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  AND2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n501), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n549), .B2(KEYINPUT6), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n266), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n456), .A2(new_n458), .A3(G97), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n252), .A2(G97), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n542), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n539), .A2(G200), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n558), .B(new_n555), .C1(new_n292), .C2(new_n539), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n528), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n463), .A2(new_n493), .A3(new_n497), .A4(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n411), .A2(new_n562), .ZN(G372));
  AND2_X1   g0363(.A1(new_n346), .A2(new_n320), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n349), .A2(new_n408), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n404), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n300), .B1(new_n566), .B2(new_n296), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n489), .A2(new_n473), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n485), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n463), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n497), .A3(new_n561), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT79), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n555), .B1(new_n542), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n540), .A2(KEYINPUT79), .A3(new_n541), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT26), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n527), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n555), .B1(new_n540), .B2(new_n541), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n521), .A3(new_n526), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT26), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n577), .A2(new_n521), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n571), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n567), .B1(new_n411), .B2(new_n583), .ZN(G369));
  INV_X1    g0384(.A(new_n497), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n251), .A2(new_n224), .A3(G13), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n586), .A2(KEYINPUT27), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(KEYINPUT27), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(G213), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G343), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n462), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n585), .B1(KEYINPUT80), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(KEYINPUT80), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n463), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n463), .A2(new_n591), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n485), .B1(new_n490), .B2(new_n491), .ZN(new_n600));
  INV_X1    g0400(.A(new_n591), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n597), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n569), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n472), .A2(new_n601), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n492), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G330), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n598), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n605), .A2(new_n612), .ZN(G399));
  INV_X1    g0413(.A(new_n208), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(G41), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n502), .A2(G116), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(G1), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n228), .B2(new_n616), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT28), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n591), .B1(new_n571), .B2(new_n581), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT29), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n560), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n557), .A2(KEYINPUT86), .A3(new_n559), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n497), .A2(new_n626), .A3(new_n526), .A4(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n600), .B1(new_n434), .B2(new_n462), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n579), .A2(new_n576), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT85), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n579), .A2(new_n633), .A3(new_n576), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n527), .A2(new_n573), .A3(KEYINPUT26), .A4(new_n574), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n521), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n601), .B1(new_n630), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT87), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n640), .B(new_n601), .C1(new_n630), .C2(new_n637), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n624), .B1(new_n642), .B2(new_n623), .ZN(new_n643));
  XOR2_X1   g0443(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n644));
  INV_X1    g0444(.A(KEYINPUT30), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(KEYINPUT82), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n487), .A2(new_n539), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n427), .A2(new_n647), .A3(new_n520), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n645), .A2(KEYINPUT82), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n648), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n513), .A2(new_n517), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n344), .A2(new_n481), .A3(new_n539), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n494), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n591), .B(new_n644), .C1(new_n651), .C2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n654), .B(KEYINPUT83), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n648), .B(new_n649), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n601), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n659), .B2(KEYINPUT31), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n562), .A2(new_n591), .ZN(new_n661));
  OAI21_X1  g0461(.A(G330), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT84), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT84), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n664), .B(G330), .C1(new_n660), .C2(new_n661), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n643), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n620), .B1(new_n669), .B2(G1), .ZN(G364));
  INV_X1    g0470(.A(new_n610), .ZN(new_n671));
  INV_X1    g0471(.A(G13), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G20), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n251), .B1(new_n673), .B2(G45), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n615), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(G330), .B2(new_n609), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n676), .B(KEYINPUT88), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n273), .A2(new_n208), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT89), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G355), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(G116), .B2(new_n208), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n249), .A2(G45), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n390), .A2(new_n614), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n423), .B2(new_n229), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(G13), .A2(G33), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G20), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n223), .B1(G20), .B2(new_n318), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n679), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n224), .A2(new_n344), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(G190), .A3(new_n525), .ZN(new_n697));
  INV_X1    g0497(.A(G322), .ZN(new_n698));
  NOR2_X1   g0498(.A1(G190), .A2(G200), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G311), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n697), .A2(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n224), .A2(G179), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n699), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n273), .B(new_n702), .C1(G329), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n696), .A2(G200), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G190), .ZN(new_n708));
  INV_X1    g0508(.A(G317), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT33), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n709), .A2(KEYINPUT33), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n292), .A2(G179), .A3(G200), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n224), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n703), .A2(G190), .A3(G200), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n715), .A2(G294), .B1(new_n717), .B2(G303), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n707), .A2(new_n292), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n703), .A2(new_n292), .A3(G200), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n719), .A2(G326), .B1(new_n721), .B2(G283), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n706), .A2(new_n712), .A3(new_n718), .A4(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n717), .A2(G87), .ZN(new_n725));
  INV_X1    g0525(.A(new_n719), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n201), .ZN(new_n727));
  INV_X1    g0527(.A(new_n708), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n203), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n273), .B1(new_n700), .B2(new_n217), .C1(new_n202), .C2(new_n697), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n720), .A2(new_n219), .ZN(new_n731));
  NOR4_X1   g0531(.A1(new_n727), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G159), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n704), .A2(KEYINPUT32), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT32), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n705), .B2(G159), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n734), .B(new_n736), .C1(G97), .C2(new_n715), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n723), .A2(new_n724), .B1(new_n732), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n724), .B2(new_n723), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n695), .B1(new_n739), .B2(new_n692), .ZN(new_n740));
  INV_X1    g0540(.A(new_n691), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n609), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n678), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(G396));
  NAND2_X1  g0544(.A1(new_n308), .A2(new_n591), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n317), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n320), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n320), .A2(new_n591), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n622), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n749), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n621), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n676), .B1(new_n667), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n667), .B2(new_n753), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n728), .A2(new_n756), .B1(new_n716), .B2(new_n219), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G97), .A2(new_n715), .B1(new_n719), .B2(G303), .ZN(new_n758));
  INV_X1    g0558(.A(new_n700), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n273), .B1(new_n759), .B2(G116), .ZN(new_n760));
  INV_X1    g0560(.A(new_n697), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n761), .A2(G294), .B1(new_n705), .B2(G311), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n758), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n757), .B(new_n763), .C1(G87), .C2(new_n721), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT91), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n721), .A2(G68), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n766), .B1(new_n201), .B2(new_n716), .C1(new_n202), .C2(new_n714), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n372), .B(new_n767), .C1(G132), .C2(new_n705), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT92), .B(G143), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n761), .A2(new_n769), .B1(new_n759), .B2(G159), .ZN(new_n770));
  INV_X1    g0570(.A(G137), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n770), .B1(new_n728), .B2(new_n261), .C1(new_n771), .C2(new_n726), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT34), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n773), .B2(new_n772), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n692), .B1(new_n765), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n679), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n692), .A2(new_n689), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n217), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n777), .B(new_n780), .C1(new_n751), .C2(new_n690), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n755), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G384));
  AND2_X1   g0583(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n784), .A2(new_n785), .A3(new_n469), .A4(new_n226), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT36), .ZN(new_n787));
  INV_X1    g0587(.A(new_n228), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n788), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n201), .A2(G68), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n251), .B(G13), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT98), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n375), .A2(new_n385), .ZN(new_n794));
  INV_X1    g0594(.A(new_n589), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(KEYINPUT94), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT94), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n384), .B1(new_n364), .B2(new_n374), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n589), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n404), .B2(new_n408), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT37), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n402), .A2(new_n396), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n407), .B(new_n802), .C1(new_n803), .C2(new_n798), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n799), .B2(new_n796), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n375), .A2(new_n406), .A3(new_n385), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT96), .B1(new_n806), .B2(new_n403), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT96), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n407), .B(new_n808), .C1(new_n803), .C2(new_n798), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n807), .A2(new_n800), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(KEYINPUT37), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT97), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n810), .A2(KEYINPUT97), .A3(KEYINPUT37), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n801), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n793), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n816), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n810), .A2(KEYINPUT97), .A3(KEYINPUT37), .ZN(new_n819));
  AOI21_X1  g0619(.A(KEYINPUT97), .B1(new_n810), .B2(KEYINPUT37), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n819), .A2(new_n820), .A3(new_n805), .ZN(new_n821));
  OAI211_X1 g0621(.A(KEYINPUT98), .B(new_n818), .C1(new_n821), .C2(new_n801), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n352), .B1(new_n368), .B2(new_n373), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n363), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n824), .A2(new_n255), .A3(new_n374), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n385), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n795), .ZN(new_n827));
  INV_X1    g0627(.A(new_n826), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n827), .B(new_n407), .C1(new_n828), .C2(new_n803), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n805), .B1(KEYINPUT37), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n827), .B1(new_n404), .B2(new_n408), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT38), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n817), .A2(new_n822), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT99), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n817), .A2(new_n822), .A3(KEYINPUT99), .A4(new_n833), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n332), .A2(new_n601), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n350), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n346), .B(new_n349), .C1(new_n332), .C2(new_n601), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n749), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT83), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n654), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n591), .B1(new_n843), .B2(new_n651), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT31), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n844), .B(new_n644), .C1(new_n562), .C2(new_n591), .ZN(new_n846));
  AND4_X1   g0646(.A1(KEYINPUT40), .A2(new_n841), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n836), .A2(new_n837), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT100), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n836), .A2(new_n850), .A3(new_n837), .A4(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n832), .B(KEYINPUT38), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n853), .A2(new_n841), .A3(new_n845), .A4(new_n846), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n845), .A2(new_n410), .A3(new_n846), .ZN(new_n858));
  OAI21_X1  g0658(.A(G330), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n858), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n813), .A2(new_n814), .ZN(new_n864));
  INV_X1    g0664(.A(new_n801), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n816), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n866), .A2(KEYINPUT98), .B1(KEYINPUT38), .B2(new_n832), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT39), .B1(new_n867), .B2(new_n817), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n343), .A2(new_n345), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n333), .A3(new_n601), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n404), .A2(new_n795), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n748), .B(KEYINPUT93), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n621), .B2(new_n751), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n839), .A2(new_n840), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n876), .B1(new_n881), .B2(new_n853), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n410), .B(new_n624), .C1(new_n642), .C2(new_n623), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n567), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n883), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n863), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT103), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n863), .A2(new_n886), .ZN(new_n889));
  OAI21_X1  g0689(.A(G1), .B1(new_n672), .B2(G20), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(KEYINPUT102), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT102), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n792), .B1(new_n892), .B2(new_n893), .ZN(G367));
  INV_X1    g0694(.A(new_n603), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n626), .B(new_n627), .C1(new_n555), .C2(new_n601), .ZN(new_n896));
  INV_X1    g0696(.A(new_n575), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n601), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n899), .A2(KEYINPUT42), .B1(new_n578), .B2(new_n601), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n597), .A2(KEYINPUT42), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n604), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n524), .A2(new_n601), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n527), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n521), .A2(new_n904), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT43), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n900), .A2(new_n909), .A3(new_n908), .A4(new_n902), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n611), .A2(new_n898), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n914), .B(new_n915), .Z(new_n916));
  XNOR2_X1  g0716(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n615), .B(new_n917), .Z(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n605), .A2(KEYINPUT45), .A3(new_n898), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT45), .B1(new_n605), .B2(new_n898), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT105), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(KEYINPUT44), .C1(new_n605), .C2(new_n898), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT44), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n898), .B1(KEYINPUT105), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n604), .B(new_n926), .C1(KEYINPUT105), .C2(new_n925), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n922), .A2(new_n928), .A3(new_n611), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n611), .B1(new_n922), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT106), .B1(new_n599), .B2(new_n602), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n671), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(new_n671), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(new_n895), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n929), .A2(new_n930), .A3(new_n669), .A4(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n919), .B1(new_n937), .B2(new_n669), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n916), .B1(new_n938), .B2(new_n675), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n693), .B1(new_n208), .B2(new_n303), .C1(new_n686), .C2(new_n240), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n679), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n728), .A2(new_n733), .B1(new_n716), .B2(new_n202), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G68), .B2(new_n715), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n697), .A2(new_n261), .B1(new_n704), .B2(new_n771), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n445), .B(new_n944), .C1(G50), .C2(new_n759), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n720), .A2(new_n217), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n719), .B2(new_n769), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n700), .A2(new_n756), .B1(new_n704), .B2(new_n709), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n372), .B1(new_n726), .B2(new_n701), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(G303), .C2(new_n761), .ZN(new_n951));
  INV_X1    g0751(.A(G294), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n728), .A2(new_n952), .B1(new_n219), .B2(new_n714), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G97), .B2(new_n721), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n716), .A2(new_n469), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n951), .B(new_n954), .C1(KEYINPUT46), .C2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n717), .A2(KEYINPUT46), .A3(G116), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT107), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n948), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT47), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n941), .B1(new_n960), .B2(new_n692), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n741), .B2(new_n907), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n939), .A2(new_n962), .ZN(G387));
  NAND2_X1  g0763(.A1(new_n936), .A2(new_n675), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n716), .A2(new_n217), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n303), .A2(new_n714), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n733), .B2(new_n726), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n965), .B(new_n968), .C1(G97), .C2(new_n721), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n708), .A2(new_n377), .B1(new_n759), .B2(G68), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n761), .A2(G50), .B1(new_n705), .B2(G150), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n390), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n720), .A2(new_n469), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n390), .B(new_n975), .C1(G326), .C2(new_n705), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n714), .A2(new_n756), .B1(new_n716), .B2(new_n952), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n761), .A2(G317), .B1(new_n759), .B2(G303), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n728), .B2(new_n701), .C1(new_n698), .C2(new_n726), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT48), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n980), .B2(new_n979), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT49), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n692), .B1(new_n974), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n237), .A2(new_n423), .ZN(new_n987));
  INV_X1    g0787(.A(new_n617), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n987), .A2(new_n685), .B1(new_n988), .B2(new_n681), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n617), .B(new_n423), .C1(new_n203), .C2(new_n217), .ZN(new_n990));
  XNOR2_X1  g0790(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n201), .B2(new_n377), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n259), .A2(new_n991), .A3(G50), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n989), .A2(new_n995), .B1(G107), .B2(new_n208), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n778), .B1(new_n996), .B2(new_n693), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n986), .B(new_n997), .C1(new_n599), .C2(new_n741), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n936), .A2(new_n669), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n615), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n936), .A2(new_n669), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n964), .B(new_n998), .C1(new_n1000), .C2(new_n1001), .ZN(G393));
  NAND2_X1  g0802(.A1(new_n929), .A2(new_n930), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n674), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n898), .A2(new_n741), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n245), .A2(new_n685), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n693), .B1(new_n465), .B2(new_n208), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n679), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n726), .A2(new_n709), .B1(new_n701), .B2(new_n697), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT52), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n273), .B(new_n731), .C1(G294), .C2(new_n759), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G116), .A2(new_n715), .B1(new_n708), .B2(G303), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n716), .A2(new_n756), .B1(new_n704), .B2(new_n698), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT111), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G150), .A2(new_n719), .B1(new_n761), .B2(G159), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT51), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n714), .A2(new_n217), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G68), .B2(new_n717), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n759), .A2(new_n377), .B1(new_n705), .B2(new_n769), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n708), .A2(G50), .B1(new_n721), .B2(G87), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1019), .A2(new_n390), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1013), .A2(new_n1015), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1008), .B1(new_n1023), .B2(new_n692), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1004), .B1(new_n1005), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1003), .A2(new_n999), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n615), .A3(new_n937), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(G390));
  NAND3_X1  g0828(.A1(new_n639), .A2(new_n641), .A3(new_n748), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n747), .A3(new_n879), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1030), .A2(new_n873), .A3(new_n836), .A4(new_n837), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n873), .B1(new_n878), .B2(new_n880), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n868), .B2(new_n870), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n666), .A2(new_n751), .A3(new_n879), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n845), .A2(new_n846), .A3(G330), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n841), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1036), .A2(new_n410), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n884), .A2(new_n567), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n878), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n879), .B1(new_n666), .B2(new_n751), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1037), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1029), .A2(new_n747), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1036), .A2(new_n751), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1034), .B(new_n1047), .C1(new_n879), .C2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1042), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1040), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1039), .A2(new_n1050), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n615), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1039), .A2(new_n675), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n778), .B1(new_n259), .B2(new_n779), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n761), .A2(G132), .B1(new_n705), .B2(G125), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT54), .B(G143), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n445), .B1(new_n759), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n716), .A2(new_n261), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT53), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n708), .A2(G137), .B1(new_n721), .B2(G50), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G159), .A2(new_n715), .B1(new_n719), .B2(G128), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G97), .A2(new_n759), .B1(new_n705), .B2(G294), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n273), .B1(new_n761), .B2(G116), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n725), .A4(new_n766), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1018), .B1(G283), .B2(new_n719), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n219), .B2(new_n728), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1066), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT112), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT112), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n692), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1056), .B1(new_n1073), .B2(new_n1075), .C1(new_n871), .C2(new_n690), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1054), .A2(new_n1055), .A3(new_n1076), .ZN(G378));
  INV_X1    g0877(.A(KEYINPUT57), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1042), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1053), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT117), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n856), .A2(G330), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n852), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n296), .A2(new_n301), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n267), .A2(new_n795), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT114), .Z(new_n1089));
  XNOR2_X1  g0889(.A(new_n1087), .B(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(KEYINPUT115), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n883), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1091), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n852), .A2(new_n1083), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n852), .B2(new_n1083), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1082), .B(new_n1091), .C1(new_n849), .C2(new_n851), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n883), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1081), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n883), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1080), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1053), .A2(new_n1079), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1093), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n1101), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n616), .B1(new_n1106), .B2(new_n1078), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n675), .B1(new_n1105), .B2(new_n1101), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1090), .A2(new_n689), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n390), .A2(G41), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n761), .A2(G107), .B1(new_n705), .B2(G283), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n303), .B2(new_n700), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n965), .B(new_n1114), .C1(G68), .C2(new_n715), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n726), .A2(new_n469), .B1(new_n720), .B2(new_n202), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G97), .B2(new_n708), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1115), .A2(new_n1117), .A3(new_n1110), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT58), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1112), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(G33), .B(G41), .C1(new_n705), .C2(G124), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n761), .A2(G128), .B1(new_n759), .B2(G137), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n716), .B2(new_n1058), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G150), .A2(new_n715), .B1(new_n719), .B2(G125), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT113), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(G132), .C2(new_n708), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT59), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1121), .B1(new_n733), .B2(new_n720), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1120), .B1(new_n1119), .B2(new_n1118), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n692), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n675), .B(new_n615), .C1(new_n201), .C2(new_n779), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1109), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1108), .A2(KEYINPUT116), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT116), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n674), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n1133), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1103), .A2(new_n1107), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(G375));
  NAND2_X1  g0940(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n880), .A2(new_n689), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n692), .A2(G68), .A3(new_n689), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n697), .A2(new_n771), .B1(new_n700), .B2(new_n261), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G128), .B2(new_n705), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G50), .A2(new_n715), .B1(new_n719), .B2(G132), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n708), .A2(new_n1059), .B1(new_n717), .B2(G159), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n372), .B1(G58), .B2(new_n721), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n719), .A2(G294), .B1(new_n759), .B2(G107), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n469), .B2(new_n728), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT118), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n717), .A2(G97), .B1(new_n705), .B2(G303), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT119), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n273), .B(new_n946), .C1(G283), .C2(new_n761), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n967), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n778), .B(new_n1143), .C1(new_n1157), .C2(new_n692), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1141), .A2(new_n675), .B1(new_n1142), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT120), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1042), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n918), .A3(new_n1051), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT121), .Z(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(G381));
  OR2_X1    g0966(.A1(G393), .A2(G396), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(G387), .A2(G390), .A3(G384), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(G375), .A2(G378), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1165), .A3(new_n1169), .ZN(G407));
  NAND2_X1  g0970(.A1(new_n590), .A2(G213), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(G407), .A2(G213), .A3(new_n1173), .ZN(G409));
  AOI22_X1  g0974(.A1(new_n1096), .A2(new_n1099), .B1(new_n1053), .B2(new_n1079), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1133), .B1(new_n1175), .B2(new_n918), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n675), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G378), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1139), .B2(G378), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT124), .B1(new_n1179), .B2(new_n1172), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT60), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1162), .B1(new_n1181), .B2(new_n1050), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1161), .A2(KEYINPUT60), .A3(new_n1042), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n615), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1160), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(G384), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1107), .A2(new_n1103), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(G378), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1190));
  INV_X1    g0990(.A(G378), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n1171), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1180), .A2(new_n1186), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT62), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT61), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1193), .A2(new_n1186), .A3(new_n1171), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT122), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT62), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1193), .A2(new_n1186), .A3(KEYINPUT122), .A4(new_n1171), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1172), .A2(G2897), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1186), .B(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1194), .B1(new_n1193), .B2(new_n1171), .ZN(new_n1207));
  AOI211_X1 g1007(.A(KEYINPUT124), .B(new_n1172), .C1(new_n1189), .C2(new_n1192), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1197), .A2(new_n1198), .A3(new_n1204), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1209), .A2(new_n1198), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1213), .A2(new_n1197), .A3(KEYINPUT125), .A4(new_n1204), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(G387), .A2(new_n1027), .A3(new_n1025), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(G393), .B(new_n743), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G390), .A2(new_n939), .A3(new_n962), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT126), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1216), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT126), .B1(new_n1225), .B2(new_n1218), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1212), .A2(new_n1214), .A3(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1206), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1229));
  AND4_X1   g1029(.A1(new_n1198), .A2(new_n1229), .A3(new_n1225), .A4(new_n1218), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1232));
  XOR2_X1   g1032(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1233));
  OAI221_X1 g1033(.A(new_n1230), .B1(new_n1231), .B2(new_n1196), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(new_n1234), .ZN(G405));
  OAI21_X1  g1035(.A(KEYINPUT127), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1220), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT127), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1225), .A2(new_n1218), .A3(KEYINPUT126), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1139), .B(G378), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(new_n1186), .Z(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1236), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(KEYINPUT127), .B(new_n1242), .C1(new_n1222), .C2(new_n1226), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(G402));
endmodule


