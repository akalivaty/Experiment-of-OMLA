//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XOR2_X1   g000(.A(KEYINPUT93), .B(G36gat), .Z(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  OR3_X1    g002(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n204));
  AOI22_X1  g003(.A1(new_n202), .A2(G29gat), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G43gat), .B(G50gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT94), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n206), .A2(new_n207), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT17), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(KEYINPUT8), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT100), .ZN(new_n217));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT7), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G99gat), .B(G106gat), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n221), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n217), .A2(new_n223), .A3(new_n219), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n213), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n222), .A2(new_n224), .ZN(new_n227));
  INV_X1    g026(.A(new_n211), .ZN(new_n228));
  AND2_X1   g027(.A1(G232gat), .A2(G233gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n227), .A2(new_n228), .B1(KEYINPUT41), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G190gat), .B(G218gat), .Z(new_n232));
  AND2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n229), .A2(KEYINPUT41), .ZN(new_n235));
  XNOR2_X1  g034(.A(G134gat), .B(G162gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OR3_X1    g037(.A1(new_n233), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n233), .B2(new_n234), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(G15gat), .B(G22gat), .Z(new_n242));
  INV_X1    g041(.A(G1gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT96), .ZN(new_n245));
  XNOR2_X1  g044(.A(G15gat), .B(G22gat), .ZN(new_n246));
  OR3_X1    g045(.A1(new_n246), .A2(KEYINPUT96), .A3(G1gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n243), .A2(KEYINPUT95), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT95), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT16), .B1(new_n249), .B2(G1gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G8gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT97), .ZN(new_n254));
  INV_X1    g053(.A(G8gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n244), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(G71gat), .A2(G78gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(G71gat), .A2(G78gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G57gat), .B(G64gat), .Z(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(KEYINPUT98), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(KEYINPUT9), .B2(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI221_X1 g062(.A(new_n260), .B1(KEYINPUT9), .B2(new_n257), .C1(new_n259), .C2(KEYINPUT98), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT99), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(KEYINPUT99), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT21), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n254), .B(new_n256), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n271), .ZN(new_n274));
  INV_X1    g073(.A(G231gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n274), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G127gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n279), .A2(new_n280), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n273), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n283), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n281), .A3(new_n272), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G155gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G183gat), .B(G211gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n284), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n290), .B1(new_n284), .B2(new_n286), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n241), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT101), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT101), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n241), .C1(new_n291), .C2(new_n292), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT102), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n269), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n269), .A2(new_n225), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n222), .A2(new_n264), .A3(new_n263), .A4(new_n224), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n300), .B(new_n301), .C1(new_n304), .C2(KEYINPUT10), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT10), .B1(new_n302), .B2(new_n303), .ZN(new_n306));
  INV_X1    g105(.A(new_n301), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT102), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G230gat), .A2(G233gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n309), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n302), .A2(KEYINPUT103), .A3(new_n311), .A4(new_n303), .ZN(new_n312));
  XNOR2_X1  g111(.A(G120gat), .B(G148gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT103), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n304), .A2(new_n311), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT105), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n307), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n309), .B(KEYINPUT104), .Z(new_n323));
  OAI21_X1  g122(.A(new_n318), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n315), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n320), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n321), .B1(new_n320), .B2(new_n326), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n299), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n213), .A2(new_n254), .A3(new_n256), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n254), .A2(new_n256), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n228), .ZN(new_n334));
  NAND2_X1  g133(.A1(G229gat), .A2(G233gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT18), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT18), .A4(new_n335), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n254), .A2(new_n211), .A3(new_n256), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n335), .B(KEYINPUT13), .Z(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n338), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G197gat), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT11), .B(G169gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n348), .B(KEYINPUT12), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n338), .A2(new_n351), .A3(new_n339), .A4(new_n343), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  INV_X1    g154(.A(G169gat), .ZN(new_n356));
  INV_X1    g155(.A(G176gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT23), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT24), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT24), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n360), .B(new_n362), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n355), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n360), .A2(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n367), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT67), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n363), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n362), .A2(KEYINPUT25), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n359), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT66), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n373), .A2(new_n378), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT68), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT27), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(G183gat), .ZN(new_n387));
  INV_X1    g186(.A(G183gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(KEYINPUT27), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n385), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(KEYINPUT27), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(G183gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT68), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT28), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(G190gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT69), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT69), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n390), .A2(new_n398), .A3(new_n393), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n391), .A2(new_n392), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n394), .B1(new_n400), .B2(G190gat), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n356), .B(new_n357), .C1(KEYINPUT71), .C2(KEYINPUT26), .ZN(new_n403));
  AND2_X1   g202(.A1(KEYINPUT71), .A2(KEYINPUT26), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n359), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT70), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT70), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n408), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n364), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT72), .B(new_n364), .C1(new_n405), .C2(new_n410), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n384), .B1(new_n402), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT1), .ZN(new_n417));
  INV_X1    g216(.A(G120gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n419));
  INV_X1    g218(.A(G134gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G127gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n280), .A2(G134gat), .ZN(new_n422));
  AND4_X1   g221(.A1(new_n417), .A2(new_n419), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(G113gat), .ZN(new_n424));
  INV_X1    g223(.A(G113gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G120gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT73), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n426), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(new_n422), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n423), .A2(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n428), .A2(new_n417), .A3(new_n434), .A4(new_n419), .ZN(new_n435));
  XNOR2_X1  g234(.A(G113gat), .B(G120gat), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n436), .B2(KEYINPUT1), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n384), .B(new_n438), .C1(new_n402), .C2(new_n415), .ZN(new_n439));
  NAND2_X1  g238(.A1(G227gat), .A2(G233gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n440), .B(KEYINPUT64), .Z(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT32), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(G15gat), .B(G43gat), .Z(new_n446));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n443), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n448), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n442), .B(KEYINPUT32), .C1(new_n444), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n439), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n440), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n441), .A2(KEYINPUT34), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n454), .A2(KEYINPUT34), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n449), .A2(new_n456), .A3(new_n451), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(G228gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G155gat), .A2(G162gat), .ZN(new_n463));
  INV_X1    g262(.A(G155gat), .ZN(new_n464));
  INV_X1    g263(.A(G162gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G141gat), .B(G148gat), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n463), .B(new_n466), .C1(new_n467), .C2(KEYINPUT2), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT3), .ZN(new_n469));
  INV_X1    g268(.A(G141gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G148gat), .ZN(new_n471));
  INV_X1    g270(.A(G148gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G141gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G155gat), .B(G162gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n463), .A2(KEYINPUT2), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n468), .A2(new_n469), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT29), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT22), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT74), .B(G218gat), .ZN(new_n482));
  INV_X1    g281(.A(G211gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G197gat), .B(G204gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G211gat), .B(G218gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n485), .ZN(new_n488));
  INV_X1    g287(.A(new_n486), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n480), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n474), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n487), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n486), .B1(new_n484), .B2(new_n485), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n479), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT82), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT3), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT29), .B1(new_n490), .B2(new_n487), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT82), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n494), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n491), .B1(new_n502), .B2(KEYINPUT83), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n468), .A2(new_n477), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n469), .B1(new_n500), .B2(KEYINPUT82), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n497), .A2(new_n498), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n462), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n468), .A2(KEYINPUT78), .A3(new_n477), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT78), .B1(new_n468), .B2(new_n477), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n500), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT78), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n492), .B2(new_n493), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n468), .A2(KEYINPUT78), .A3(new_n477), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n469), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n462), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n490), .A2(new_n487), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT75), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n480), .B(KEYINPUT84), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G78gat), .B(G106gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT31), .B(G50gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT85), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n510), .A2(new_n524), .A3(new_n528), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(G22gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n502), .A2(KEYINPUT83), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n507), .A2(new_n508), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n491), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n523), .B1(new_n536), .B2(new_n462), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n533), .B1(new_n537), .B2(new_n528), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n530), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(G22gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n533), .A3(new_n528), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n537), .A2(new_n528), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(KEYINPUT85), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n460), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G1gat), .B(G29gat), .Z(new_n545));
  XNOR2_X1  g344(.A(G57gat), .B(G85gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G225gat), .A2(G233gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n432), .B1(new_n515), .B2(new_n516), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n438), .A2(new_n504), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n478), .A2(new_n438), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n551), .B1(new_n517), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT4), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n494), .A2(new_n432), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT4), .B1(new_n438), .B2(new_n504), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(KEYINPUT5), .B(new_n555), .C1(new_n557), .C2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT3), .B1(new_n511), .B2(new_n512), .ZN(new_n563));
  INV_X1    g362(.A(new_n556), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT80), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n567), .B(KEYINPUT4), .C1(new_n438), .C2(new_n504), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n552), .A2(KEYINPUT5), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n550), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT6), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT81), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT6), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n570), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(new_n549), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(new_n571), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n416), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G226gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(new_n276), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n384), .B(KEYINPUT76), .C1(new_n402), .C2(new_n415), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(KEYINPUT29), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n416), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n521), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n589), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n584), .B2(new_n587), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n416), .A2(new_n585), .A3(new_n276), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n520), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n588), .A2(KEYINPUT77), .A3(new_n521), .A4(new_n590), .ZN(new_n598));
  XNOR2_X1  g397(.A(G8gat), .B(G36gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G64gat), .B(G92gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  NAND4_X1  g400(.A1(new_n593), .A2(new_n597), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT30), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n597), .A2(new_n598), .ZN(new_n605));
  INV_X1    g404(.A(new_n601), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(new_n603), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n593), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n606), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n582), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n544), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT35), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT86), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n604), .A2(new_n608), .A3(new_n610), .A4(KEYINPUT86), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT89), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n562), .A2(new_n619), .A3(new_n570), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n562), .B2(new_n570), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n620), .A2(new_n621), .A3(new_n550), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n575), .B(new_n574), .C1(new_n622), .C2(new_n579), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n624));
  NAND4_X1  g423(.A1(new_n623), .A2(new_n459), .A3(new_n458), .A4(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n539), .B2(new_n543), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT92), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n618), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n618), .B2(new_n626), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n614), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n552), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT87), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(KEYINPUT87), .A3(new_n552), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n553), .A2(new_n554), .A3(new_n552), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n634), .A2(KEYINPUT39), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(KEYINPUT88), .A3(new_n550), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT88), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT39), .B1(new_n634), .B2(new_n635), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n549), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n638), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n622), .B1(new_n646), .B2(KEYINPUT40), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT88), .B1(new_n641), .B2(new_n550), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n644), .A2(new_n643), .A3(new_n549), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n637), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n616), .A2(new_n647), .A3(new_n617), .A4(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n595), .A2(new_n520), .A3(new_n596), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n521), .B1(new_n588), .B2(new_n590), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT37), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT90), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n601), .B1(new_n605), .B2(new_n593), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT37), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n601), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n659), .B(new_n660), .C1(new_n661), .C2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n609), .B2(new_n606), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n605), .B2(new_n593), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT38), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT90), .B1(new_n665), .B2(new_n658), .ZN(new_n668));
  INV_X1    g467(.A(new_n602), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n623), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n664), .A2(new_n667), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n539), .A2(new_n543), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n653), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n581), .A2(new_n604), .A3(new_n610), .A4(new_n608), .ZN(new_n675));
  INV_X1    g474(.A(new_n460), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT36), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT36), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n460), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n674), .A2(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n354), .B1(new_n630), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n331), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n581), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n243), .ZN(G1324gat));
  INV_X1    g484(.A(new_n618), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n687), .A2(KEYINPUT106), .A3(new_n330), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT106), .B1(new_n687), .B2(new_n330), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(G8gat), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n330), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(KEYINPUT42), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n692), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n688), .B2(new_n689), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n690), .B(new_n693), .C1(new_n695), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g495(.A(new_n683), .ZN(new_n697));
  AOI21_X1  g496(.A(G15gat), .B1(new_n697), .B2(new_n676), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n677), .A2(new_n679), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT107), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n698), .B1(new_n697), .B2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n683), .A2(new_n672), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  AOI21_X1  g505(.A(new_n241), .B1(new_n630), .B2(new_n681), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n291), .A2(new_n292), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n329), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n354), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(G29gat), .A3(new_n581), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT45), .Z(new_n713));
  NOR2_X1   g512(.A1(new_n241), .A2(KEYINPUT44), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(new_n612), .B2(new_n672), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n674), .A2(new_n717), .A3(new_n675), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n673), .A2(new_n699), .A3(new_n716), .A4(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n715), .B1(new_n630), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n241), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT35), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n544), .B2(new_n612), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n618), .A2(new_n626), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT92), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n618), .A2(new_n626), .A3(new_n627), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n673), .A2(new_n680), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n721), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n720), .B1(new_n729), .B2(KEYINPUT44), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n710), .ZN(new_n732));
  OAI21_X1  g531(.A(G29gat), .B1(new_n732), .B2(new_n581), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n733), .ZN(G1328gat));
  OAI21_X1  g533(.A(new_n202), .B1(new_n732), .B2(new_n618), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n687), .A2(new_n202), .A3(new_n241), .A4(new_n709), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(KEYINPUT109), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n735), .B(new_n738), .C1(new_n736), .C2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n460), .A2(G43gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n711), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n731), .A2(new_n700), .A3(new_n710), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(G43gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1330gat));
  NOR3_X1   g548(.A1(new_n711), .A2(G50gat), .A3(new_n672), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n731), .A2(new_n674), .A3(new_n710), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G50gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n752), .B(new_n753), .Z(G1331gat));
  NAND2_X1  g553(.A1(new_n630), .A2(new_n719), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n295), .A2(new_n298), .A3(new_n353), .A4(new_n329), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n582), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g559(.A1(new_n757), .A2(new_n618), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(G1333gat));
  NAND3_X1  g564(.A1(new_n758), .A2(G71gat), .A3(new_n700), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n757), .A2(new_n460), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n768));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n767), .B2(KEYINPUT112), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n766), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n758), .A2(new_n674), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n708), .A2(new_n354), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n329), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT113), .B1(new_n730), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n707), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n779), .B(new_n776), .C1(new_n781), .C2(new_n720), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n582), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G85gat), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n775), .A2(new_n241), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n755), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n329), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n581), .A2(G85gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT114), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n784), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1336gat));
  NAND2_X1  g595(.A1(new_n787), .A2(new_n788), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n618), .A2(G92gat), .A3(new_n329), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(G92gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n730), .A2(new_n618), .A3(new_n777), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n778), .A2(new_n686), .A3(new_n782), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n798), .B(KEYINPUT115), .Z(new_n804));
  AOI22_X1  g603(.A1(new_n803), .A2(G92gat), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(G1337gat));
  NAND3_X1  g606(.A1(new_n778), .A2(new_n700), .A3(new_n782), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G99gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n789), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n460), .A2(G99gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(G1338gat));
  NOR2_X1   g611(.A1(new_n672), .A2(G106gat), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n789), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n674), .B(new_n776), .C1(new_n781), .C2(new_n720), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n778), .A2(new_n674), .A3(new_n782), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n821), .A2(G106gat), .B1(new_n789), .B2(new_n813), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n341), .A2(new_n342), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n335), .B1(new_n332), .B2(new_n334), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n348), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n352), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n327), .B2(new_n328), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n322), .B2(new_n323), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n310), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n323), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n831), .B(new_n834), .C1(new_n306), .C2(new_n307), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT117), .A3(new_n325), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT117), .B1(new_n835), .B2(new_n325), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n839), .A2(new_n840), .B1(new_n350), .B2(new_n352), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n835), .A2(new_n325), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n844), .A2(new_n836), .B1(new_n310), .B2(new_n832), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(KEYINPUT55), .B1(new_n310), .B2(new_n319), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n825), .A2(new_n830), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n829), .B(KEYINPUT118), .C1(new_n327), .C2(new_n328), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n721), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n839), .A2(new_n840), .ZN(new_n850));
  AND4_X1   g649(.A1(new_n721), .A2(new_n846), .A3(new_n829), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n708), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n294), .A2(new_n329), .A3(new_n354), .A4(new_n297), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n674), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n854), .A2(new_n582), .A3(new_n618), .A4(new_n676), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n354), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(new_n425), .ZN(G1340gat));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n329), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(new_n418), .ZN(G1341gat));
  NOR2_X1   g658(.A1(new_n855), .A2(new_n708), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(new_n280), .ZN(G1342gat));
  NOR4_X1   g660(.A1(new_n241), .A2(new_n460), .A3(new_n581), .A4(G134gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n618), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT119), .Z(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n855), .B2(new_n241), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n865), .B(new_n866), .C1(KEYINPUT56), .C2(new_n863), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n830), .A2(new_n825), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n845), .A2(KEYINPUT55), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(new_n850), .A3(new_n353), .A4(new_n320), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n848), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n851), .B1(new_n872), .B2(new_n241), .ZN(new_n873));
  INV_X1    g672(.A(new_n708), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n853), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n674), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n700), .A2(new_n686), .A3(new_n581), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n470), .A3(new_n353), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n830), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n829), .B(KEYINPUT120), .C1(new_n327), .C2(new_n328), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n871), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n851), .B1(new_n884), .B2(new_n241), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n853), .B1(new_n885), .B2(new_n874), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n674), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n875), .A2(new_n889), .A3(new_n674), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n888), .A2(new_n353), .A3(new_n890), .A4(new_n877), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT122), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n891), .A2(KEYINPUT122), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n868), .B(new_n880), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n891), .A2(G141gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n880), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT121), .B1(new_n897), .B2(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n899), .B(new_n868), .C1(new_n896), .C2(new_n880), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n895), .B1(new_n898), .B2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(new_n329), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n879), .A2(new_n472), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n878), .B1(new_n887), .B2(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n890), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(new_n329), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(KEYINPUT59), .A3(new_n472), .ZN(new_n907));
  XNOR2_X1  g706(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n886), .A2(new_n889), .A3(new_n674), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n672), .B1(new_n852), .B2(new_n853), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n889), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n911), .A2(new_n329), .A3(new_n878), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n908), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n903), .B1(new_n907), .B2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n905), .B2(new_n708), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n879), .A2(new_n464), .A3(new_n874), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n905), .B2(new_n241), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n879), .A2(new_n465), .A3(new_n721), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n686), .A2(new_n581), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n875), .A2(new_n544), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n353), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(new_n356), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT125), .ZN(G1348gat));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n902), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n390), .A2(new_n393), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n925), .A2(new_n874), .ZN(new_n932));
  MUX2_X1   g731(.A(new_n931), .B(new_n388), .S(new_n932), .Z(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n933), .B(new_n934), .ZN(G1350gat));
  NOR2_X1   g734(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n925), .B2(new_n721), .ZN(new_n937));
  NAND2_X1  g736(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n937), .B(new_n938), .Z(G1351gat));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n700), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n876), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(G197gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n353), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n886), .A2(new_n889), .A3(new_n674), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n889), .B1(new_n875), .B2(new_n674), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT126), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n909), .B(new_n948), .C1(new_n910), .C2(new_n889), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n354), .B(new_n941), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  OAI21_X1  g750(.A(G197gat), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n941), .B1(new_n947), .B2(new_n949), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(new_n951), .A3(new_n353), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n944), .B1(new_n952), .B2(new_n954), .ZN(G1352gat));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n942), .A2(new_n956), .A3(new_n902), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  AND2_X1   g757(.A1(new_n953), .A2(new_n902), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n956), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n483), .A3(new_n874), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n911), .A2(new_n708), .A3(new_n941), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n942), .B2(new_n721), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n241), .A2(new_n482), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n953), .B2(new_n967), .ZN(G1355gat));
endmodule


