//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(new_n202), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n225), .A2(new_n210), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n213), .B(new_n219), .C1(new_n220), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n220), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n227), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT76), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(G274), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G232), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT74), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT74), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G190), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G87), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT73), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT73), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G33), .A3(G87), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT70), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n262), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G223), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G226), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(G1698), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n267), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n261), .B1(new_n277), .B2(new_n252), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n260), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n264), .A2(new_n266), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n270), .A2(G33), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n262), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT70), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(G1698), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G223), .B2(G1698), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n280), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n252), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n256), .ZN(new_n290));
  AOI21_X1  g0090(.A(G200), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n247), .B1(new_n279), .B2(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n289), .A2(new_n261), .A3(new_n258), .A4(new_n259), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n273), .A2(new_n276), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n252), .B1(new_n295), .B2(new_n280), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n294), .B1(new_n296), .B2(new_n256), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(KEYINPUT76), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g0099(.A(KEYINPUT8), .B(G58), .Z(new_n300));
  NAND2_X1  g0100(.A1(new_n207), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n304), .A2(new_n217), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n302), .B2(KEYINPUT72), .ZN(new_n308));
  INV_X1    g0108(.A(new_n306), .ZN(new_n309));
  INV_X1    g0109(.A(new_n300), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n303), .A2(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(G58), .A2(G68), .ZN(new_n313));
  OAI21_X1  g0113(.A(G20), .B1(new_n313), .B2(new_n202), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G20), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G159), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n271), .A2(new_n272), .ZN(new_n319));
  AOI21_X1  g0119(.A(G20), .B1(new_n319), .B2(new_n281), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT7), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT7), .B1(new_n273), .B2(G20), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n305), .B1(new_n324), .B2(KEYINPUT16), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT16), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT71), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n270), .B2(G33), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n262), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n281), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n321), .B1(new_n330), .B2(new_n208), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n332));
  AOI211_X1 g0132(.A(KEYINPUT7), .B(G20), .C1(new_n281), .C2(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n331), .A2(new_n318), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n326), .B1(new_n334), .B2(new_n317), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n312), .B1(new_n325), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n299), .A2(new_n336), .A3(KEYINPUT17), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT17), .B1(new_n299), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n256), .B1(new_n287), .B2(new_n288), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n277), .B2(new_n252), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n340), .A2(G169), .B1(new_n260), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n304), .A2(new_n217), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n284), .A2(new_n321), .A3(new_n208), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(new_n323), .A3(G68), .ZN(new_n346));
  INV_X1    g0146(.A(new_n317), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n335), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n349), .B2(new_n311), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI211_X1 g0152(.A(KEYINPUT18), .B(new_n343), .C1(new_n349), .C2(new_n311), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT75), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT75), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT18), .B1(new_n336), .B2(new_n343), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n350), .A2(new_n351), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n339), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n281), .A2(new_n332), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G222), .A2(G1698), .ZN(new_n362));
  INV_X1    g0162(.A(G1698), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G223), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n288), .C1(G77), .C2(new_n361), .ZN(new_n366));
  INV_X1    g0166(.A(new_n253), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n252), .A2(new_n254), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(G226), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n370), .A3(G190), .ZN(new_n371));
  XOR2_X1   g0171(.A(new_n371), .B(KEYINPUT68), .Z(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n301), .A2(G50), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n307), .A2(new_n374), .B1(G50), .B2(new_n306), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n262), .A2(G20), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n300), .A2(new_n376), .B1(G150), .B2(new_n315), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n203), .A2(G20), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n375), .B1(new_n379), .B2(new_n344), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(KEYINPUT9), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n366), .A2(new_n370), .ZN(new_n382));
  AOI22_X1  g0182(.A1(G200), .A2(new_n382), .B1(new_n380), .B2(KEYINPUT9), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n372), .A2(new_n373), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n371), .B(KEYINPUT68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n381), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT10), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G169), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n380), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G179), .B2(new_n382), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n300), .A2(new_n315), .B1(G20), .B2(G77), .ZN(new_n393));
  INV_X1    g0193(.A(new_n376), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT15), .B(G87), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G77), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n396), .A2(new_n344), .B1(new_n397), .B2(new_n309), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT67), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n305), .A2(new_n399), .A3(new_n306), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT67), .B1(new_n309), .B2(new_n344), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(G77), .A3(new_n301), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G244), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n253), .B1(new_n405), .B2(new_n368), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n361), .A2(G238), .A3(G1698), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n361), .A2(G232), .A3(new_n363), .ZN(new_n408));
  INV_X1    g0208(.A(G107), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(new_n361), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n406), .B1(new_n410), .B2(new_n288), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G190), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n404), .B(new_n412), .C1(new_n294), .C2(new_n411), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n341), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n398), .A2(new_n403), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(G169), .C2(new_n411), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n315), .A2(G50), .B1(G20), .B2(new_n318), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n394), .B2(new_n397), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(new_n344), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(KEYINPUT11), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n402), .A2(G68), .A3(new_n301), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n309), .A2(new_n318), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT12), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(KEYINPUT11), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G238), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n253), .B1(new_n427), .B2(new_n368), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n275), .A2(new_n363), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n232), .A2(G1698), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n281), .A2(new_n429), .A3(new_n332), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n252), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n435), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n428), .B2(new_n433), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n389), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n436), .B(G179), .C1(new_n442), .C2(new_n434), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n439), .B2(new_n440), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n426), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n294), .B1(new_n436), .B2(new_n438), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n434), .A2(new_n442), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n435), .B2(new_n434), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n448), .B2(G190), .ZN(new_n449));
  INV_X1    g0249(.A(new_n426), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n417), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n359), .A2(new_n392), .A3(new_n452), .ZN(new_n453));
  MUX2_X1   g0253(.A(G257), .B(G264), .S(G1698), .Z(new_n454));
  NAND2_X1  g0254(.A1(new_n273), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n360), .A2(G303), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n252), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n207), .B(G45), .C1(new_n248), .C2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G41), .ZN(new_n460));
  OAI211_X1 g0260(.A(G270), .B(new_n252), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n252), .A2(G274), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT78), .B1(new_n459), .B2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT78), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n248), .A3(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n459), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n249), .A2(G1), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n463), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n461), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(G169), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n207), .A2(new_n471), .A3(G13), .A4(G20), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT81), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n304), .A2(new_n217), .B1(G20), .B2(new_n471), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n208), .C1(G33), .C2(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n474), .A2(KEYINPUT20), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT20), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n471), .B1(new_n207), .B2(G33), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n400), .A2(new_n401), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT82), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n479), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n474), .A2(KEYINPUT20), .A3(new_n477), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n400), .A2(new_n401), .A3(new_n481), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n473), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n470), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n483), .A2(new_n489), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n468), .A2(new_n462), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n273), .A2(new_n454), .B1(G303), .B2(new_n360), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n461), .C1(new_n493), .C2(new_n252), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n341), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n490), .A2(KEYINPUT21), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(G200), .ZN(new_n498));
  INV_X1    g0298(.A(new_n457), .ZN(new_n499));
  INV_X1    g0299(.A(new_n469), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(G190), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n470), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n491), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n496), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT83), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT83), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n496), .A2(new_n502), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n273), .A2(new_n208), .A3(G68), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT19), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n376), .A2(new_n513), .A3(G97), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n263), .B1(new_n432), .B2(new_n208), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(new_n513), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n344), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n395), .A2(new_n309), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n207), .A2(G33), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n306), .A2(new_n521), .A3(new_n217), .A4(new_n304), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n395), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(KEYINPUT79), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n522), .B2(new_n395), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n519), .A2(new_n520), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  INV_X1    g0330(.A(G274), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n467), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n252), .C1(G250), .C2(new_n467), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G238), .A2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n405), .B2(G1698), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n273), .A2(new_n535), .B1(G33), .B2(G116), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n536), .B2(new_n252), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G169), .ZN(new_n538));
  OAI211_X1 g0338(.A(G179), .B(new_n533), .C1(new_n536), .C2(new_n252), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n529), .A2(new_n530), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n518), .A2(new_n344), .B1(new_n309), .B2(new_n395), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(KEYINPUT80), .A3(new_n528), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n405), .A2(G1698), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT4), .B1(new_n273), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n281), .A2(new_n332), .A3(G250), .A4(G1698), .ZN(new_n546));
  AND2_X1   g0346(.A1(KEYINPUT4), .A2(G244), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n281), .A2(new_n332), .A3(new_n547), .A4(new_n363), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n548), .A3(new_n475), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n288), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n252), .B1(new_n458), .B2(new_n460), .ZN(new_n551));
  INV_X1    g0351(.A(G257), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n551), .A2(new_n552), .B1(new_n468), .B2(new_n462), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(G169), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n550), .A2(new_n341), .A3(new_n554), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n331), .A2(new_n409), .A3(new_n333), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n476), .A2(KEYINPUT6), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g0362(.A(KEYINPUT77), .B(G107), .Z(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g0364(.A(KEYINPUT77), .B(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n561), .A3(new_n560), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(G20), .B1(G77), .B2(new_n315), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n305), .B1(new_n559), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n306), .A2(G97), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n522), .B2(new_n476), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n556), .B(new_n557), .C1(new_n569), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(G20), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n315), .A2(G77), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n344), .B1(new_n576), .B2(new_n558), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n550), .A2(new_n554), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  INV_X1    g0379(.A(new_n572), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n550), .A2(G190), .A3(new_n554), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n577), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n537), .A2(G200), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n523), .A2(G87), .ZN(new_n584));
  OAI211_X1 g0384(.A(G190), .B(new_n533), .C1(new_n536), .C2(new_n252), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n583), .A2(new_n541), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n543), .A2(new_n573), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n273), .A2(KEYINPUT22), .A3(new_n208), .A4(G87), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n281), .A2(new_n332), .A3(new_n208), .A4(G87), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n589), .A2(new_n590), .B1(G116), .B2(new_n376), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT84), .B1(new_n208), .B2(G107), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT23), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n588), .A2(new_n591), .A3(new_n596), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n344), .ZN(new_n599));
  OAI211_X1 g0399(.A(G264), .B(new_n252), .C1(new_n458), .C2(new_n460), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n552), .A2(G1698), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G250), .B2(G1698), .ZN(new_n603));
  INV_X1    g0403(.A(G294), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n284), .A2(new_n603), .B1(new_n262), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n601), .B1(new_n605), .B2(new_n288), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n261), .A3(new_n492), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G250), .A2(G1698), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n552), .B2(G1698), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n273), .A2(new_n609), .B1(G33), .B2(G294), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n492), .B(new_n600), .C1(new_n610), .C2(new_n252), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n294), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT25), .B1(new_n309), .B2(new_n409), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n309), .A2(KEYINPUT25), .A3(new_n409), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(G107), .B2(new_n523), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n599), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n606), .A2(G179), .A3(new_n492), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(G169), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n305), .B1(new_n595), .B2(new_n597), .ZN(new_n622));
  INV_X1    g0422(.A(new_n617), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT85), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n618), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n587), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n453), .A2(new_n511), .A3(new_n629), .ZN(G372));
  NAND3_X1  g0430(.A1(new_n496), .A2(new_n506), .A3(new_n624), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n573), .A2(new_n582), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n538), .A2(new_n539), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n529), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n586), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n631), .A2(new_n632), .A3(new_n618), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n543), .A2(new_n586), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT26), .B1(new_n637), .B2(new_n573), .ZN(new_n638));
  INV_X1    g0438(.A(new_n634), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n586), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n573), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n636), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n453), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n391), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n352), .A2(new_n353), .ZN(new_n647));
  INV_X1    g0447(.A(new_n445), .ZN(new_n648));
  INV_X1    g0448(.A(new_n416), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n451), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT17), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n293), .A2(KEYINPUT76), .A3(new_n297), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT76), .B1(new_n293), .B2(new_n297), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n349), .A2(new_n311), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n299), .A2(new_n336), .A3(KEYINPUT17), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n647), .B1(new_n650), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n646), .B1(new_n659), .B2(new_n388), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT86), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(G213), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n511), .B1(new_n497), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n496), .A2(new_n506), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n491), .A3(new_n668), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n670), .B2(new_n673), .ZN(new_n675));
  OAI21_X1  g0475(.A(G330), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n599), .A2(new_n617), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n668), .ZN(new_n678));
  INV_X1    g0478(.A(new_n628), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n627), .B1(new_n618), .B2(new_n624), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n677), .A2(new_n621), .A3(new_n668), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT88), .Z(new_n683));
  AOI21_X1  g0483(.A(new_n676), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n672), .A2(new_n669), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n683), .B2(new_n681), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n677), .A2(new_n621), .A3(new_n669), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n211), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR4_X1   g0494(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n215), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT89), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n494), .B2(new_n341), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT89), .A4(G179), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n550), .A2(new_n554), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n600), .B1(new_n610), .B2(new_n252), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n537), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n701), .A2(new_n702), .A3(new_n703), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT90), .ZN(new_n709));
  INV_X1    g0509(.A(new_n611), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n703), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n578), .A2(KEYINPUT90), .A3(new_n611), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n494), .A2(new_n341), .A3(new_n537), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n578), .A2(new_n704), .A3(new_n537), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT30), .A3(new_n702), .A4(new_n701), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n708), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n717), .B2(new_n668), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n708), .A2(new_n714), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT91), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n708), .A2(new_n714), .A3(KEYINPUT91), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n716), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n668), .A2(KEYINPUT31), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n511), .A2(new_n629), .A3(new_n669), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n699), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n644), .A2(new_n669), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(new_n631), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n635), .A2(new_n618), .A3(new_n573), .A4(new_n582), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n583), .A2(new_n585), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n541), .A2(new_n584), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n540), .A2(new_n542), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n573), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n642), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n577), .A2(new_n580), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n555), .B1(new_n341), .B2(new_n703), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n634), .A4(new_n586), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT26), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n634), .B(KEYINPUT92), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n737), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n669), .B1(new_n732), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n727), .A2(new_n729), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n698), .B1(new_n746), .B2(G1), .ZN(G364));
  AND2_X1   g0547(.A1(new_n208), .A2(G13), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n207), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n693), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n676), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n674), .A2(new_n675), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n699), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n751), .B(KEYINPUT93), .Z(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n217), .B1(G20), .B2(new_n389), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n208), .A2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n361), .B1(new_n767), .B2(G329), .ZN(new_n768));
  INV_X1    g0568(.A(G303), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  NAND2_X1  g0572(.A1(G20), .A2(G179), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n765), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n261), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n772), .A2(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n341), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n764), .A2(new_n261), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n782), .A2(new_n604), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n771), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT98), .B(G326), .Z(new_n788));
  NAND3_X1  g0588(.A1(new_n774), .A2(new_n261), .A3(G200), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI221_X1 g0590(.A(new_n786), .B1(new_n787), .B2(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n361), .B1(new_n409), .B2(new_n783), .C1(new_n775), .C2(new_n397), .ZN(new_n792));
  INV_X1    g0592(.A(new_n777), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(G58), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  OR3_X1    g0595(.A1(new_n766), .A2(KEYINPUT32), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(KEYINPUT32), .B1(new_n766), .B2(new_n795), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(new_n263), .C2(new_n770), .ZN(new_n798));
  INV_X1    g0598(.A(new_n787), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(G50), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n789), .A2(new_n318), .B1(new_n782), .B2(new_n476), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT97), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n794), .A2(new_n800), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n763), .B1(new_n791), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n758), .A2(new_n762), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n211), .A2(new_n361), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(KEYINPUT94), .B2(G355), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(KEYINPUT94), .B2(G355), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n692), .A2(new_n273), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n216), .A2(new_n249), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n245), .C2(new_n249), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n812), .B(new_n815), .C1(G116), .C2(new_n211), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n761), .B(new_n806), .C1(new_n809), .C2(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n753), .A2(new_n755), .B1(new_n759), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n762), .A2(new_n756), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n761), .B1(new_n397), .B2(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n360), .B1(new_n766), .B2(new_n772), .C1(new_n782), .C2(new_n476), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n784), .A2(new_n789), .B1(new_n787), .B2(new_n769), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n471), .A2(new_n775), .B1(new_n777), .B2(new_n604), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n263), .A2(new_n783), .B1(new_n770), .B2(new_n409), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n775), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G143), .A2(new_n793), .B1(new_n827), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n787), .C1(new_n830), .C2(new_n789), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT34), .ZN(new_n832));
  INV_X1    g0632(.A(new_n783), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G68), .A2(new_n833), .B1(new_n781), .B2(G58), .ZN(new_n834));
  INV_X1    g0634(.A(G50), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n770), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n284), .B(new_n836), .C1(G132), .C2(new_n767), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n826), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n413), .B1(new_n404), .B2(new_n669), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n416), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n649), .A2(new_n669), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n821), .B1(new_n838), .B2(new_n763), .C1(new_n843), .C2(new_n757), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n728), .A2(new_n842), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT99), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n417), .A2(new_n669), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n644), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n644), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n727), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n752), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n852), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n844), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT100), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  OR3_X1    g0658(.A1(new_n215), .A2(new_n397), .A3(new_n313), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n201), .A2(G68), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n207), .B(G13), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT101), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n218), .A2(G116), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n567), .B2(KEYINPUT35), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(KEYINPUT35), .B2(new_n567), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT36), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  INV_X1    g0669(.A(new_n841), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n643), .A2(new_n638), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n848), .B1(new_n871), .B2(new_n732), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT99), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n644), .A2(new_n846), .A3(new_n848), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n445), .A2(KEYINPUT102), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n450), .A2(new_n669), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n449), .B2(new_n450), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n426), .C1(new_n441), .C2(new_n444), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n441), .A2(new_n444), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n451), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n877), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n869), .B1(new_n875), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n841), .B1(new_n849), .B2(new_n850), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(KEYINPUT103), .A3(new_n885), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n348), .A2(new_n344), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT16), .B1(new_n346), .B2(new_n347), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n311), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n666), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT75), .B1(new_n352), .B2(new_n353), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n356), .A2(new_n355), .A3(new_n357), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n898), .B2(new_n339), .ZN(new_n899));
  INV_X1    g0699(.A(new_n343), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n655), .A2(KEYINPUT104), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n349), .B(new_n311), .C1(new_n652), .C2(new_n653), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n655), .A2(new_n894), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n350), .B2(KEYINPUT104), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n893), .A2(new_n900), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n908), .A3(new_n895), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n904), .A2(new_n907), .B1(KEYINPUT37), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n890), .B1(new_n899), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n658), .B1(new_n896), .B2(new_n897), .ZN(new_n915));
  OAI211_X1 g0715(.A(KEYINPUT38), .B(new_n914), .C1(new_n915), .C2(new_n895), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n887), .A2(new_n889), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n666), .B1(new_n352), .B2(new_n353), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n903), .B1(new_n339), .B2(new_n647), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n655), .A2(new_n900), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n902), .A2(new_n921), .A3(new_n903), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n904), .A2(new_n907), .B1(KEYINPUT37), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n890), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n911), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n876), .A2(new_n880), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n927), .A2(new_n928), .A3(new_n669), .A4(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n918), .A2(new_n919), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n453), .B1(new_n745), .B2(new_n729), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n660), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n931), .B(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n656), .A2(new_n657), .A3(new_n356), .A4(new_n357), .ZN(new_n935));
  INV_X1    g0735(.A(new_n903), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n902), .A2(new_n921), .A3(new_n903), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n938), .A2(new_n905), .B1(new_n913), .B2(new_n906), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n895), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n910), .B1(new_n359), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n942), .B2(KEYINPUT38), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n717), .A2(new_n724), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n718), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n726), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n842), .B1(new_n881), .B2(new_n884), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT40), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n917), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n453), .A2(new_n946), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT105), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n699), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n953), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n934), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n207), .B2(new_n748), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n934), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n868), .B1(new_n959), .B2(new_n960), .ZN(G367));
  AOI21_X1  g0761(.A(new_n808), .B1(new_n692), .B2(new_n524), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n813), .A2(new_n238), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n761), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n758), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n734), .A2(new_n669), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n639), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n640), .B2(new_n966), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n770), .A2(new_n471), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT46), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT110), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(KEYINPUT46), .B2(new_n969), .C1(new_n604), .C2(new_n789), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT111), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(KEYINPUT111), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n784), .A2(new_n775), .B1(new_n777), .B2(new_n769), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G97), .A2(new_n833), .B1(new_n781), .B2(G107), .ZN(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n284), .C1(new_n977), .C2(new_n766), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n975), .B(new_n978), .C1(G311), .C2(new_n799), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n973), .A2(new_n974), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT112), .Z(new_n981));
  INV_X1    g0781(.A(new_n201), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G150), .A2(new_n793), .B1(new_n827), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n781), .A2(G68), .ZN(new_n984));
  INV_X1    g0784(.A(new_n770), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n985), .A2(G58), .B1(new_n767), .B2(G137), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G143), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n988), .A2(new_n787), .B1(new_n789), .B2(new_n795), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n361), .B1(new_n783), .B2(new_n397), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT113), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n987), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n981), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n993), .A2(KEYINPUT47), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n762), .B1(new_n993), .B2(KEYINPUT47), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n964), .B1(new_n965), .B2(new_n968), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n683), .A2(new_n681), .ZN(new_n997));
  INV_X1    g0797(.A(new_n686), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n676), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n676), .A2(new_n999), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n746), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n738), .A2(new_n668), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n632), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n736), .A2(new_n668), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n690), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(KEYINPUT107), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1007), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n687), .A2(KEYINPUT107), .A3(new_n689), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1012), .A3(KEYINPUT45), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT107), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n690), .B2(new_n1007), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1014), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1010), .B1(new_n687), .B2(new_n689), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1013), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT108), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n1022), .A3(new_n684), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1021), .A2(new_n684), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n684), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT108), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1003), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n746), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n693), .B(KEYINPUT41), .Z(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n750), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n687), .A2(new_n1007), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT42), .Z(new_n1033));
  OAI21_X1  g0833(.A(new_n573), .B1(new_n1005), .B2(new_n624), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n669), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n1036), .A2(KEYINPUT106), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT106), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n684), .A2(new_n1007), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n996), .B1(new_n1031), .B2(new_n1044), .ZN(G387));
  OAI22_X1  g0845(.A1(new_n810), .A2(new_n695), .B1(G107), .B2(new_n211), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n235), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n300), .A2(new_n835), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n695), .B(new_n249), .C1(new_n318), .C2(new_n397), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n813), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1047), .A2(G45), .B1(KEYINPUT114), .B2(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1046), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n760), .B1(new_n1054), .B2(new_n808), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n782), .A2(new_n395), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G97), .B2(new_n833), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n397), .B2(new_n770), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n789), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1058), .B1(new_n300), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n273), .B1(new_n830), .B2(new_n766), .C1(new_n775), .C2(new_n318), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G50), .B2(new_n793), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(new_n795), .C2(new_n787), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n782), .A2(new_n784), .B1(new_n770), .B2(new_n604), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G303), .A2(new_n827), .B1(new_n793), .B2(G317), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n772), .B2(new_n789), .C1(new_n778), .C2(new_n787), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT49), .Z(new_n1070));
  OAI221_X1 g0870(.A(new_n284), .B1(new_n783), .B2(new_n471), .C1(new_n766), .C2(new_n788), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1063), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1055), .B1(new_n1072), .B2(new_n762), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n997), .B2(new_n965), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT115), .Z(new_n1075));
  AND2_X1   g0875(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1075), .B1(new_n750), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n693), .B1(new_n1076), .B2(new_n746), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1003), .B2(new_n1078), .ZN(G393));
  OAI21_X1  g0879(.A(new_n809), .B1(new_n476), .B2(new_n211), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n242), .A2(new_n692), .A3(new_n273), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n760), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n360), .B1(new_n766), .B2(new_n778), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n782), .A2(new_n471), .B1(new_n770), .B2(new_n784), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(G107), .C2(new_n833), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n604), .B2(new_n775), .C1(new_n769), .C2(new_n789), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n787), .A2(new_n977), .B1(new_n777), .B2(new_n772), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT52), .Z(new_n1088));
  OAI22_X1  g0888(.A1(new_n787), .A2(new_n830), .B1(new_n777), .B2(new_n795), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT51), .Z(new_n1090));
  NOR2_X1   g0890(.A1(new_n783), .A2(new_n263), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n782), .A2(new_n397), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G68), .C2(new_n985), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1059), .A2(new_n982), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n827), .A2(new_n300), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n284), .B1(G143), .B2(new_n767), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1086), .A2(new_n1088), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1082), .B1(new_n1098), .B2(new_n762), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1007), .B2(new_n965), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n749), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1002), .B(KEYINPUT109), .Z(new_n1103));
  AOI21_X1  g0903(.A(new_n694), .B1(new_n1103), .B2(new_n1101), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n1027), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  AOI21_X1  g0906(.A(new_n885), .B1(new_n727), .B2(new_n843), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n946), .A2(G330), .A3(new_n947), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n888), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n727), .A2(new_n843), .A3(new_n885), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n839), .A2(new_n416), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n841), .B1(new_n744), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n699), .B(new_n842), .C1(new_n726), .C2(new_n945), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1110), .B(new_n1113), .C1(new_n885), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n453), .A2(G330), .A3(new_n946), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n932), .A2(new_n1117), .A3(new_n660), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT116), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n888), .A2(new_n885), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n929), .A2(new_n669), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1121), .A2(new_n1122), .B1(new_n927), .B2(new_n928), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1112), .A2(new_n885), .B1(new_n669), .B2(new_n929), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n925), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1110), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1123), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1108), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n927), .A2(new_n928), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1122), .B1(new_n875), .B2(new_n886), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1132), .B2(new_n1125), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1120), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1108), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1125), .A3(new_n1110), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1118), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1136), .C1(KEYINPUT116), .C2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1138), .A3(new_n693), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1135), .A2(new_n1136), .A3(new_n750), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1130), .A2(new_n756), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n820), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n760), .B1(new_n300), .B2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n360), .B1(new_n766), .B2(new_n604), .C1(new_n263), .C2(new_n770), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1144), .B(new_n1092), .C1(G68), .C2(new_n833), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G97), .A2(new_n827), .B1(new_n793), .B2(G116), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G107), .A2(new_n1059), .B1(new_n799), .B2(G283), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n361), .B1(new_n766), .B2(new_n1149), .C1(new_n782), .C2(new_n795), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n982), .B2(new_n833), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  AOI22_X1  g0952(.A1(new_n1059), .A2(G137), .B1(new_n827), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT117), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n985), .A2(G150), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1156), .A2(KEYINPUT53), .B1(new_n777), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(KEYINPUT53), .B2(new_n1156), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n799), .A2(G128), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1151), .A2(new_n1155), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1148), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1143), .B1(new_n1163), .B2(new_n762), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1141), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1140), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1139), .A2(new_n1166), .ZN(G378));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n380), .A2(new_n666), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n392), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n392), .A2(new_n1170), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1169), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n392), .A2(new_n1170), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n1171), .A3(new_n1168), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n953), .B2(G330), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n699), .B(new_n1177), .C1(new_n949), .C2(new_n952), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n931), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n885), .A2(new_n843), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n726), .B2(new_n945), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n925), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1184), .A2(KEYINPUT40), .B1(new_n917), .B2(new_n951), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1177), .B1(new_n1185), .B2(new_n699), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n930), .A2(new_n919), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n917), .A2(new_n951), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n950), .B1(new_n1183), .B2(new_n925), .ZN(new_n1189));
  OAI211_X1 g0989(.A(G330), .B(new_n1178), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n918), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1181), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1135), .A2(new_n1136), .A3(new_n1116), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1119), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n694), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1192), .A2(new_n1194), .A3(KEYINPUT121), .A4(KEYINPUT57), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1192), .A2(new_n1194), .A3(KEYINPUT57), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1197), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n751), .B1(new_n982), .B2(new_n1142), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n793), .A2(G128), .B1(new_n985), .B2(new_n1152), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT119), .Z(new_n1205));
  OAI22_X1  g1005(.A1(new_n830), .A2(new_n782), .B1(new_n775), .B2(new_n829), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G132), .B2(new_n1059), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(new_n1149), .C2(new_n787), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n795), .B2(new_n783), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n273), .A2(G41), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n835), .B1(G33), .B2(G41), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n833), .A2(G58), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n397), .B2(new_n770), .C1(new_n784), .C2(new_n766), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1214), .B1(new_n777), .B2(new_n409), .C1(new_n395), .C2(new_n775), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G97), .C2(new_n1059), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n984), .B1(new_n787), .B2(new_n471), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT118), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT58), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1216), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1224), .B2(new_n1223), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n762), .B1(new_n1213), .B2(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT120), .Z(new_n1228));
  AOI211_X1 g1028(.A(new_n1203), .B(new_n1228), .C1(new_n756), .C2(new_n1177), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1192), .B2(new_n750), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1202), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT122), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT122), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1202), .A2(new_n1233), .A3(new_n1230), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(G375));
  AND2_X1   g1036(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1118), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1137), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1030), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n886), .A2(new_n756), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n760), .B1(G68), .B2(new_n1142), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n360), .B1(new_n766), .B2(new_n769), .C1(new_n397), .C2(new_n783), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1243), .B(new_n1056), .C1(G97), .C2(new_n985), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G107), .A2(new_n827), .B1(new_n793), .B2(G283), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G116), .A2(new_n1059), .B1(new_n799), .B2(G294), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n799), .A2(G132), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT123), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1059), .A2(new_n1152), .B1(new_n793), .B2(G137), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT124), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1217), .B1(new_n782), .B2(new_n835), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G159), .B2(new_n985), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n284), .B1(G128), .B2(new_n767), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n830), .C2(new_n775), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1247), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1242), .B1(new_n1257), .B2(new_n762), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1116), .A2(new_n750), .B1(new_n1241), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1240), .A2(new_n1259), .ZN(G381));
  OAI211_X1 g1060(.A(new_n996), .B(new_n1105), .C1(new_n1031), .C2(new_n1044), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G378), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1139), .A2(KEYINPUT125), .A3(new_n1166), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(G393), .A2(G396), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1266), .A2(new_n857), .A3(new_n1259), .A4(new_n1240), .ZN(new_n1267));
  OR4_X1    g1067(.A1(G375), .A2(new_n1261), .A3(new_n1265), .A4(new_n1267), .ZN(G407));
  INV_X1    g1068(.A(new_n1265), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1235), .A2(G213), .A3(new_n667), .A4(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1270), .ZN(G409));
  NAND3_X1  g1071(.A1(new_n1202), .A2(G378), .A3(new_n1230), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1192), .A2(new_n1194), .A3(new_n1030), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1230), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1263), .A2(new_n1274), .A3(new_n1264), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT126), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1263), .A2(new_n1274), .A3(new_n1277), .A4(new_n1264), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1272), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n667), .A2(G213), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1238), .B1(new_n1281), .B2(new_n1137), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1237), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n693), .A3(new_n1283), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1284), .A2(G384), .A3(new_n1259), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1284), .B2(new_n1259), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1279), .A2(new_n1280), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT62), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n667), .A2(G213), .A3(G2897), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1287), .B(new_n1291), .Z(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1279), .A2(new_n1295), .A3(new_n1280), .A4(new_n1287), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1289), .A2(new_n1293), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1298), .A2(new_n1266), .A3(KEYINPUT127), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT127), .B1(new_n1298), .B2(new_n1266), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1261), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1044), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1029), .B1(new_n1027), .B2(new_n746), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n750), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1105), .B1(new_n1304), .B2(new_n996), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1299), .B1(new_n1301), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G387), .A2(G390), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1299), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1307), .A2(new_n1261), .A3(new_n1308), .A4(new_n1300), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1297), .A2(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1288), .A2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1279), .A2(KEYINPUT63), .A3(new_n1280), .A4(new_n1287), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1311), .A2(new_n1317), .ZN(G405));
  INV_X1    g1118(.A(new_n1287), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1232), .A2(new_n1234), .A3(new_n1269), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1320), .B2(new_n1272), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1272), .A3(new_n1319), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1312), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1323), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1310), .B1(new_n1325), .B2(new_n1321), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1326), .ZN(G402));
endmodule


