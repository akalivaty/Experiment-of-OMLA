

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795;

  NAND2_X1 U379 ( .A1(n411), .A2(G210), .ZN(n741) );
  NAND2_X1 U380 ( .A1(n422), .A2(KEYINPUT2), .ZN(n425) );
  NAND2_X1 U381 ( .A1(n359), .A2(n358), .ZN(n422) );
  INV_X1 U382 ( .A(n446), .ZN(n360) );
  NAND2_X1 U383 ( .A1(n385), .A2(n386), .ZN(n443) );
  AND2_X1 U384 ( .A1(n788), .A2(n444), .ZN(n388) );
  NOR2_X1 U385 ( .A1(n723), .A2(n649), .ZN(n362) );
  XNOR2_X1 U386 ( .A(n510), .B(n361), .ZN(n694) );
  XNOR2_X1 U387 ( .A(n511), .B(KEYINPUT1), .ZN(n361) );
  XNOR2_X1 U388 ( .A(n523), .B(n507), .ZN(n777) );
  BUF_X1 U389 ( .A(G143), .Z(n357) );
  XNOR2_X1 U390 ( .A(G116), .B(KEYINPUT3), .ZN(n470) );
  INV_X1 U391 ( .A(G953), .ZN(n781) );
  NAND2_X1 U392 ( .A1(n458), .A2(n457), .ZN(n674) );
  AND2_X2 U393 ( .A1(n462), .A2(n461), .ZN(n458) );
  XNOR2_X2 U394 ( .A(n499), .B(n520), .ZN(n568) );
  INV_X1 U395 ( .A(n657), .ZN(n358) );
  XNOR2_X2 U396 ( .A(n447), .B(n360), .ZN(n359) );
  XNOR2_X1 U397 ( .A(n362), .B(KEYINPUT34), .ZN(n638) );
  XNOR2_X2 U398 ( .A(n633), .B(KEYINPUT83), .ZN(n368) );
  XNOR2_X2 U399 ( .A(n514), .B(G134), .ZN(n523) );
  INV_X1 U400 ( .A(n696), .ZN(n652) );
  XNOR2_X1 U401 ( .A(n777), .B(G146), .ZN(n574) );
  XNOR2_X2 U402 ( .A(n452), .B(n519), .ZN(n463) );
  XNOR2_X2 U403 ( .A(n471), .B(n569), .ZN(n452) );
  INV_X1 U404 ( .A(n534), .ZN(n466) );
  XOR2_X1 U405 ( .A(G125), .B(G146), .Z(n534) );
  INV_X1 U406 ( .A(KEYINPUT72), .ZN(n495) );
  INV_X1 U407 ( .A(KEYINPUT35), .ZN(n366) );
  AND2_X1 U408 ( .A1(n644), .A2(n449), .ZN(n448) );
  NAND2_X1 U409 ( .A1(n611), .A2(n684), .ZN(n428) );
  XNOR2_X1 U410 ( .A(n599), .B(n598), .ZN(n710) );
  XNOR2_X1 U411 ( .A(n748), .B(n747), .ZN(n750) );
  XNOR2_X1 U412 ( .A(n467), .B(n534), .ZN(n779) );
  XNOR2_X1 U413 ( .A(n768), .B(n495), .ZN(n471) );
  XNOR2_X1 U414 ( .A(n470), .B(G119), .ZN(n499) );
  NOR2_X1 U415 ( .A1(n758), .A2(n759), .ZN(n760) );
  NOR2_X1 U416 ( .A1(n663), .A2(n759), .ZN(n665) );
  XNOR2_X1 U417 ( .A(n465), .B(n463), .ZN(n369) );
  INV_X1 U418 ( .A(n395), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n657), .B(n656), .ZN(n780) );
  NAND2_X1 U420 ( .A1(n365), .A2(n624), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n438), .B(n587), .ZN(n365) );
  XNOR2_X2 U422 ( .A(n367), .B(n366), .ZN(n788) );
  NAND2_X1 U423 ( .A1(n638), .A2(n637), .ZN(n367) );
  XNOR2_X2 U424 ( .A(n604), .B(KEYINPUT39), .ZN(n611) );
  XNOR2_X2 U425 ( .A(n428), .B(n427), .ZN(n795) );
  XNOR2_X1 U426 ( .A(n463), .B(n465), .ZN(n738) );
  NAND2_X2 U427 ( .A1(n480), .A2(n478), .ZN(n438) );
  XNOR2_X1 U428 ( .A(n509), .B(n494), .ZN(n745) );
  XNOR2_X1 U429 ( .A(n574), .B(n508), .ZN(n509) );
  INV_X1 U430 ( .A(KEYINPUT102), .ZN(n598) );
  INV_X1 U431 ( .A(KEYINPUT84), .ZN(n483) );
  NAND2_X1 U432 ( .A1(n445), .A2(KEYINPUT44), .ZN(n444) );
  AND2_X1 U433 ( .A1(n593), .A2(n592), .ZN(n416) );
  XNOR2_X1 U434 ( .A(G902), .B(KEYINPUT15), .ZN(n548) );
  XOR2_X1 U435 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n516) );
  XOR2_X1 U436 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n513) );
  NAND2_X1 U437 ( .A1(n371), .A2(n658), .ZN(n486) );
  INV_X1 U438 ( .A(KEYINPUT5), .ZN(n571) );
  XNOR2_X1 U439 ( .A(n775), .B(G101), .ZN(n569) );
  XOR2_X1 U440 ( .A(G137), .B(G131), .Z(n507) );
  XNOR2_X1 U441 ( .A(n437), .B(n436), .ZN(n467) );
  INV_X1 U442 ( .A(G140), .ZN(n436) );
  XNOR2_X1 U443 ( .A(KEYINPUT69), .B(KEYINPUT10), .ZN(n437) );
  XNOR2_X1 U444 ( .A(G128), .B(G119), .ZN(n553) );
  XNOR2_X1 U445 ( .A(n501), .B(G137), .ZN(n500) );
  INV_X1 U446 ( .A(G110), .ZN(n501) );
  XNOR2_X1 U447 ( .A(n503), .B(n552), .ZN(n502) );
  INV_X1 U448 ( .A(KEYINPUT24), .ZN(n552) );
  XNOR2_X1 U449 ( .A(KEYINPUT91), .B(KEYINPUT23), .ZN(n503) );
  XNOR2_X1 U450 ( .A(n434), .B(n531), .ZN(n555) );
  XNOR2_X1 U451 ( .A(n530), .B(n435), .ZN(n434) );
  INV_X1 U452 ( .A(KEYINPUT79), .ZN(n435) );
  XNOR2_X1 U453 ( .A(n557), .B(n374), .ZN(n505) );
  INV_X1 U454 ( .A(KEYINPUT22), .ZN(n497) );
  XNOR2_X1 U455 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n605) );
  OR2_X1 U456 ( .A1(G902), .A2(G237), .ZN(n522) );
  INV_X1 U457 ( .A(n482), .ZN(n481) );
  AND2_X1 U458 ( .A1(n707), .A2(n483), .ZN(n482) );
  XNOR2_X1 U459 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U460 ( .A(n420), .B(n419), .ZN(n698) );
  XNOR2_X1 U461 ( .A(KEYINPUT21), .B(KEYINPUT94), .ZN(n419) );
  NAND2_X1 U462 ( .A1(n551), .A2(G221), .ZN(n420) );
  XNOR2_X1 U463 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n775) );
  NAND2_X1 U464 ( .A1(n442), .A2(n440), .ZN(n439) );
  AND2_X1 U465 ( .A1(n441), .A2(KEYINPUT73), .ZN(n440) );
  INV_X1 U466 ( .A(KEYINPUT44), .ZN(n441) );
  XOR2_X1 U467 ( .A(KEYINPUT97), .B(G104), .Z(n542) );
  XNOR2_X1 U468 ( .A(G113), .B(G122), .ZN(n541) );
  XNOR2_X1 U469 ( .A(KEYINPUT95), .B(KEYINPUT12), .ZN(n537) );
  INV_X1 U470 ( .A(KEYINPUT45), .ZN(n446) );
  INV_X1 U471 ( .A(n548), .ZN(n658) );
  XNOR2_X1 U472 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U473 ( .A1(G237), .A2(G234), .ZN(n558) );
  XNOR2_X1 U474 ( .A(n492), .B(n491), .ZN(n723) );
  INV_X1 U475 ( .A(KEYINPUT33), .ZN(n491) );
  XNOR2_X1 U476 ( .A(n646), .B(KEYINPUT105), .ZN(n493) );
  XNOR2_X1 U477 ( .A(n575), .B(n573), .ZN(n430) );
  XNOR2_X1 U478 ( .A(n572), .B(n571), .ZN(n573) );
  INV_X1 U479 ( .A(G104), .ZN(n472) );
  XNOR2_X1 U480 ( .A(KEYINPUT16), .B(G122), .ZN(n521) );
  XNOR2_X1 U481 ( .A(G107), .B(KEYINPUT9), .ZN(n524) );
  XOR2_X1 U482 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n525) );
  XNOR2_X1 U483 ( .A(G116), .B(G122), .ZN(n527) );
  XNOR2_X1 U484 ( .A(n581), .B(n580), .ZN(n584) );
  XNOR2_X1 U485 ( .A(n579), .B(KEYINPUT110), .ZN(n580) );
  AND2_X1 U486 ( .A1(n418), .A2(n392), .ZN(n594) );
  XNOR2_X1 U487 ( .A(n547), .B(n469), .ZN(n597) );
  XNOR2_X1 U488 ( .A(KEYINPUT13), .B(G475), .ZN(n469) );
  XNOR2_X1 U489 ( .A(n556), .B(n372), .ZN(n756) );
  NOR2_X1 U490 ( .A1(G952), .A2(n781), .ZN(n759) );
  INV_X1 U491 ( .A(KEYINPUT40), .ZN(n427) );
  INV_X1 U492 ( .A(KEYINPUT36), .ZN(n407) );
  NAND2_X1 U493 ( .A1(n632), .A2(KEYINPUT32), .ZN(n460) );
  NOR2_X1 U494 ( .A1(n632), .A2(KEYINPUT32), .ZN(n459) );
  NOR2_X1 U495 ( .A1(n370), .A2(n379), .ZN(n461) );
  INV_X1 U496 ( .A(KEYINPUT82), .ZN(n431) );
  AND2_X1 U497 ( .A1(n694), .A2(KEYINPUT104), .ZN(n370) );
  AND2_X1 U498 ( .A1(G210), .A2(n522), .ZN(n371) );
  AND2_X1 U499 ( .A1(n555), .A2(G221), .ZN(n372) );
  AND2_X1 U500 ( .A1(n487), .A2(n486), .ZN(n373) );
  XOR2_X1 U501 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n374) );
  NOR2_X1 U502 ( .A1(n612), .A2(n399), .ZN(n375) );
  AND2_X1 U503 ( .A1(n658), .A2(n732), .ZN(n376) );
  AND2_X1 U504 ( .A1(n416), .A2(n415), .ZN(n377) );
  NOR2_X1 U505 ( .A1(n707), .A2(n483), .ZN(n378) );
  NAND2_X1 U506 ( .A1(n696), .A2(n629), .ZN(n379) );
  OR2_X1 U507 ( .A1(n476), .A2(n378), .ZN(n380) );
  OR2_X1 U508 ( .A1(n658), .A2(n371), .ZN(n381) );
  XOR2_X1 U509 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n382) );
  XOR2_X1 U510 ( .A(n740), .B(n739), .Z(n383) );
  XOR2_X1 U511 ( .A(KEYINPUT48), .B(KEYINPUT70), .Z(n384) );
  INV_X1 U512 ( .A(KEYINPUT74), .ZN(n424) );
  NAND2_X1 U513 ( .A1(n368), .A2(n388), .ZN(n385) );
  OR2_X1 U514 ( .A1(n387), .A2(n445), .ZN(n386) );
  INV_X1 U515 ( .A(n444), .ZN(n387) );
  NAND2_X1 U516 ( .A1(n504), .A2(n620), .ZN(n657) );
  XNOR2_X2 U517 ( .A(n617), .B(KEYINPUT38), .ZN(n708) );
  OR2_X1 U518 ( .A1(n640), .A2(n389), .ZN(n457) );
  OR2_X1 U519 ( .A1(n694), .A2(KEYINPUT104), .ZN(n389) );
  NAND2_X1 U520 ( .A1(n368), .A2(n788), .ZN(n390) );
  BUF_X1 U521 ( .A(n723), .Z(n391) );
  XNOR2_X1 U522 ( .A(n510), .B(n511), .ZN(n392) );
  NOR2_X2 U523 ( .A1(n682), .A2(n712), .ZN(n608) );
  XNOR2_X1 U524 ( .A(n364), .B(n382), .ZN(n393) );
  XNOR2_X1 U525 ( .A(n498), .B(n382), .ZN(n645) );
  NOR2_X1 U526 ( .A1(n650), .A2(n583), .ZN(n468) );
  AND2_X1 U527 ( .A1(n485), .A2(KEYINPUT84), .ZN(n479) );
  AND2_X1 U528 ( .A1(n369), .A2(n394), .ZN(n477) );
  AND2_X1 U529 ( .A1(n371), .A2(n482), .ZN(n394) );
  NAND2_X1 U530 ( .A1(n780), .A2(n424), .ZN(n396) );
  NAND2_X1 U531 ( .A1(n395), .A2(KEYINPUT74), .ZN(n397) );
  NAND2_X1 U532 ( .A1(n396), .A2(n397), .ZN(n421) );
  INV_X1 U533 ( .A(n780), .ZN(n395) );
  BUF_X1 U534 ( .A(n574), .Z(n398) );
  NAND2_X1 U535 ( .A1(n480), .A2(n478), .ZN(n399) );
  NAND2_X1 U536 ( .A1(n693), .A2(n694), .ZN(n646) );
  XNOR2_X1 U537 ( .A(n399), .B(n587), .ZN(n400) );
  XNOR2_X1 U538 ( .A(n438), .B(n587), .ZN(n625) );
  XNOR2_X1 U539 ( .A(n412), .B(n384), .ZN(n504) );
  NAND2_X1 U540 ( .A1(n377), .A2(n413), .ZN(n412) );
  NAND2_X1 U541 ( .A1(n443), .A2(n439), .ZN(n401) );
  NAND2_X1 U542 ( .A1(n443), .A2(n439), .ZN(n451) );
  XNOR2_X1 U543 ( .A(n432), .B(n431), .ZN(n641) );
  XNOR2_X1 U544 ( .A(n464), .B(n502), .ZN(n554) );
  XNOR2_X1 U545 ( .A(n500), .B(n553), .ZN(n464) );
  NAND2_X1 U546 ( .A1(n458), .A2(n457), .ZN(n402) );
  AND2_X2 U547 ( .A1(n426), .A2(n376), .ZN(n408) );
  NAND2_X1 U548 ( .A1(n423), .A2(n425), .ZN(n403) );
  NAND2_X1 U549 ( .A1(n425), .A2(n423), .ZN(n426) );
  XNOR2_X1 U550 ( .A(n414), .B(n605), .ZN(n413) );
  NAND2_X1 U551 ( .A1(n455), .A2(n453), .ZN(n404) );
  NAND2_X1 U552 ( .A1(n455), .A2(n453), .ZN(n789) );
  NAND2_X1 U553 ( .A1(n454), .A2(n459), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n405), .B(n406), .ZN(n752) );
  XNOR2_X1 U555 ( .A(n523), .B(n529), .ZN(n405) );
  AND2_X1 U556 ( .A1(G217), .A2(n555), .ZN(n406) );
  XNOR2_X1 U557 ( .A(n407), .B(n375), .ZN(n578) );
  AND2_X2 U558 ( .A1(n403), .A2(n376), .ZN(n411) );
  NAND2_X1 U559 ( .A1(n401), .A2(n448), .ZN(n409) );
  XNOR2_X1 U560 ( .A(n409), .B(n446), .ZN(n410) );
  NAND2_X1 U561 ( .A1(n408), .A2(G217), .ZN(n757) );
  NAND2_X1 U562 ( .A1(n411), .A2(G475), .ZN(n749) );
  NAND2_X1 U563 ( .A1(n408), .A2(G472), .ZN(n662) );
  NAND2_X1 U564 ( .A1(n408), .A2(G478), .ZN(n753) );
  NAND2_X1 U565 ( .A1(n408), .A2(G469), .ZN(n490) );
  NOR2_X2 U566 ( .A1(n795), .A2(n792), .ZN(n414) );
  NAND2_X1 U567 ( .A1(n610), .A2(n609), .ZN(n415) );
  XNOR2_X2 U568 ( .A(n417), .B(KEYINPUT76), .ZN(n682) );
  NAND2_X1 U569 ( .A1(n594), .A2(n400), .ZN(n417) );
  XNOR2_X1 U570 ( .A(n590), .B(KEYINPUT28), .ZN(n418) );
  NAND2_X1 U571 ( .A1(n421), .A2(n727), .ZN(n423) );
  INV_X1 U572 ( .A(n425), .ZN(n729) );
  AND2_X1 U573 ( .A1(n456), .A2(n460), .ZN(n455) );
  NOR2_X1 U574 ( .A1(n751), .A2(n759), .ZN(n429) );
  NOR2_X1 U575 ( .A1(n742), .A2(n759), .ZN(n743) );
  XNOR2_X1 U576 ( .A(n429), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U577 ( .A(KEYINPUT73), .ZN(n445) );
  NOR2_X1 U578 ( .A1(n433), .A2(n584), .ZN(n603) );
  XNOR2_X1 U579 ( .A(n430), .B(n398), .ZN(n659) );
  NOR2_X1 U580 ( .A1(n640), .A2(n639), .ZN(n432) );
  NOR2_X1 U581 ( .A1(n655), .A2(n450), .ZN(n449) );
  XNOR2_X1 U582 ( .A(n468), .B(KEYINPUT75), .ZN(n433) );
  NAND2_X1 U583 ( .A1(n410), .A2(n727), .ZN(n732) );
  INV_X1 U584 ( .A(n390), .ZN(n442) );
  NAND2_X1 U585 ( .A1(n451), .A2(n448), .ZN(n447) );
  INV_X1 U586 ( .A(n666), .ZN(n450) );
  XNOR2_X1 U587 ( .A(n452), .B(G140), .ZN(n494) );
  INV_X1 U588 ( .A(n640), .ZN(n454) );
  NAND2_X1 U589 ( .A1(n640), .A2(KEYINPUT32), .ZN(n456) );
  NAND2_X1 U590 ( .A1(n789), .A2(n674), .ZN(n633) );
  NAND2_X1 U591 ( .A1(n640), .A2(KEYINPUT104), .ZN(n462) );
  NOR2_X2 U592 ( .A1(n745), .A2(G902), .ZN(n510) );
  NAND2_X1 U593 ( .A1(n484), .A2(n482), .ZN(n474) );
  XNOR2_X2 U594 ( .A(n767), .B(n466), .ZN(n465) );
  OR2_X2 U595 ( .A1(n756), .A2(G902), .ZN(n506) );
  NAND2_X1 U596 ( .A1(n493), .A2(n639), .ZN(n492) );
  INV_X1 U597 ( .A(n710), .ZN(n627) );
  XNOR2_X1 U598 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X2 U599 ( .A(n473), .B(n472), .ZN(n768) );
  XNOR2_X2 U600 ( .A(G107), .B(G110), .ZN(n473) );
  AND2_X2 U601 ( .A1(n475), .A2(n474), .ZN(n480) );
  NOR2_X1 U602 ( .A1(n477), .A2(n380), .ZN(n475) );
  NOR2_X1 U603 ( .A1(n481), .A2(n486), .ZN(n476) );
  NAND2_X1 U604 ( .A1(n373), .A2(n485), .ZN(n595) );
  NAND2_X1 U605 ( .A1(n479), .A2(n373), .ZN(n478) );
  INV_X1 U606 ( .A(n485), .ZN(n484) );
  OR2_X2 U607 ( .A1(n738), .A2(n381), .ZN(n485) );
  NAND2_X1 U608 ( .A1(n369), .A2(n371), .ZN(n487) );
  NOR2_X1 U609 ( .A1(n488), .A2(n759), .ZN(G54) );
  XNOR2_X1 U610 ( .A(n490), .B(n489), .ZN(n488) );
  XNOR2_X1 U611 ( .A(n745), .B(n744), .ZN(n489) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n746) );
  XNOR2_X2 U613 ( .A(n496), .B(n497), .ZN(n640) );
  NOR2_X2 U614 ( .A1(n645), .A2(n628), .ZN(n496) );
  NAND2_X1 U615 ( .A1(n625), .A2(n624), .ZN(n498) );
  XNOR2_X2 U616 ( .A(n568), .B(n521), .ZN(n767) );
  XNOR2_X2 U617 ( .A(n506), .B(n505), .ZN(n629) );
  XNOR2_X1 U618 ( .A(n741), .B(n383), .ZN(n742) );
  XNOR2_X1 U619 ( .A(KEYINPUT71), .B(G113), .ZN(n520) );
  XNOR2_X1 U620 ( .A(n518), .B(n517), .ZN(n519) );
  INV_X1 U621 ( .A(KEYINPUT81), .ZN(n656) );
  INV_X1 U622 ( .A(n636), .ZN(n637) );
  XNOR2_X1 U623 ( .A(n659), .B(n660), .ZN(n661) );
  XNOR2_X1 U624 ( .A(n662), .B(n661), .ZN(n663) );
  INV_X1 U625 ( .A(n694), .ZN(n643) );
  INV_X1 U626 ( .A(G469), .ZN(n511) );
  XNOR2_X2 U627 ( .A(G128), .B(G143), .ZN(n514) );
  AND2_X1 U628 ( .A1(G227), .A2(n781), .ZN(n508) );
  NAND2_X1 U629 ( .A1(G224), .A2(n781), .ZN(n512) );
  XNOR2_X1 U630 ( .A(n513), .B(n512), .ZN(n518) );
  INV_X1 U631 ( .A(n514), .ZN(n515) );
  NAND2_X1 U632 ( .A1(G214), .A2(n522), .ZN(n707) );
  XNOR2_X1 U633 ( .A(KEYINPUT101), .B(G478), .ZN(n533) );
  XNOR2_X1 U634 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U635 ( .A(n526), .B(KEYINPUT7), .Z(n528) );
  XNOR2_X1 U636 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U637 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n531) );
  NAND2_X1 U638 ( .A1(G234), .A2(n781), .ZN(n530) );
  NOR2_X1 U639 ( .A1(G902), .A2(n752), .ZN(n532) );
  XNOR2_X1 U640 ( .A(n533), .B(n532), .ZN(n596) );
  INV_X1 U641 ( .A(n596), .ZN(n586) );
  XNOR2_X1 U642 ( .A(n779), .B(n357), .ZN(n546) );
  XOR2_X1 U643 ( .A(G131), .B(KEYINPUT11), .Z(n536) );
  NOR2_X1 U644 ( .A1(G953), .A2(G237), .ZN(n570) );
  NAND2_X1 U645 ( .A1(n570), .A2(G214), .ZN(n535) );
  XNOR2_X1 U646 ( .A(n535), .B(n536), .ZN(n540) );
  XOR2_X1 U647 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n538) );
  XNOR2_X1 U648 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U649 ( .A(n540), .B(n539), .Z(n544) );
  XNOR2_X1 U650 ( .A(n542), .B(n541), .ZN(n543) );
  NOR2_X1 U651 ( .A1(G902), .A2(n746), .ZN(n547) );
  NAND2_X1 U652 ( .A1(n586), .A2(n597), .ZN(n681) );
  INV_X1 U653 ( .A(n681), .ZN(n684) );
  NAND2_X1 U654 ( .A1(n548), .A2(G234), .ZN(n550) );
  XNOR2_X1 U655 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n549) );
  INV_X1 U656 ( .A(n698), .ZN(n626) );
  NAND2_X1 U657 ( .A1(n551), .A2(G217), .ZN(n557) );
  XOR2_X1 U658 ( .A(n779), .B(n554), .Z(n556) );
  AND2_X1 U659 ( .A1(n626), .A2(n629), .ZN(n567) );
  XNOR2_X1 U660 ( .A(n558), .B(KEYINPUT14), .ZN(n560) );
  NAND2_X1 U661 ( .A1(G952), .A2(n560), .ZN(n721) );
  NOR2_X1 U662 ( .A1(G953), .A2(n721), .ZN(n559) );
  XOR2_X1 U663 ( .A(KEYINPUT88), .B(n559), .Z(n623) );
  INV_X1 U664 ( .A(n623), .ZN(n565) );
  NAND2_X1 U665 ( .A1(n560), .A2(G902), .ZN(n561) );
  XNOR2_X1 U666 ( .A(n561), .B(KEYINPUT89), .ZN(n621) );
  NAND2_X1 U667 ( .A1(G953), .A2(n621), .ZN(n562) );
  NOR2_X1 U668 ( .A1(G900), .A2(n562), .ZN(n563) );
  XNOR2_X1 U669 ( .A(n563), .B(KEYINPUT106), .ZN(n564) );
  NOR2_X1 U670 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U671 ( .A(KEYINPUT77), .B(n566), .ZN(n582) );
  NAND2_X1 U672 ( .A1(n567), .A2(n582), .ZN(n589) );
  XNOR2_X1 U673 ( .A(n568), .B(n569), .ZN(n575) );
  NAND2_X1 U674 ( .A1(n570), .A2(G210), .ZN(n572) );
  NOR2_X1 U675 ( .A1(n659), .A2(G902), .ZN(n576) );
  XNOR2_X2 U676 ( .A(n576), .B(G472), .ZN(n696) );
  XOR2_X1 U677 ( .A(KEYINPUT6), .B(n696), .Z(n634) );
  NOR2_X1 U678 ( .A1(n589), .A2(n634), .ZN(n577) );
  NAND2_X1 U679 ( .A1(n684), .A2(n577), .ZN(n612) );
  NOR2_X1 U680 ( .A1(n643), .A2(n578), .ZN(n690) );
  NAND2_X1 U681 ( .A1(n596), .A2(n597), .ZN(n636) );
  NAND2_X1 U682 ( .A1(n652), .A2(n707), .ZN(n581) );
  XOR2_X1 U683 ( .A(KEYINPUT30), .B(KEYINPUT109), .Z(n579) );
  INV_X1 U684 ( .A(n582), .ZN(n583) );
  NOR2_X2 U685 ( .A1(n629), .A2(n698), .ZN(n693) );
  NAND2_X1 U686 ( .A1(n392), .A2(n693), .ZN(n650) );
  NAND2_X1 U687 ( .A1(n595), .A2(n603), .ZN(n585) );
  NOR2_X1 U688 ( .A1(n636), .A2(n585), .ZN(n679) );
  NOR2_X1 U689 ( .A1(n690), .A2(n679), .ZN(n593) );
  NOR2_X1 U690 ( .A1(n597), .A2(n586), .ZN(n687) );
  NOR2_X1 U691 ( .A1(n684), .A2(n687), .ZN(n712) );
  XNOR2_X1 U692 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n587) );
  NOR2_X1 U693 ( .A1(n589), .A2(n696), .ZN(n590) );
  NOR2_X1 U694 ( .A1(n682), .A2(KEYINPUT78), .ZN(n591) );
  NAND2_X1 U695 ( .A1(n712), .A2(n591), .ZN(n592) );
  INV_X1 U696 ( .A(n594), .ZN(n601) );
  INV_X1 U697 ( .A(n595), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U699 ( .A1(n597), .A2(n596), .ZN(n599) );
  NOR2_X1 U700 ( .A1(n711), .A2(n710), .ZN(n600) );
  XNOR2_X1 U701 ( .A(n600), .B(KEYINPUT41), .ZN(n722) );
  NOR2_X1 U702 ( .A1(n601), .A2(n722), .ZN(n602) );
  XNOR2_X1 U703 ( .A(n602), .B(KEYINPUT42), .ZN(n792) );
  NAND2_X1 U704 ( .A1(n708), .A2(n603), .ZN(n604) );
  INV_X1 U705 ( .A(KEYINPUT47), .ZN(n607) );
  NAND2_X1 U706 ( .A1(n608), .A2(KEYINPUT78), .ZN(n606) );
  NAND2_X1 U707 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U708 ( .A1(n608), .A2(KEYINPUT47), .ZN(n609) );
  NAND2_X1 U709 ( .A1(n611), .A2(n687), .ZN(n692) );
  XOR2_X1 U710 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n615) );
  NOR2_X1 U711 ( .A1(n612), .A2(n694), .ZN(n613) );
  NAND2_X1 U712 ( .A1(n613), .A2(n707), .ZN(n614) );
  XNOR2_X1 U713 ( .A(n615), .B(n614), .ZN(n616) );
  NAND2_X1 U714 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U715 ( .A(KEYINPUT108), .B(n618), .Z(n791) );
  INV_X1 U716 ( .A(n791), .ZN(n619) );
  AND2_X1 U717 ( .A1(n692), .A2(n619), .ZN(n620) );
  NOR2_X1 U718 ( .A1(G898), .A2(n781), .ZN(n771) );
  NAND2_X1 U719 ( .A1(n621), .A2(n771), .ZN(n622) );
  NAND2_X1 U720 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U721 ( .A1(n627), .A2(n626), .ZN(n628) );
  INV_X1 U722 ( .A(n634), .ZN(n639) );
  XOR2_X1 U723 ( .A(KEYINPUT103), .B(n629), .Z(n699) );
  INV_X1 U724 ( .A(n699), .ZN(n630) );
  NOR2_X1 U725 ( .A1(n643), .A2(n630), .ZN(n631) );
  NAND2_X1 U726 ( .A1(n634), .A2(n631), .ZN(n632) );
  XNOR2_X1 U727 ( .A(n393), .B(KEYINPUT90), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n390), .A2(KEYINPUT44), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n699), .A2(n641), .ZN(n642) );
  NAND2_X1 U730 ( .A1(n643), .A2(n642), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n712), .B(KEYINPUT78), .ZN(n654) );
  INV_X1 U732 ( .A(n393), .ZN(n647) );
  NOR2_X1 U733 ( .A1(n696), .A2(n646), .ZN(n704) );
  NAND2_X1 U734 ( .A1(n647), .A2(n704), .ZN(n648) );
  XNOR2_X1 U735 ( .A(n648), .B(KEYINPUT31), .ZN(n688) );
  OR2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n671) );
  NOR2_X1 U738 ( .A1(n688), .A2(n671), .ZN(n653) );
  NOR2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n655) );
  INV_X1 U740 ( .A(KEYINPUT2), .ZN(n727) );
  XOR2_X1 U741 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n660) );
  INV_X1 U742 ( .A(KEYINPUT63), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(G57) );
  XNOR2_X1 U744 ( .A(n666), .B(G101), .ZN(G3) );
  NAND2_X1 U745 ( .A1(n671), .A2(n684), .ZN(n667) );
  XNOR2_X1 U746 ( .A(n667), .B(G104), .ZN(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n669) );
  XNOR2_X1 U748 ( .A(G107), .B(KEYINPUT112), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U750 ( .A(KEYINPUT26), .B(n670), .Z(n673) );
  NAND2_X1 U751 ( .A1(n671), .A2(n687), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n673), .B(n672), .ZN(G9) );
  XNOR2_X1 U753 ( .A(n402), .B(G110), .ZN(G12) );
  INV_X1 U754 ( .A(n687), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n682), .A2(n675), .ZN(n677) );
  XNOR2_X1 U756 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U758 ( .A(G128), .B(n678), .ZN(G30) );
  XNOR2_X1 U759 ( .A(n357), .B(n679), .ZN(n680) );
  XNOR2_X1 U760 ( .A(n680), .B(KEYINPUT115), .ZN(G45) );
  NOR2_X1 U761 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U762 ( .A(G146), .B(n683), .Z(G48) );
  NAND2_X1 U763 ( .A1(n688), .A2(n684), .ZN(n685) );
  XNOR2_X1 U764 ( .A(n685), .B(KEYINPUT116), .ZN(n686) );
  XNOR2_X1 U765 ( .A(G113), .B(n686), .ZN(G15) );
  NAND2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U767 ( .A(n689), .B(G116), .ZN(G18) );
  XNOR2_X1 U768 ( .A(G125), .B(n690), .ZN(n691) );
  XNOR2_X1 U769 ( .A(n691), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U770 ( .A(G134), .B(n692), .ZN(G36) );
  OR2_X1 U771 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U772 ( .A(n695), .B(KEYINPUT50), .ZN(n697) );
  NAND2_X1 U773 ( .A1(n697), .A2(n696), .ZN(n702) );
  NAND2_X1 U774 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U775 ( .A(KEYINPUT49), .B(n700), .ZN(n701) );
  NOR2_X1 U776 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U778 ( .A(KEYINPUT51), .B(n705), .Z(n706) );
  NOR2_X1 U779 ( .A1(n722), .A2(n706), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U781 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U783 ( .A(KEYINPUT117), .B(n713), .Z(n714) );
  NOR2_X1 U784 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U785 ( .A1(n716), .A2(n391), .ZN(n717) );
  NOR2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U787 ( .A(n719), .B(KEYINPUT52), .ZN(n720) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n725) );
  NOR2_X1 U789 ( .A1(n722), .A2(n391), .ZN(n724) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U791 ( .A(n726), .B(KEYINPUT118), .ZN(n735) );
  XOR2_X1 U792 ( .A(KEYINPUT80), .B(n363), .Z(n728) );
  NAND2_X1 U793 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U794 ( .A1(n729), .A2(KEYINPUT80), .ZN(n730) );
  NAND2_X1 U795 ( .A1(n731), .A2(n730), .ZN(n733) );
  NAND2_X1 U796 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U797 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U798 ( .A1(n736), .A2(G953), .ZN(n737) );
  XNOR2_X1 U799 ( .A(n737), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U800 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n740) );
  XNOR2_X1 U801 ( .A(n369), .B(KEYINPUT85), .ZN(n739) );
  XNOR2_X1 U802 ( .A(KEYINPUT56), .B(n743), .ZN(G51) );
  XOR2_X1 U803 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n744) );
  XNOR2_X1 U804 ( .A(KEYINPUT59), .B(KEYINPUT120), .ZN(n748) );
  XNOR2_X1 U805 ( .A(n746), .B(KEYINPUT119), .ZN(n747) );
  XNOR2_X1 U806 ( .A(n750), .B(n749), .ZN(n751) );
  XOR2_X1 U807 ( .A(n752), .B(KEYINPUT121), .Z(n754) );
  XNOR2_X1 U808 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U809 ( .A1(n759), .A2(n755), .ZN(G63) );
  XNOR2_X1 U810 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X1 U811 ( .A(n760), .B(KEYINPUT122), .ZN(G66) );
  OR2_X1 U812 ( .A1(G953), .A2(n410), .ZN(n765) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n762) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n762), .ZN(n763) );
  NAND2_X1 U815 ( .A1(n763), .A2(G898), .ZN(n764) );
  NAND2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n766), .B(KEYINPUT124), .ZN(n773) );
  XNOR2_X1 U818 ( .A(n767), .B(G101), .ZN(n769) );
  XNOR2_X1 U819 ( .A(n768), .B(n769), .ZN(n770) );
  NOR2_X1 U820 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U821 ( .A(n773), .B(n772), .Z(n774) );
  XNOR2_X1 U822 ( .A(KEYINPUT123), .B(n774), .ZN(G69) );
  XOR2_X1 U823 ( .A(KEYINPUT125), .B(n775), .Z(n776) );
  XNOR2_X1 U824 ( .A(n777), .B(n776), .ZN(n778) );
  XNOR2_X1 U825 ( .A(n779), .B(n778), .ZN(n783) );
  XNOR2_X1 U826 ( .A(n363), .B(n783), .ZN(n782) );
  NAND2_X1 U827 ( .A1(n782), .A2(n781), .ZN(n787) );
  XNOR2_X1 U828 ( .A(G227), .B(n783), .ZN(n784) );
  NAND2_X1 U829 ( .A1(n784), .A2(G900), .ZN(n785) );
  NAND2_X1 U830 ( .A1(n785), .A2(G953), .ZN(n786) );
  NAND2_X1 U831 ( .A1(n787), .A2(n786), .ZN(G72) );
  XNOR2_X1 U832 ( .A(n788), .B(G122), .ZN(G24) );
  XNOR2_X1 U833 ( .A(n404), .B(G119), .ZN(n790) );
  XNOR2_X1 U834 ( .A(n790), .B(KEYINPUT126), .ZN(G21) );
  XOR2_X1 U835 ( .A(G140), .B(n791), .Z(G42) );
  XNOR2_X1 U836 ( .A(G137), .B(KEYINPUT127), .ZN(n794) );
  BUF_X1 U837 ( .A(n792), .Z(n793) );
  XNOR2_X1 U838 ( .A(n794), .B(n793), .ZN(G39) );
  XOR2_X1 U839 ( .A(n795), .B(G131), .Z(G33) );
endmodule

