//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G78gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(G127gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n215), .B(new_n216), .C1(G1gat), .C2(new_n213), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n217), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n208), .B2(new_n207), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n212), .B(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G183gat), .B(G211gat), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n226), .B(new_n227), .Z(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n223), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G43gat), .B(G50gat), .Z(new_n231));
  INV_X1    g030(.A(KEYINPUT15), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G29gat), .A2(G36gat), .ZN(new_n234));
  INV_X1    g033(.A(G29gat), .ZN(new_n235));
  INV_X1    g034(.A(G36gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT14), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT14), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G29gat), .B2(G36gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n234), .B1(new_n240), .B2(KEYINPUT91), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT91), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n233), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n231), .A2(new_n232), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n234), .B(KEYINPUT92), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n231), .A2(new_n232), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n244), .A2(new_n240), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT17), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255));
  INV_X1    g054(.A(G85gat), .ZN(new_n256));
  INV_X1    g055(.A(G92gat), .ZN(new_n257));
  AOI22_X1  g056(.A1(KEYINPUT8), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G99gat), .B(G106gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n254), .B(new_n258), .C1(KEYINPUT96), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(KEYINPUT96), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n250), .A2(new_n252), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT96), .ZN(new_n264));
  INV_X1    g063(.A(new_n259), .ZN(new_n265));
  AOI211_X1 g064(.A(new_n264), .B(new_n265), .C1(new_n254), .C2(new_n258), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n260), .B1(KEYINPUT96), .B2(new_n259), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n248), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n268), .A2(KEYINPUT97), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT97), .B1(new_n268), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n263), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G134gat), .B(G162gat), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n273), .ZN(new_n275));
  XOR2_X1   g074(.A(G190gat), .B(G218gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT98), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n274), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n274), .B2(new_n275), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n262), .A2(new_n207), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT10), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n206), .B1(new_n267), .B2(new_n266), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT10), .B(new_n206), .C1(new_n267), .C2(new_n266), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G230gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n283), .A2(new_n285), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(new_n292), .ZN(new_n295));
  XNOR2_X1  g094(.A(G120gat), .B(G148gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G176gat), .B(G204gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n293), .B(new_n298), .C1(new_n294), .C2(new_n292), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT99), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT99), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n230), .A2(new_n282), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n307));
  INV_X1    g106(.A(G169gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n310), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  AND2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(KEYINPUT23), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT23), .ZN(new_n324));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT66), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n320), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n329), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(G183gat), .B(G190gat), .C1(KEYINPUT68), .C2(KEYINPUT24), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(new_n308), .A3(new_n309), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(KEYINPUT23), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n317), .A2(new_n334), .ZN(new_n347));
  AND4_X1   g146(.A1(new_n315), .A2(new_n342), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n335), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n351), .A2(KEYINPUT70), .B1(G127gat), .B2(G134gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(G127gat), .A2(G134gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n351), .B1(G113gat), .B2(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(G113gat), .A2(G120gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n352), .B(new_n354), .C1(new_n356), .C2(new_n358), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT26), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n363), .A3(new_n345), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n317), .B1(new_n310), .B2(KEYINPUT26), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT27), .B(G183gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT28), .B1(new_n367), .B2(new_n339), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n338), .A2(KEYINPUT27), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G183gat), .ZN(new_n371));
  AND4_X1   g170(.A1(KEYINPUT28), .A2(new_n369), .A3(new_n371), .A4(new_n339), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n366), .B(new_n329), .C1(new_n368), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT69), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n371), .A3(new_n339), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(KEYINPUT28), .A3(new_n339), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT69), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n329), .A4(new_n366), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n350), .A2(new_n362), .A3(new_n374), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n360), .A2(new_n361), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n374), .A2(new_n381), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n348), .B1(new_n333), .B2(new_n334), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT64), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G15gat), .B(G43gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(KEYINPUT33), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(KEYINPUT32), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n389), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n382), .B2(new_n386), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT32), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n400), .A2(KEYINPUT33), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n398), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n382), .A2(new_n386), .A3(new_n399), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT34), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n307), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n390), .A2(KEYINPUT32), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n410), .A3(new_n394), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n405), .B(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n411), .A2(KEYINPUT73), .A3(new_n413), .A4(new_n398), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT74), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n404), .A2(new_n406), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(new_n414), .A3(KEYINPUT74), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT36), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n413), .B1(new_n411), .B2(new_n398), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT72), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n415), .A2(new_n424), .A3(KEYINPUT36), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429));
  INV_X1    g228(.A(G141gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G148gat), .ZN(new_n431));
  INV_X1    g230(.A(G148gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G141gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n431), .A2(new_n433), .B1(KEYINPUT2), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  NOR2_X1   g235(.A1(G155gat), .A2(G162gat), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT81), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G162gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n225), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n431), .A2(new_n433), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT2), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n436), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n225), .A2(new_n439), .A3(KEYINPUT80), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(G155gat), .B2(G162gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n435), .A2(new_n443), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT3), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n383), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT81), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n441), .B1(new_n440), .B2(new_n434), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n435), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G141gat), .B(G148gat), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n450), .B(new_n434), .C1(KEYINPUT2), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n429), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(KEYINPUT5), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n456), .A2(new_n458), .A3(new_n360), .A4(new_n361), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n362), .A2(KEYINPUT83), .A3(new_n456), .A4(new_n458), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT4), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  INV_X1    g268(.A(new_n463), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n468), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n462), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n451), .B2(new_n362), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n479), .A3(new_n383), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n429), .B1(new_n467), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT5), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n429), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n459), .A2(new_n479), .A3(new_n383), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n479), .B1(new_n459), .B2(new_n383), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n466), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n470), .A2(new_n471), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n461), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT86), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  AOI211_X1 g298(.A(new_n499), .B(new_n496), .C1(new_n484), .C2(new_n491), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n476), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G1gat), .B(G29gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT0), .ZN(new_n503));
  XNOR2_X1  g302(.A(G57gat), .B(G85gat), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n503), .B(new_n504), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n476), .C1(new_n498), .C2(new_n500), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT29), .ZN(new_n511));
  INV_X1    g310(.A(new_n373), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n385), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G226gat), .A2(G233gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT77), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT22), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n517), .A2(KEYINPUT75), .B1(G211gat), .B2(G218gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(KEYINPUT75), .B2(new_n517), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(KEYINPUT76), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(KEYINPUT76), .ZN(new_n521));
  XNOR2_X1  g320(.A(G197gat), .B(G204gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G211gat), .B(G218gat), .Z(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n528), .A3(new_n514), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n350), .A2(new_n374), .A3(new_n381), .ZN(new_n530));
  INV_X1    g329(.A(new_n514), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n516), .A2(new_n527), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT37), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n385), .A2(new_n514), .A3(new_n512), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n531), .A2(KEYINPUT29), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n527), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n516), .A2(new_n538), .A3(new_n529), .A4(new_n532), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n534), .B1(new_n537), .B2(new_n527), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT38), .ZN(new_n544));
  XOR2_X1   g343(.A(G8gat), .B(G36gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT78), .ZN(new_n546));
  XNOR2_X1  g345(.A(G64gat), .B(G92gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n546), .B(new_n547), .Z(new_n548));
  NAND4_X1  g347(.A1(new_n540), .A2(new_n543), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n539), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n539), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT37), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n548), .A3(new_n540), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(KEYINPUT38), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n506), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n510), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G228gat), .A2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G22gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G50gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n538), .B1(KEYINPUT29), .B2(new_n460), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT29), .B1(new_n525), .B2(new_n526), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n459), .B1(new_n565), .B2(KEYINPUT3), .ZN(new_n566));
  XNOR2_X1  g365(.A(G78gat), .B(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n564), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n564), .B2(new_n566), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n563), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n566), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n567), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n564), .A2(new_n566), .A3(new_n568), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(new_n562), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n467), .A2(new_n481), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT39), .B1(new_n577), .B2(new_n485), .ZN(new_n578));
  OAI22_X1  g377(.A1(new_n474), .A2(new_n475), .B1(new_n460), .B2(new_n453), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(new_n485), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n582), .A3(new_n485), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n581), .A2(KEYINPUT40), .A3(new_n505), .A4(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n505), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(new_n580), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n551), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n550), .B1(new_n533), .B2(new_n539), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n589), .B2(new_n551), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n588), .B1(new_n551), .B2(new_n589), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n584), .A2(new_n587), .A3(new_n594), .A4(new_n507), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n558), .A2(new_n576), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n507), .A2(KEYINPUT88), .A3(new_n508), .A4(new_n509), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n501), .B(new_n506), .C1(new_n598), .C2(KEYINPUT6), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n594), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n428), .B(new_n596), .C1(new_n600), .C2(new_n576), .ZN(new_n601));
  AND4_X1   g400(.A1(new_n576), .A2(new_n415), .A3(new_n426), .A4(new_n424), .ZN(new_n602));
  INV_X1    g401(.A(new_n594), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n509), .A2(KEYINPUT88), .A3(new_n508), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n492), .A2(new_n497), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n499), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n497), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n505), .B1(new_n608), .B2(new_n476), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n599), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n602), .B(new_n603), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n420), .A2(KEYINPUT89), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n571), .A2(new_n575), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(new_n590), .A3(new_n593), .A4(new_n592), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n510), .B2(new_n557), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n423), .B1(new_n415), .B2(new_n416), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT89), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n419), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n601), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n221), .A2(new_n249), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n220), .A2(new_n633), .A3(new_n248), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n220), .B2(new_n248), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n220), .A2(new_n248), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT94), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n634), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n250), .A2(new_n221), .A3(new_n252), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT18), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n631), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n643), .A2(new_n644), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(KEYINPUT18), .A3(new_n638), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n651), .A2(new_n652), .A3(new_n640), .A4(new_n630), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n624), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n624), .A2(KEYINPUT95), .A3(new_n654), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n306), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n597), .A2(new_n599), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G8gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n659), .A2(new_n594), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n306), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT95), .B1(new_n624), .B2(new_n654), .ZN(new_n668));
  INV_X1    g467(.A(new_n654), .ZN(new_n669));
  AOI211_X1 g468(.A(new_n656), .B(new_n669), .C1(new_n601), .C2(new_n623), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n594), .B(new_n667), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n671), .A2(G8gat), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n671), .A2(new_n664), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT100), .B1(new_n675), .B2(KEYINPUT42), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n671), .A2(new_n677), .A3(new_n673), .A4(new_n664), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n674), .B1(new_n676), .B2(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  AND4_X1   g479(.A1(new_n620), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n620), .B1(new_n619), .B2(new_n419), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n659), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n427), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n421), .B2(new_n420), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n659), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n688), .B2(new_n680), .ZN(G1326gat));
  INV_X1    g488(.A(new_n576), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n659), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n282), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT44), .B1(new_n624), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  AOI211_X1 g495(.A(new_n696), .B(new_n282), .C1(new_n601), .C2(new_n623), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n305), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n230), .A2(new_n669), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n660), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n223), .B(new_n228), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n694), .A3(new_n305), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n657), .B2(new_n658), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n235), .A3(new_n661), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n707));
  AND2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n702), .B1(new_n708), .B2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n705), .A2(new_n236), .A3(new_n594), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n701), .B2(new_n603), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  INV_X1    g515(.A(new_n683), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n705), .B2(new_n718), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n558), .A2(new_n576), .A3(new_n595), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n576), .B1(new_n660), .B2(new_n603), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n686), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n683), .A2(new_n618), .B1(new_n612), .B2(KEYINPUT35), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n694), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n696), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n624), .A2(KEYINPUT44), .A3(new_n694), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n725), .A2(new_n686), .A3(new_n726), .A4(new_n700), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT103), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G43gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n727), .A2(KEYINPUT103), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n719), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n705), .A2(new_n718), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(G43gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n731), .A2(new_n736), .ZN(G1330gat));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n705), .A2(new_n738), .A3(new_n690), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n725), .A2(new_n690), .A3(new_n726), .A4(new_n700), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n739), .A2(KEYINPUT48), .A3(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1331gat));
  NOR4_X1   g545(.A1(new_n703), .A2(new_n654), .A3(new_n694), .A4(new_n305), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n624), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n660), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(G57gat), .Z(G1332gat));
  NAND2_X1  g549(.A1(new_n748), .A2(KEYINPUT104), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n624), .A2(new_n752), .A3(new_n747), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(new_n594), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  XNOR2_X1  g558(.A(new_n683), .B(KEYINPUT105), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n748), .A2(G71gat), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n751), .A2(new_n686), .A3(new_n753), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(G71gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n754), .A2(new_n690), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g565(.A1(new_n230), .A2(new_n654), .A3(new_n305), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n725), .A2(new_n661), .A3(new_n726), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G85gat), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n230), .A2(new_n654), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n694), .B(new_n770), .C1(new_n722), .C2(new_n723), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n624), .A2(KEYINPUT51), .A3(new_n694), .A4(new_n770), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n661), .A2(new_n256), .A3(new_n699), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n769), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT106), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n769), .B(new_n779), .C1(new_n775), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1336gat));
  NAND4_X1  g580(.A1(new_n725), .A2(new_n594), .A3(new_n726), .A4(new_n767), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n699), .A2(new_n594), .A3(new_n257), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT52), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n783), .B(new_n787), .C1(new_n775), .C2(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1337gat));
  NAND3_X1  g588(.A1(new_n698), .A2(new_n686), .A3(new_n767), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G99gat), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n717), .A2(G99gat), .A3(new_n305), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n775), .B2(new_n792), .ZN(G1338gat));
  NAND4_X1  g592(.A1(new_n725), .A2(new_n690), .A3(new_n726), .A4(new_n767), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n773), .A2(new_n774), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n305), .A2(new_n576), .A3(G106gat), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT107), .Z(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT53), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n698), .A2(KEYINPUT109), .A3(new_n690), .A4(new_n767), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n794), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n803), .A2(new_n805), .A3(G106gat), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT108), .B1(new_n796), .B2(new_n799), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n809), .B(new_n798), .C1(new_n773), .C2(new_n774), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n802), .B1(new_n806), .B2(new_n811), .ZN(G1339gat));
  NAND3_X1  g611(.A1(new_n286), .A2(new_n287), .A3(new_n291), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n293), .A2(new_n813), .A3(KEYINPUT54), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n291), .B1(new_n286), .B2(new_n287), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n816));
  AOI21_X1  g615(.A(new_n298), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n301), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(KEYINPUT111), .A3(new_n301), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n293), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n824));
  INV_X1    g623(.A(new_n816), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n299), .B1(new_n293), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n654), .A2(new_n821), .A3(new_n822), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT112), .B1(new_n637), .B2(new_n639), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n638), .B2(new_n650), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n637), .A2(KEYINPUT112), .A3(new_n639), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n629), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(new_n653), .A3(new_n304), .A4(new_n302), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n694), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n821), .A2(new_n822), .A3(new_n827), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n832), .B(new_n653), .C1(new_n280), .C2(new_n281), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n703), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n230), .A2(new_n669), .A3(new_n282), .A4(new_n305), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n660), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n603), .A3(new_n602), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT114), .Z(new_n842));
  INV_X1    g641(.A(G113gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n654), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n838), .A2(new_n839), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n576), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT113), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n661), .A2(new_n603), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n717), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n669), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n851), .ZN(G1340gat));
  INV_X1    g651(.A(G120gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n853), .A3(new_n699), .ZN(new_n854));
  OAI21_X1  g653(.A(G120gat), .B1(new_n850), .B2(new_n305), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n850), .B2(new_n703), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n703), .A2(G127gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n841), .B2(new_n858), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n850), .B2(new_n282), .ZN(new_n860));
  INV_X1    g659(.A(G134gat), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n594), .A2(new_n282), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n840), .A2(new_n861), .A3(new_n602), .A4(new_n862), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT56), .Z(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(KEYINPUT115), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n848), .A2(new_n686), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n690), .A2(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n824), .B2(new_n826), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n814), .A2(KEYINPUT117), .A3(new_n817), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n823), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n819), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n654), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n694), .B1(new_n877), .B2(new_n833), .ZN(new_n878));
  OAI22_X1  g677(.A1(new_n878), .A2(KEYINPUT118), .B1(new_n835), .B2(new_n836), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n880), .B(new_n694), .C1(new_n877), .C2(new_n833), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n703), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n882), .A2(new_n883), .B1(new_n669), .B2(new_n667), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT119), .B(new_n703), .C1(new_n879), .C2(new_n881), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n871), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n576), .B1(new_n838), .B2(new_n839), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n654), .B(new_n870), .C1(new_n886), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n686), .A2(KEYINPUT120), .A3(new_n576), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT120), .B1(new_n686), .B2(new_n576), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n893), .A2(new_n840), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(new_n430), .A3(new_n654), .A4(new_n603), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n892), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n703), .B1(new_n878), .B2(new_n837), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n839), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n576), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(KEYINPUT122), .A3(new_n839), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n888), .A2(new_n889), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n305), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n870), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n902), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n870), .B1(new_n886), .B2(new_n890), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n305), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n902), .A2(G148gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n603), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n699), .A2(new_n432), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n913), .A2(new_n917), .B1(new_n921), .B2(new_n922), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n914), .B2(new_n703), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n230), .A2(new_n225), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n918), .B2(new_n925), .ZN(G1346gat));
  OAI211_X1 g725(.A(new_n694), .B(new_n870), .C1(new_n886), .C2(new_n890), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n439), .B1(new_n927), .B2(KEYINPUT123), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(KEYINPUT123), .B2(new_n927), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n895), .A2(new_n439), .A3(new_n862), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1347gat));
  NAND4_X1  g730(.A1(new_n845), .A2(new_n660), .A3(new_n594), .A4(new_n602), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n654), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n760), .A2(new_n661), .A3(new_n603), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT113), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n846), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n669), .A2(new_n308), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  OR2_X1    g739(.A1(new_n935), .A2(new_n937), .ZN(new_n941));
  OAI21_X1  g740(.A(G176gat), .B1(new_n941), .B2(new_n305), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n933), .A2(new_n309), .A3(new_n699), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1349gat));
  OAI21_X1  g743(.A(G183gat), .B1(new_n941), .B2(new_n703), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n933), .A2(new_n367), .A3(new_n230), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n338), .B1(new_n938), .B2(new_n230), .ZN(new_n949));
  INV_X1    g748(.A(new_n947), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT60), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n948), .A2(new_n951), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n339), .A3(new_n694), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n694), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(G190gat), .ZN(new_n956));
  AOI211_X1 g755(.A(KEYINPUT61), .B(new_n339), .C1(new_n938), .C2(new_n694), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G1351gat));
  NOR3_X1   g757(.A1(new_n686), .A2(new_n661), .A3(new_n603), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n887), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n654), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n908), .A2(new_n909), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(new_n959), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n654), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  INV_X1    g765(.A(G204gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n967), .B1(new_n911), .B2(new_n959), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n887), .A2(new_n967), .A3(new_n959), .A4(new_n699), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n966), .B1(new_n968), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n699), .A3(new_n959), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G204gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(KEYINPUT125), .A3(new_n976), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n978), .A2(new_n981), .ZN(G1353gat));
  OAI211_X1 g781(.A(new_n230), .B(new_n959), .C1(new_n908), .C2(new_n909), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT63), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n983), .A2(new_n984), .A3(G211gat), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n703), .A2(G211gat), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n960), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n984), .B1(new_n983), .B2(G211gat), .ZN(new_n991));
  OAI21_X1  g790(.A(KEYINPUT127), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(new_n991), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n993), .A2(new_n994), .A3(new_n985), .A4(new_n989), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n992), .A2(new_n995), .ZN(G1354gat));
  INV_X1    g795(.A(G218gat), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n960), .A2(new_n997), .A3(new_n694), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n963), .A2(new_n694), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n999), .B2(new_n997), .ZN(G1355gat));
endmodule


