//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  XNOR2_X1  g001(.A(G141gat), .B(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n207), .C1(new_n203), .C2(KEYINPUT2), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n202), .B1(new_n213), .B2(KEYINPUT3), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT79), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n218));
  INV_X1    g017(.A(G127gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G134gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT70), .B(G134gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(new_n219), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT71), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT71), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n220), .C1(new_n221), .C2(new_n219), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  INV_X1    g025(.A(G120gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G113gat), .A2(G120gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n223), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n235));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n236), .A3(new_n229), .ZN(new_n237));
  XNOR2_X1  g036(.A(G127gat), .B(G134gat), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(KEYINPUT72), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n217), .A2(new_n218), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n222), .A2(KEYINPUT71), .B1(new_n232), .B2(new_n231), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n246), .A2(new_n225), .B1(new_n240), .B2(new_n239), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n211), .A2(new_n212), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AND4_X1   g048(.A1(new_n245), .A2(new_n234), .A3(new_n248), .A4(new_n241), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n245), .A3(new_n248), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n248), .A3(new_n241), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT81), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n243), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT5), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n247), .A2(new_n248), .ZN(new_n261));
  INV_X1    g060(.A(new_n253), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n217), .A2(new_n242), .A3(new_n218), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n258), .A3(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n249), .A2(new_n250), .A3(new_n264), .ZN(new_n268));
  OAI211_X1 g067(.A(KEYINPUT5), .B(new_n263), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT0), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G57gat), .ZN(new_n273));
  INV_X1    g072(.A(G85gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n275), .A3(new_n269), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n281));
  INV_X1    g080(.A(new_n267), .ZN(new_n282));
  INV_X1    g081(.A(new_n268), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n258), .A2(new_n257), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n285), .B(new_n243), .C1(new_n251), .C2(new_n255), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT6), .B(new_n276), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n290), .A2(KEYINPUT91), .ZN(new_n291));
  OR3_X1    g090(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(KEYINPUT91), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n294), .A2(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(KEYINPUT92), .B2(new_n294), .ZN(new_n296));
  XOR2_X1   g095(.A(G43gat), .B(G50gat), .Z(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(KEYINPUT90), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(KEYINPUT90), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n298), .A2(KEYINPUT15), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT93), .B(KEYINPUT15), .Z(new_n302));
  AOI22_X1  g101(.A1(new_n297), .A2(new_n302), .B1(G29gat), .B2(G36gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n292), .A2(new_n290), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT17), .ZN(new_n308));
  XNOR2_X1  g107(.A(G15gat), .B(G22gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT16), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(G1gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n311), .B(new_n312), .C1(G1gat), .C2(new_n309), .ZN(new_n313));
  NOR2_X1   g112(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n301), .A2(new_n306), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n308), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n307), .A2(new_n315), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G229gat), .A2(G233gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT18), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n316), .B(new_n315), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n322), .B(KEYINPUT13), .Z(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n322), .A3(new_n320), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT18), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G141gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT11), .ZN(new_n333));
  INV_X1    g132(.A(G169gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(G197gat), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT89), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(KEYINPUT89), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n337), .A2(KEYINPUT12), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT12), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n331), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n339), .A2(new_n340), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n323), .A2(new_n342), .A3(new_n327), .A4(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G15gat), .B(G43gat), .Z(new_n346));
  XNOR2_X1  g145(.A(G71gat), .B(G99gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT67), .B(G190gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n353));
  NAND2_X1  g152(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n356), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n357), .A2(KEYINPUT26), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(KEYINPUT26), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n352), .B2(new_n353), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n355), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G183gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(KEYINPUT24), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n334), .A2(new_n356), .B1(new_n373), .B2(KEYINPUT65), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT65), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT23), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n374), .A2(new_n376), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n378));
  INV_X1    g177(.A(new_n357), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(KEYINPUT23), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n373), .A2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n334), .A2(KEYINPUT64), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT64), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G169gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n373), .A2(KEYINPUT65), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n357), .A2(new_n376), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n389), .A3(new_n359), .ZN(new_n390));
  NOR2_X1   g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n368), .B2(new_n370), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n378), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT66), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT66), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(new_n378), .C1(new_n390), .C2(new_n392), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n382), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT68), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n365), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g198(.A(KEYINPUT68), .B(new_n382), .C1(new_n394), .C2(new_n396), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n242), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT74), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n403), .B(new_n242), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  INV_X1    g203(.A(new_n392), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n377), .A3(new_n387), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n395), .B1(new_n406), .B2(new_n378), .ZN(new_n407));
  INV_X1    g206(.A(new_n396), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n381), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n364), .B1(new_n409), .B2(KEYINPUT68), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n397), .A2(new_n398), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n247), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n404), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n349), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT32), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(new_n413), .B2(new_n415), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  AOI221_X4 g221(.A(new_n419), .B1(KEYINPUT33), .B2(new_n348), .C1(new_n413), .C2(new_n415), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n413), .B2(new_n415), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n399), .A2(new_n400), .A3(new_n242), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(KEYINPUT74), .B2(new_n401), .ZN(new_n428));
  INV_X1    g227(.A(new_n425), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n414), .A3(new_n404), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n422), .A2(new_n424), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT33), .B1(new_n413), .B2(new_n415), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n420), .A2(new_n434), .A3(new_n349), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n423), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n431), .A2(KEYINPUT76), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n426), .A2(new_n430), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n433), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT36), .ZN(new_n442));
  XNOR2_X1  g241(.A(G78gat), .B(G106gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT31), .ZN(new_n444));
  INV_X1    g243(.A(G50gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G197gat), .B(G204gat), .ZN(new_n447));
  AND2_X1   g246(.A1(G211gat), .A2(G218gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n447), .B1(KEYINPUT22), .B2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G211gat), .B(G218gat), .Z(new_n450));
  AND2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n449), .A2(new_n450), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT29), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT3), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n214), .B2(new_n216), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n449), .B(new_n450), .ZN(new_n459));
  OAI22_X1  g258(.A1(new_n457), .A2(new_n248), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G228gat), .ZN(new_n461));
  INV_X1    g260(.A(G233gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT82), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT3), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  OAI221_X1 g266(.A(new_n463), .B1(new_n248), .B2(new_n467), .C1(new_n458), .C2(new_n459), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n446), .B1(new_n469), .B2(G22gat), .ZN(new_n470));
  INV_X1    g269(.A(G22gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n465), .A2(new_n474), .A3(new_n471), .A4(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n470), .A2(new_n473), .A3(KEYINPUT85), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n469), .A2(G22gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n478), .A2(new_n479), .B1(new_n481), .B2(new_n446), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n410), .A2(KEYINPUT78), .A3(new_n411), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n399), .B2(new_n400), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n485), .A3(new_n466), .ZN(new_n486));
  NAND2_X1  g285(.A1(G226gat), .A2(G233gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT77), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n397), .A2(new_n364), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n489), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n453), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n489), .B1(new_n491), .B2(KEYINPUT29), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n459), .A3(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G64gat), .ZN(new_n498));
  INV_X1    g297(.A(G92gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n493), .A2(KEYINPUT30), .A3(new_n496), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n492), .B1(new_n486), .B2(new_n489), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n496), .B1(new_n502), .B2(new_n459), .ZN(new_n503));
  INV_X1    g302(.A(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n496), .B(new_n500), .C1(new_n502), .C2(new_n459), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n482), .B1(new_n509), .B2(new_n289), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n432), .B1(new_n422), .B2(new_n424), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n433), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n442), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n442), .A2(new_n514), .A3(KEYINPUT86), .A4(new_n510), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n503), .A2(KEYINPUT37), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n504), .B1(new_n503), .B2(KEYINPUT37), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT38), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n493), .A2(new_n522), .A3(new_n496), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n494), .A2(new_n453), .A3(new_n495), .ZN(new_n524));
  OAI211_X1 g323(.A(KEYINPUT37), .B(new_n524), .C1(new_n502), .C2(new_n453), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .A4(new_n504), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n287), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n270), .A2(KEYINPUT88), .A3(KEYINPUT6), .A4(new_n276), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n280), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n506), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n521), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n255), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT81), .B1(new_n252), .B2(new_n254), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n266), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT39), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n260), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n261), .A2(new_n262), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n540), .B2(new_n258), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n256), .B2(new_n258), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n542), .A3(new_n275), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT40), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n277), .ZN(new_n546));
  OR3_X1    g345(.A1(new_n543), .A2(KEYINPUT87), .A3(new_n544), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT87), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n482), .B1(new_n509), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n517), .A2(new_n518), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n482), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n437), .B(new_n439), .C1(new_n435), .C2(new_n423), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n433), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n501), .A2(new_n505), .A3(new_n508), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n288), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT35), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n435), .A2(new_n423), .A3(new_n431), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n559), .A2(new_n511), .A3(new_n482), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n531), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n509), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n345), .B1(new_n552), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n274), .B2(new_n499), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G99gat), .B(G106gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n308), .A2(new_n318), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n574), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n573), .B(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n316), .A2(new_n578), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G134gat), .B(G162gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n583), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n591), .A2(KEYINPUT95), .ZN(new_n592));
  XOR2_X1   g391(.A(G57gat), .B(G64gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(KEYINPUT95), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G71gat), .B(G78gat), .Z(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n590), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n575), .A2(new_n599), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n604), .A3(new_n602), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n578), .A2(new_n600), .A3(KEYINPUT100), .A4(KEYINPUT10), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n601), .A2(new_n604), .ZN(new_n612));
  INV_X1    g411(.A(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G176gat), .ZN(new_n616));
  INV_X1    g415(.A(G204gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n607), .A2(KEYINPUT101), .A3(new_n608), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n611), .A2(new_n614), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n609), .A2(new_n614), .ZN(new_n621));
  INV_X1    g420(.A(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(KEYINPUT102), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT21), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n315), .B1(new_n629), .B2(new_n599), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G183gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n599), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT97), .B(G211gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT98), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n635), .B(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n589), .A2(new_n628), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT103), .B1(new_n566), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n509), .A2(new_n289), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n646), .A2(new_n553), .A3(new_n433), .A4(new_n554), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n647), .A2(KEYINPUT35), .B1(new_n560), .B2(new_n563), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n534), .A2(new_n550), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n515), .B2(new_n516), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n650), .B2(new_n518), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652));
  INV_X1    g451(.A(new_n644), .ZN(new_n653));
  NOR4_X1   g452(.A1(new_n651), .A2(new_n652), .A3(new_n345), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n289), .B1(new_n645), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT16), .B(G8gat), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n509), .B(new_n659), .C1(new_n645), .C2(new_n654), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n552), .A2(new_n565), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n344), .A3(new_n644), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n652), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n566), .A2(KEYINPUT103), .A3(new_n644), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n556), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n667), .A2(KEYINPUT104), .A3(KEYINPUT42), .A4(new_n659), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n509), .B1(new_n645), .B2(new_n654), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n661), .B1(new_n669), .B2(G8gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n660), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n662), .B(new_n668), .C1(new_n670), .C2(new_n671), .ZN(G1325gat));
  NOR2_X1   g471(.A1(new_n645), .A2(new_n654), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n442), .A2(new_n514), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G15gat), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n512), .A2(new_n433), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n673), .B2(new_n678), .ZN(G1326gat));
  OAI21_X1  g478(.A(new_n482), .B1(new_n645), .B2(new_n654), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT105), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n680), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(new_n643), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n628), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n588), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n688), .A2(G29gat), .A3(new_n288), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n566), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n686), .A2(new_n345), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n551), .A2(new_n510), .A3(new_n442), .A4(new_n514), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n588), .B1(new_n565), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n589), .A2(KEYINPUT44), .ZN(new_n695));
  OAI221_X1 g494(.A(new_n692), .B1(new_n694), .B2(KEYINPUT44), .C1(new_n651), .C2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n288), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n691), .A2(new_n697), .ZN(G1328gat));
  OAI21_X1  g497(.A(G36gat), .B1(new_n696), .B2(new_n556), .ZN(new_n699));
  INV_X1    g498(.A(new_n566), .ZN(new_n700));
  NOR4_X1   g499(.A1(new_n700), .A2(G36gat), .A3(new_n556), .A4(new_n688), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(G1329gat));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n696), .B2(new_n675), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n695), .B1(new_n552), .B2(new_n565), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n565), .A2(new_n693), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT44), .B1(new_n707), .B2(new_n589), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n674), .A4(new_n692), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n705), .A2(G43gat), .A3(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n688), .A2(G43gat), .A3(new_n677), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n566), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT47), .ZN(new_n715));
  OAI21_X1  g514(.A(G43gat), .B1(new_n696), .B2(new_n675), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(new_n714), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n712), .A2(new_n715), .B1(new_n717), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g517(.A1(new_n566), .A2(new_n445), .A3(new_n482), .A4(new_n687), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n696), .A2(new_n553), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(new_n445), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g522(.A(KEYINPUT48), .B(new_n719), .C1(new_n720), .C2(new_n445), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1331gat));
  INV_X1    g524(.A(new_n628), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n589), .A2(new_n726), .A3(new_n643), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n345), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n288), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT107), .B(G57gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1332gat));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n556), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  AND2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n732), .B2(new_n733), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n728), .A2(new_n737), .A3(new_n675), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT108), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n728), .B2(new_n677), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT50), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(new_n743), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1334gat));
  NOR2_X1   g544(.A1(new_n728), .A2(new_n553), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g546(.A1(new_n344), .A2(new_n684), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n628), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n706), .A2(new_n708), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n288), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n707), .A2(new_n589), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT51), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n694), .A2(new_n754), .A3(new_n748), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n628), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n274), .A3(new_n289), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n757), .ZN(G1336gat));
  NOR2_X1   g557(.A1(new_n556), .A2(G92gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR4_X1   g559(.A1(new_n706), .A2(new_n708), .A3(new_n556), .A4(new_n749), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n499), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n760), .B(new_n764), .C1(new_n499), .C2(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1337gat));
  INV_X1    g565(.A(new_n677), .ZN(new_n767));
  AOI21_X1  g566(.A(G99gat), .B1(new_n756), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n750), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n674), .A2(G99gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(G1338gat));
  OAI21_X1  g570(.A(G106gat), .B1(new_n750), .B2(new_n553), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n553), .A2(G106gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n753), .A2(new_n628), .A3(new_n755), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n776));
  NAND4_X1  g575(.A1(new_n772), .A2(new_n773), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NOR4_X1   g576(.A1(new_n706), .A2(new_n708), .A3(new_n553), .A4(new_n749), .ZN(new_n778));
  INV_X1    g577(.A(G106gat), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n775), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n777), .A2(new_n781), .A3(new_n783), .ZN(G1339gat));
  NAND4_X1  g583(.A1(new_n603), .A2(new_n605), .A3(new_n613), .A4(new_n606), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(KEYINPUT54), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n611), .A2(new_n786), .A3(new_n619), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n607), .A2(new_n608), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n618), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT55), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n790), .A3(KEYINPUT55), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n620), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(KEYINPUT111), .A3(new_n620), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n344), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n321), .A2(new_n322), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n324), .A2(new_n326), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n324), .A2(KEYINPUT112), .A3(new_n326), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n336), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n628), .A2(new_n343), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n589), .B1(new_n797), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n804), .A2(new_n343), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n589), .A2(new_n795), .A3(new_n807), .A4(new_n796), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n643), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n644), .A2(new_n345), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n288), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n555), .A2(new_n509), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n344), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n810), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n560), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n509), .A2(new_n288), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT113), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n345), .A2(new_n226), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n814), .B1(new_n819), .B2(new_n820), .ZN(G1340gat));
  AOI21_X1  g620(.A(G120gat), .B1(new_n813), .B2(new_n628), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n726), .A2(new_n227), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n819), .B2(new_n823), .ZN(G1341gat));
  NAND3_X1  g623(.A1(new_n813), .A2(new_n219), .A3(new_n684), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n819), .A2(new_n684), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n219), .ZN(G1342gat));
  NAND2_X1  g626(.A1(new_n819), .A2(new_n589), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G134gat), .ZN(new_n829));
  INV_X1    g628(.A(new_n221), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n830), .A3(new_n589), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT56), .Z(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1343gat));
  NOR3_X1   g632(.A1(new_n674), .A2(new_n288), .A3(new_n509), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT57), .B1(new_n815), .B2(new_n482), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n793), .B2(new_n791), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n787), .A2(new_n790), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(KEYINPUT114), .A3(new_n620), .A4(new_n792), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n344), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n589), .B1(new_n843), .B2(new_n805), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n643), .B1(new_n844), .B2(new_n808), .ZN(new_n845));
  AOI211_X1 g644(.A(new_n836), .B(new_n553), .C1(new_n845), .C2(new_n810), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n834), .B1(new_n835), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G141gat), .B1(new_n847), .B2(new_n345), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n674), .A2(new_n553), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n811), .A2(new_n556), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n345), .A2(G141gat), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT115), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT58), .ZN(G1344gat));
  OR3_X1    g654(.A1(new_n850), .A2(G148gat), .A3(new_n726), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n845), .A2(new_n810), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT116), .B(new_n836), .C1(new_n858), .C2(new_n553), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n553), .B1(new_n845), .B2(new_n810), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(KEYINPUT57), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n815), .A2(KEYINPUT57), .A3(new_n482), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n628), .A3(new_n834), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n857), .B1(new_n865), .B2(G148gat), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n628), .B(new_n834), .C1(new_n835), .C2(new_n846), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n867), .A2(new_n857), .A3(G148gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n856), .B1(new_n866), .B2(new_n868), .ZN(G1345gat));
  NOR2_X1   g668(.A1(new_n643), .A2(new_n205), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT117), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n847), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n205), .B1(new_n850), .B2(new_n643), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n847), .B2(new_n588), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n206), .A3(new_n589), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT118), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n509), .A2(new_n288), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT120), .Z(new_n880));
  NAND2_X1  g679(.A1(new_n816), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881), .B2(new_n345), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n555), .A2(new_n556), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT119), .Z(new_n884));
  AOI21_X1  g683(.A(new_n289), .B1(new_n809), .B2(new_n810), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(new_n344), .A3(new_n384), .A4(new_n386), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n882), .A2(new_n887), .ZN(G1348gat));
  OAI21_X1  g687(.A(G176gat), .B1(new_n881), .B2(new_n726), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n356), .A3(new_n628), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1349gat));
  OAI21_X1  g690(.A(G183gat), .B1(new_n881), .B2(new_n643), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT122), .B1(new_n893), .B2(KEYINPUT60), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n886), .A2(new_n351), .A3(new_n684), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n892), .A2(new_n897), .A3(new_n895), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(new_n894), .ZN(G1350gat));
  NAND4_X1  g698(.A1(new_n815), .A2(new_n560), .A3(new_n589), .A4(new_n880), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G190gat), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT61), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(KEYINPUT61), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n901), .B2(KEYINPUT61), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n903), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n350), .A3(new_n589), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1351gat));
  AND2_X1   g710(.A1(new_n880), .A2(new_n675), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n864), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G197gat), .B1(new_n913), .B2(new_n345), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n885), .A2(new_n509), .A3(new_n849), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(G197gat), .A3(new_n345), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT125), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(G1352gat));
  NOR2_X1   g717(.A1(new_n726), .A2(G204gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n885), .A2(new_n509), .A3(new_n849), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT62), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(KEYINPUT126), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(KEYINPUT126), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n920), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT127), .B1(new_n920), .B2(KEYINPUT62), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n922), .A2(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n864), .A2(new_n628), .A3(new_n912), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n617), .B2(new_n927), .ZN(G1353gat));
  OR3_X1    g727(.A1(new_n915), .A2(G211gat), .A3(new_n643), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n864), .A2(new_n684), .A3(new_n912), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n913), .A2(new_n934), .A3(new_n588), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n915), .A2(new_n588), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(G1355gat));
endmodule


