

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597;

  XNOR2_X1 U326 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U327 ( .A(n443), .B(n383), .ZN(n384) );
  XOR2_X1 U328 ( .A(n491), .B(KEYINPUT101), .Z(n294) );
  XOR2_X1 U329 ( .A(KEYINPUT91), .B(KEYINPUT3), .Z(n295) );
  XOR2_X1 U330 ( .A(n333), .B(n332), .Z(n296) );
  XOR2_X1 U331 ( .A(KEYINPUT100), .B(n422), .Z(n297) );
  XOR2_X1 U332 ( .A(n481), .B(n480), .Z(n298) );
  XNOR2_X1 U333 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n467) );
  XNOR2_X1 U334 ( .A(n468), .B(n467), .ZN(n470) );
  INV_X1 U335 ( .A(KEYINPUT20), .ZN(n396) );
  XNOR2_X1 U336 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U337 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U338 ( .A(n334), .B(n296), .ZN(n335) );
  XNOR2_X1 U339 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U340 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U341 ( .A(n407), .B(n406), .ZN(n409) );
  XNOR2_X1 U342 ( .A(n414), .B(n413), .ZN(n582) );
  NOR2_X1 U343 ( .A1(n535), .A2(n485), .ZN(n570) );
  INV_X1 U344 ( .A(G183GAT), .ZN(n486) );
  XOR2_X1 U345 ( .A(KEYINPUT110), .B(n511), .Z(n517) );
  XOR2_X1 U346 ( .A(n377), .B(n376), .Z(n525) );
  XNOR2_X1 U347 ( .A(n486), .B(KEYINPUT124), .ZN(n487) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n465) );
  XNOR2_X1 U349 ( .A(n488), .B(n487), .ZN(G1350GAT) );
  XNOR2_X1 U350 ( .A(n466), .B(n465), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(G43GAT), .B(G29GAT), .Z(n300) );
  XNOR2_X1 U352 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U354 ( .A(n301), .B(KEYINPUT70), .Z(n303) );
  XNOR2_X1 U355 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n459) );
  XOR2_X1 U357 ( .A(G197GAT), .B(G8GAT), .Z(n373) );
  XOR2_X1 U358 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n305) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n373), .B(n306), .ZN(n316) );
  XOR2_X1 U362 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n308) );
  XOR2_X1 U363 ( .A(G141GAT), .B(G22GAT), .Z(n380) );
  XOR2_X1 U364 ( .A(KEYINPUT71), .B(G1GAT), .Z(n438) );
  XNOR2_X1 U365 ( .A(n380), .B(n438), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U367 ( .A(n309), .B(G113GAT), .Z(n314) );
  XOR2_X1 U368 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n311) );
  XNOR2_X1 U369 ( .A(KEYINPUT69), .B(G15GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(n312), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U374 ( .A(n459), .B(n317), .Z(n554) );
  XOR2_X1 U375 ( .A(KEYINPUT73), .B(n554), .Z(n566) );
  XOR2_X1 U376 ( .A(G148GAT), .B(KEYINPUT75), .Z(n319) );
  XNOR2_X1 U377 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n338) );
  XOR2_X1 U379 ( .A(G120GAT), .B(G71GAT), .Z(n399) );
  XOR2_X1 U380 ( .A(G64GAT), .B(G92GAT), .Z(n321) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n323) );
  INV_X1 U383 ( .A(n323), .ZN(n322) );
  NAND2_X1 U384 ( .A1(n399), .A2(n322), .ZN(n326) );
  INV_X1 U385 ( .A(n399), .ZN(n324) );
  NAND2_X1 U386 ( .A1(n324), .A2(n323), .ZN(n325) );
  NAND2_X1 U387 ( .A1(n326), .A2(n325), .ZN(n328) );
  NAND2_X1 U388 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n336) );
  XOR2_X1 U390 ( .A(G85GAT), .B(G106GAT), .Z(n330) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(KEYINPUT76), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n447) );
  XNOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n331), .B(KEYINPUT74), .ZN(n430) );
  XNOR2_X1 U395 ( .A(n447), .B(n430), .ZN(n334) );
  XOR2_X1 U396 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n333) );
  XNOR2_X1 U397 ( .A(G78GAT), .B(KEYINPUT33), .ZN(n332) );
  XOR2_X1 U398 ( .A(n338), .B(n337), .Z(n474) );
  INV_X1 U399 ( .A(n474), .ZN(n588) );
  NAND2_X1 U400 ( .A1(n566), .A2(n588), .ZN(n492) );
  XOR2_X1 U401 ( .A(G57GAT), .B(G85GAT), .Z(n340) );
  XNOR2_X1 U402 ( .A(G134GAT), .B(G120GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U404 ( .A(G155GAT), .B(G127GAT), .Z(n342) );
  XNOR2_X1 U405 ( .A(G141GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U407 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U408 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n346) );
  NAND2_X1 U409 ( .A1(G225GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U411 ( .A(KEYINPUT93), .B(n347), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n358) );
  XOR2_X1 U413 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n351) );
  XNOR2_X1 U414 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n356) );
  XNOR2_X1 U416 ( .A(G148GAT), .B(KEYINPUT2), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n295), .B(n352), .ZN(n385) );
  XOR2_X1 U418 ( .A(n385), .B(G162GAT), .Z(n354) );
  XOR2_X1 U419 ( .A(G113GAT), .B(KEYINPUT0), .Z(n401) );
  XNOR2_X1 U420 ( .A(G29GAT), .B(n401), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U422 ( .A(n356), .B(n355), .Z(n357) );
  XOR2_X1 U423 ( .A(n358), .B(n357), .Z(n581) );
  XOR2_X1 U424 ( .A(KEYINPUT19), .B(G176GAT), .Z(n360) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U427 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n361) );
  XOR2_X1 U428 ( .A(n362), .B(n361), .Z(n408) );
  INV_X1 U429 ( .A(n408), .ZN(n377) );
  XOR2_X1 U430 ( .A(KEYINPUT82), .B(G92GAT), .Z(n444) );
  XOR2_X1 U431 ( .A(G183GAT), .B(G64GAT), .Z(n429) );
  XOR2_X1 U432 ( .A(n444), .B(n429), .Z(n364) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U435 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n366) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(G190GAT), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U438 ( .A(n368), .B(n367), .Z(n375) );
  XOR2_X1 U439 ( .A(KEYINPUT90), .B(G218GAT), .Z(n370) );
  XNOR2_X1 U440 ( .A(G211GAT), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U442 ( .A(KEYINPUT21), .B(n371), .Z(n393) );
  INV_X1 U443 ( .A(n393), .ZN(n372) );
  XOR2_X1 U444 ( .A(n373), .B(n372), .Z(n374) );
  XNOR2_X1 U445 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U446 ( .A(KEYINPUT27), .B(n525), .Z(n415) );
  NOR2_X1 U447 ( .A1(n581), .A2(n415), .ZN(n550) );
  XOR2_X1 U448 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n379) );
  XNOR2_X1 U449 ( .A(KEYINPUT24), .B(KEYINPUT89), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n391) );
  XOR2_X1 U451 ( .A(G78GAT), .B(G155GAT), .Z(n425) );
  XOR2_X1 U452 ( .A(KEYINPUT22), .B(n425), .Z(n382) );
  XNOR2_X1 U453 ( .A(G197GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U454 ( .A(n382), .B(n381), .ZN(n387) );
  XOR2_X1 U455 ( .A(KEYINPUT79), .B(G162GAT), .Z(n443) );
  AND2_X1 U456 ( .A1(G228GAT), .A2(G233GAT), .ZN(n383) );
  XOR2_X1 U457 ( .A(n387), .B(n386), .Z(n389) );
  XNOR2_X1 U458 ( .A(G50GAT), .B(G106GAT), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U460 ( .A(n391), .B(n390), .Z(n392) );
  XOR2_X1 U461 ( .A(n393), .B(n392), .Z(n482) );
  XOR2_X1 U462 ( .A(n482), .B(KEYINPUT28), .Z(n394) );
  XOR2_X1 U463 ( .A(KEYINPUT65), .B(n394), .Z(n529) );
  INV_X1 U464 ( .A(n529), .ZN(n395) );
  NAND2_X1 U465 ( .A1(n550), .A2(n395), .ZN(n534) );
  NAND2_X1 U466 ( .A1(G227GAT), .A2(G233GAT), .ZN(n397) );
  XOR2_X1 U467 ( .A(G190GAT), .B(G134GAT), .Z(n455) );
  XOR2_X1 U468 ( .A(n400), .B(n455), .Z(n407) );
  XOR2_X1 U469 ( .A(G15GAT), .B(G127GAT), .Z(n426) );
  XNOR2_X1 U470 ( .A(n426), .B(n401), .ZN(n405) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(G183GAT), .Z(n403) );
  XNOR2_X1 U472 ( .A(G43GAT), .B(G99GAT), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U474 ( .A(n409), .B(n408), .Z(n535) );
  INV_X1 U475 ( .A(n535), .ZN(n527) );
  XNOR2_X1 U476 ( .A(KEYINPUT88), .B(n527), .ZN(n410) );
  NOR2_X1 U477 ( .A1(n534), .A2(n410), .ZN(n421) );
  INV_X1 U478 ( .A(n581), .ZN(n522) );
  NAND2_X1 U479 ( .A1(n527), .A2(n525), .ZN(n411) );
  NAND2_X1 U480 ( .A1(n482), .A2(n411), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n412), .B(KEYINPUT25), .ZN(n417) );
  OR2_X1 U482 ( .A1(n482), .A2(n527), .ZN(n414) );
  XOR2_X1 U483 ( .A(KEYINPUT98), .B(KEYINPUT26), .Z(n413) );
  INV_X1 U484 ( .A(n582), .ZN(n553) );
  NOR2_X1 U485 ( .A1(n415), .A2(n553), .ZN(n416) );
  OR2_X1 U486 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U487 ( .A(KEYINPUT99), .B(n418), .ZN(n419) );
  NOR2_X1 U488 ( .A1(n522), .A2(n419), .ZN(n420) );
  NOR2_X1 U489 ( .A1(n421), .A2(n420), .ZN(n422) );
  XOR2_X1 U490 ( .A(KEYINPUT85), .B(KEYINPUT12), .Z(n424) );
  XNOR2_X1 U491 ( .A(G22GAT), .B(G71GAT), .ZN(n423) );
  XNOR2_X1 U492 ( .A(n424), .B(n423), .ZN(n442) );
  XOR2_X1 U493 ( .A(n425), .B(G211GAT), .Z(n428) );
  XNOR2_X1 U494 ( .A(G8GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n434) );
  XOR2_X1 U496 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U497 ( .A1(G231GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U499 ( .A(n434), .B(n433), .Z(n440) );
  XOR2_X1 U500 ( .A(KEYINPUT14), .B(KEYINPUT83), .Z(n436) );
  XNOR2_X1 U501 ( .A(KEYINPUT15), .B(KEYINPUT84), .ZN(n435) );
  XNOR2_X1 U502 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U505 ( .A(n442), .B(n441), .Z(n560) );
  INV_X1 U506 ( .A(n560), .ZN(n591) );
  NAND2_X1 U507 ( .A1(n297), .A2(n591), .ZN(n460) );
  XOR2_X1 U508 ( .A(KEYINPUT9), .B(n443), .Z(n446) );
  XNOR2_X1 U509 ( .A(G218GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n451) );
  XOR2_X1 U511 ( .A(KEYINPUT11), .B(n447), .Z(n449) );
  NAND2_X1 U512 ( .A1(G232GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U514 ( .A(n451), .B(n450), .Z(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT10), .B(KEYINPUT81), .Z(n453) );
  XNOR2_X1 U516 ( .A(KEYINPUT80), .B(KEYINPUT64), .ZN(n452) );
  XNOR2_X1 U517 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U518 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n564) );
  XOR2_X1 U521 ( .A(KEYINPUT36), .B(n564), .Z(n594) );
  NOR2_X1 U522 ( .A1(n460), .A2(n594), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n461), .B(KEYINPUT37), .ZN(n521) );
  NOR2_X1 U524 ( .A1(n492), .A2(n521), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n462), .B(KEYINPUT38), .ZN(n508) );
  NAND2_X1 U526 ( .A1(n508), .A2(n525), .ZN(n464) );
  XNOR2_X1 U527 ( .A(G36GAT), .B(KEYINPUT108), .ZN(n463) );
  XNOR2_X1 U528 ( .A(n464), .B(n463), .ZN(G1329GAT) );
  NAND2_X1 U529 ( .A1(n508), .A2(n527), .ZN(n466) );
  XOR2_X1 U530 ( .A(KEYINPUT41), .B(n474), .Z(n569) );
  NAND2_X1 U531 ( .A1(n569), .A2(n554), .ZN(n468) );
  INV_X1 U532 ( .A(n564), .ZN(n578) );
  XOR2_X1 U533 ( .A(KEYINPUT114), .B(n560), .Z(n543) );
  NAND2_X1 U534 ( .A1(n578), .A2(n543), .ZN(n469) );
  NOR2_X1 U535 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n471), .B(KEYINPUT47), .ZN(n478) );
  NOR2_X1 U537 ( .A1(n594), .A2(n591), .ZN(n472) );
  XOR2_X1 U538 ( .A(KEYINPUT45), .B(n472), .Z(n473) );
  NOR2_X1 U539 ( .A1(n474), .A2(n473), .ZN(n476) );
  INV_X1 U540 ( .A(n566), .ZN(n475) );
  NAND2_X1 U541 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U542 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U543 ( .A(KEYINPUT48), .B(n479), .ZN(n551) );
  AND2_X1 U544 ( .A1(n551), .A2(n525), .ZN(n481) );
  XNOR2_X1 U545 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n480) );
  AND2_X1 U546 ( .A1(n482), .A2(n581), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n298), .A2(n483), .ZN(n484) );
  XOR2_X1 U548 ( .A(KEYINPUT55), .B(n484), .Z(n485) );
  INV_X1 U549 ( .A(n570), .ZN(n577) );
  NOR2_X1 U550 ( .A1(n577), .A2(n543), .ZN(n488) );
  NOR2_X1 U551 ( .A1(n564), .A2(n591), .ZN(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(n489), .ZN(n490) );
  NAND2_X1 U553 ( .A1(n490), .A2(n297), .ZN(n491) );
  NOR2_X1 U554 ( .A1(n492), .A2(n294), .ZN(n501) );
  NAND2_X1 U555 ( .A1(n522), .A2(n501), .ZN(n496) );
  XOR2_X1 U556 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n494) );
  XNOR2_X1 U557 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U560 ( .A1(n525), .A2(n501), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U563 ( .A1(n501), .A2(n527), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(n500), .ZN(G1326GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n503) );
  NAND2_X1 U567 ( .A1(n501), .A2(n529), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U569 ( .A(G22GAT), .B(n504), .ZN(G1327GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n522), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NAND2_X1 U574 ( .A1(n508), .A2(n529), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n513) );
  INV_X1 U577 ( .A(n554), .ZN(n584) );
  NAND2_X1 U578 ( .A1(n584), .A2(n569), .ZN(n510) );
  XOR2_X1 U579 ( .A(n510), .B(KEYINPUT109), .Z(n520) );
  OR2_X1 U580 ( .A1(n294), .A2(n520), .ZN(n511) );
  NAND2_X1 U581 ( .A1(n522), .A2(n517), .ZN(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U583 ( .A(G64GAT), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U584 ( .A1(n517), .A2(n525), .ZN(n514) );
  XNOR2_X1 U585 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U586 ( .A1(n517), .A2(n527), .ZN(n516) );
  XNOR2_X1 U587 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U589 ( .A1(n529), .A2(n517), .ZN(n518) );
  XNOR2_X1 U590 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U591 ( .A1(n521), .A2(n520), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n530), .A2(n522), .ZN(n523) );
  XNOR2_X1 U593 ( .A(KEYINPUT112), .B(n523), .ZN(n524) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n532) );
  NAND2_X1 U600 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U604 ( .A1(n536), .A2(n551), .ZN(n537) );
  XNOR2_X1 U605 ( .A(KEYINPUT116), .B(n537), .ZN(n542) );
  INV_X1 U606 ( .A(n542), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n547), .A2(n566), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n540) );
  NAND2_X1 U610 ( .A1(n569), .A2(n547), .ZN(n539) );
  XNOR2_X1 U611 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U612 ( .A(G120GAT), .B(n541), .Z(G1341GAT) );
  XNOR2_X1 U613 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n545) );
  NOR2_X1 U614 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U615 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U616 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U618 ( .A1(n547), .A2(n564), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n563), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U625 ( .A1(n563), .A2(n569), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT119), .Z(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(KEYINPUT120), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n560), .A2(n563), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n572) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT56), .Z(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n576) );
  XNOR2_X1 U643 ( .A(G190GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n576), .B(n575), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U646 ( .A(n580), .B(n579), .Z(G1351GAT) );
  AND2_X1 U647 ( .A1(n298), .A2(n581), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n593) );
  NOR2_X1 U649 ( .A1(n584), .A2(n593), .ZN(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(n587), .ZN(G1352GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n593), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  NOR2_X1 U656 ( .A1(n591), .A2(n593), .ZN(n592) );
  XOR2_X1 U657 ( .A(G211GAT), .B(n592), .Z(G1354GAT) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X1 U659 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

