

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733;

  XOR2_X1 U367 ( .A(n464), .B(n505), .Z(n714) );
  INV_X1 U368 ( .A(G953), .ZN(n720) );
  NOR2_X1 U369 ( .A1(n688), .A2(G953), .ZN(n689) );
  XNOR2_X2 U370 ( .A(n363), .B(n356), .ZN(n596) );
  AND2_X2 U371 ( .A1(n612), .A2(n610), .ZN(n695) );
  NOR2_X2 U372 ( .A1(n543), .A2(n563), .ZN(n631) );
  NOR2_X1 U373 ( .A1(n699), .A2(n617), .ZN(n620) );
  NAND2_X1 U374 ( .A1(n695), .A2(G210), .ZN(n408) );
  AND2_X1 U375 ( .A1(G475), .A2(n610), .ZN(n611) );
  XNOR2_X1 U376 ( .A(n402), .B(n602), .ZN(n707) );
  XNOR2_X1 U377 ( .A(n514), .B(n425), .ZN(n547) );
  XNOR2_X1 U378 ( .A(n429), .B(G119), .ZN(n487) );
  XNOR2_X1 U379 ( .A(G113), .B(KEYINPUT3), .ZN(n429) );
  NOR2_X2 U380 ( .A1(n707), .A2(n719), .ZN(n609) );
  BUF_X1 U381 ( .A(n595), .Z(n345) );
  XNOR2_X2 U382 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n716) );
  INV_X1 U383 ( .A(n642), .ZN(n358) );
  XNOR2_X1 U384 ( .A(n444), .B(n443), .ZN(n550) );
  NAND2_X1 U385 ( .A1(n608), .A2(n607), .ZN(n612) );
  NOR2_X1 U386 ( .A1(n657), .A2(n521), .ZN(n523) );
  XNOR2_X1 U387 ( .A(n534), .B(KEYINPUT74), .ZN(n549) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n502) );
  NOR2_X1 U389 ( .A1(n389), .A2(n387), .ZN(n386) );
  INV_X1 U390 ( .A(n393), .ZN(n387) );
  XNOR2_X1 U391 ( .A(n489), .B(n417), .ZN(n621) );
  XNOR2_X1 U392 ( .A(n488), .B(n418), .ZN(n417) );
  AND2_X1 U393 ( .A1(n415), .A2(n357), .ZN(n371) );
  NOR2_X1 U394 ( .A1(n412), .A2(n358), .ZN(n357) );
  XOR2_X1 U395 ( .A(G122), .B(G104), .Z(n507) );
  XNOR2_X1 U396 ( .A(G143), .B(G113), .ZN(n506) );
  XNOR2_X1 U397 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n499) );
  XOR2_X1 U398 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n500) );
  XNOR2_X1 U399 ( .A(n409), .B(n350), .ZN(n564) );
  NAND2_X1 U400 ( .A1(n394), .A2(G902), .ZN(n393) );
  NAND2_X1 U401 ( .A1(n621), .A2(n394), .ZN(n388) );
  OR2_X1 U402 ( .A1(n621), .A2(n391), .ZN(n390) );
  NAND2_X1 U403 ( .A1(n490), .A2(n392), .ZN(n391) );
  INV_X1 U404 ( .A(G902), .ZN(n392) );
  INV_X1 U405 ( .A(n695), .ZN(n377) );
  XNOR2_X1 U406 ( .A(G128), .B(G119), .ZN(n463) );
  OR2_X1 U407 ( .A1(n713), .A2(KEYINPUT24), .ZN(n455) );
  XNOR2_X1 U408 ( .A(n411), .B(n410), .ZN(n456) );
  XNOR2_X1 U409 ( .A(KEYINPUT94), .B(KEYINPUT80), .ZN(n411) );
  XNOR2_X1 U410 ( .A(G110), .B(G140), .ZN(n410) );
  XNOR2_X1 U411 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n459) );
  INV_X1 U412 ( .A(G134), .ZN(n419) );
  XNOR2_X1 U413 ( .A(KEYINPUT7), .B(KEYINPUT103), .ZN(n491) );
  XOR2_X1 U414 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n492) );
  XNOR2_X1 U415 ( .A(n359), .B(KEYINPUT41), .ZN(n681) );
  AND2_X1 U416 ( .A1(n673), .A2(n665), .ZN(n359) );
  INV_X1 U417 ( .A(n567), .ZN(n367) );
  BUF_X1 U418 ( .A(n550), .Z(n362) );
  XNOR2_X1 U419 ( .A(KEYINPUT70), .B(G469), .ZN(n400) );
  NOR2_X1 U420 ( .A1(n577), .A2(n346), .ZN(n585) );
  XNOR2_X1 U421 ( .A(n467), .B(n469), .ZN(n424) );
  NAND2_X1 U422 ( .A1(n384), .A2(n382), .ZN(n381) );
  NOR2_X1 U423 ( .A1(n383), .A2(n699), .ZN(n382) );
  NOR2_X1 U424 ( .A1(n421), .A2(G472), .ZN(n383) );
  INV_X1 U425 ( .A(G137), .ZN(n481) );
  XNOR2_X1 U426 ( .A(G131), .B(G116), .ZN(n482) );
  INV_X1 U427 ( .A(n487), .ZN(n418) );
  XNOR2_X1 U428 ( .A(n413), .B(KEYINPUT72), .ZN(n412) );
  XNOR2_X1 U429 ( .A(n580), .B(KEYINPUT87), .ZN(n581) );
  XOR2_X1 U430 ( .A(KEYINPUT17), .B(KEYINPUT90), .Z(n433) );
  XOR2_X1 U431 ( .A(KEYINPUT18), .B(KEYINPUT88), .Z(n427) );
  OR2_X1 U432 ( .A1(G237), .A2(G902), .ZN(n517) );
  XNOR2_X1 U433 ( .A(G902), .B(KEYINPUT15), .ZN(n604) );
  XNOR2_X1 U434 ( .A(n423), .B(n422), .ZN(n521) );
  INV_X1 U435 ( .A(KEYINPUT69), .ZN(n422) );
  NAND2_X1 U436 ( .A1(n653), .A2(n531), .ZN(n423) );
  NAND2_X1 U437 ( .A1(n385), .A2(n390), .ZN(n528) );
  AND2_X1 U438 ( .A1(n388), .A2(n386), .ZN(n385) );
  NOR2_X1 U439 ( .A1(n645), .A2(n369), .ZN(n368) );
  INV_X1 U440 ( .A(n644), .ZN(n369) );
  INV_X1 U441 ( .A(KEYINPUT45), .ZN(n602) );
  XNOR2_X1 U442 ( .A(G110), .B(G104), .ZN(n700) );
  XNOR2_X1 U443 ( .A(n511), .B(n510), .ZN(n614) );
  XNOR2_X1 U444 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U445 ( .A(G107), .B(KEYINPUT93), .Z(n446) );
  INV_X1 U446 ( .A(G146), .ZN(n449) );
  INV_X1 U447 ( .A(KEYINPUT0), .ZN(n356) );
  XNOR2_X1 U448 ( .A(n515), .B(KEYINPUT105), .ZN(n545) );
  NAND2_X1 U449 ( .A1(n390), .A2(n349), .ZN(n657) );
  XNOR2_X1 U450 ( .A(n462), .B(n360), .ZN(n697) );
  XNOR2_X1 U451 ( .A(n461), .B(n465), .ZN(n360) );
  XNOR2_X1 U452 ( .A(n496), .B(n361), .ZN(n693) );
  XNOR2_X1 U453 ( .A(n495), .B(n497), .ZN(n361) );
  XNOR2_X1 U454 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n646) );
  XNOR2_X1 U455 ( .A(KEYINPUT115), .B(KEYINPUT42), .ZN(n526) );
  NOR2_X1 U456 ( .A1(n540), .A2(n539), .ZN(n541) );
  INV_X1 U457 ( .A(KEYINPUT35), .ZN(n570) );
  XNOR2_X1 U458 ( .A(n355), .B(n353), .ZN(n731) );
  NAND2_X1 U459 ( .A1(n585), .A2(n575), .ZN(n355) );
  XNOR2_X1 U460 ( .A(n365), .B(n364), .ZN(n729) );
  INV_X1 U461 ( .A(KEYINPUT113), .ZN(n364) );
  OR2_X1 U462 ( .A1(n549), .A2(n366), .ZN(n365) );
  XNOR2_X1 U463 ( .A(n545), .B(KEYINPUT110), .ZN(n636) );
  AND2_X1 U464 ( .A1(n375), .A2(n379), .ZN(n374) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n397) );
  NAND2_X1 U466 ( .A1(n695), .A2(G469), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n657), .B(KEYINPUT6), .ZN(n346) );
  OR2_X1 U468 ( .A1(KEYINPUT47), .A2(n553), .ZN(n347) );
  AND2_X1 U469 ( .A1(n380), .A2(n378), .ZN(n348) );
  AND2_X1 U470 ( .A1(n388), .A2(n393), .ZN(n349) );
  XOR2_X1 U471 ( .A(KEYINPUT75), .B(KEYINPUT19), .Z(n350) );
  AND2_X1 U472 ( .A1(n421), .A2(G472), .ZN(n351) );
  INV_X1 U473 ( .A(n624), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n623), .B(n622), .ZN(n624) );
  INV_X1 U475 ( .A(n665), .ZN(n389) );
  XOR2_X1 U476 ( .A(n439), .B(n438), .Z(n352) );
  XOR2_X1 U477 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n353) );
  NOR2_X1 U478 ( .A1(G952), .A2(n720), .ZN(n699) );
  INV_X1 U479 ( .A(n699), .ZN(n420) );
  XOR2_X1 U480 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n354) );
  INV_X1 U481 ( .A(n596), .ZN(n590) );
  NAND2_X1 U482 ( .A1(n596), .A2(n573), .ZN(n574) );
  NAND2_X1 U483 ( .A1(n732), .A2(n733), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n527), .B(n526), .ZN(n732) );
  XNOR2_X1 U485 ( .A(n408), .B(n352), .ZN(n407) );
  OR2_X2 U486 ( .A1(n691), .A2(G902), .ZN(n401) );
  XNOR2_X1 U487 ( .A(n451), .B(n452), .ZN(n691) );
  XNOR2_X2 U488 ( .A(n556), .B(n555), .ZN(n595) );
  XNOR2_X1 U489 ( .A(n371), .B(KEYINPUT48), .ZN(n370) );
  NAND2_X1 U490 ( .A1(n414), .A2(n347), .ZN(n413) );
  NAND2_X1 U491 ( .A1(n370), .A2(n368), .ZN(n719) );
  NAND2_X1 U492 ( .A1(n564), .A2(n565), .ZN(n363) );
  NAND2_X1 U493 ( .A1(n407), .A2(n420), .ZN(n406) );
  NAND2_X1 U494 ( .A1(n731), .A2(n630), .ZN(n582) );
  NAND2_X1 U495 ( .A1(n367), .A2(n362), .ZN(n366) );
  NAND2_X1 U496 ( .A1(n374), .A2(n372), .ZN(G57) );
  NAND2_X1 U497 ( .A1(n348), .A2(n373), .ZN(n372) );
  INV_X1 U498 ( .A(n381), .ZN(n373) );
  NAND2_X1 U499 ( .A1(n381), .A2(KEYINPUT63), .ZN(n375) );
  NAND2_X1 U500 ( .A1(n695), .A2(n351), .ZN(n384) );
  NAND2_X1 U501 ( .A1(n377), .A2(n624), .ZN(n380) );
  NAND2_X1 U502 ( .A1(n377), .A2(n376), .ZN(n379) );
  AND2_X1 U503 ( .A1(n624), .A2(KEYINPUT63), .ZN(n376) );
  INV_X1 U504 ( .A(KEYINPUT63), .ZN(n378) );
  INV_X1 U505 ( .A(n490), .ZN(n394) );
  NOR2_X2 U506 ( .A1(n682), .A2(n590), .ZN(n566) );
  XNOR2_X2 U507 ( .A(n395), .B(n557), .ZN(n682) );
  NAND2_X1 U508 ( .A1(n396), .A2(n346), .ZN(n395) );
  XNOR2_X1 U509 ( .A(n595), .B(KEYINPUT109), .ZN(n396) );
  NOR2_X1 U510 ( .A1(n397), .A2(n699), .ZN(G54) );
  XNOR2_X1 U511 ( .A(n691), .B(n690), .ZN(n398) );
  XNOR2_X2 U512 ( .A(n591), .B(KEYINPUT1), .ZN(n586) );
  XNOR2_X2 U513 ( .A(n401), .B(n400), .ZN(n591) );
  NAND2_X1 U514 ( .A1(n403), .A2(n601), .ZN(n402) );
  NAND2_X1 U515 ( .A1(n404), .A2(n584), .ZN(n403) );
  NAND2_X1 U516 ( .A1(n583), .A2(n730), .ZN(n404) );
  NAND2_X1 U517 ( .A1(n405), .A2(KEYINPUT78), .ZN(n647) );
  INV_X1 U518 ( .A(n609), .ZN(n405) );
  XNOR2_X1 U519 ( .A(n406), .B(n354), .ZN(G51) );
  INV_X1 U520 ( .A(n564), .ZN(n563) );
  NAND2_X1 U521 ( .A1(n550), .A2(n665), .ZN(n409) );
  XNOR2_X1 U522 ( .A(n552), .B(KEYINPUT79), .ZN(n414) );
  XNOR2_X1 U523 ( .A(n416), .B(n538), .ZN(n415) );
  XNOR2_X2 U524 ( .A(n718), .B(n449), .ZN(n488) );
  XNOR2_X2 U525 ( .A(n448), .B(n419), .ZN(n718) );
  XNOR2_X2 U526 ( .A(n468), .B(n424), .ZN(n653) );
  XOR2_X1 U527 ( .A(n513), .B(n512), .Z(n425) );
  XNOR2_X1 U528 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U529 ( .A(n484), .B(n483), .ZN(n486) );
  INV_X1 U530 ( .A(n453), .ZN(n434) );
  INV_X1 U531 ( .A(n604), .ZN(n603) );
  XNOR2_X1 U532 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U533 ( .A(n456), .B(KEYINPUT23), .ZN(n457) );
  XNOR2_X1 U534 ( .A(n450), .B(n435), .ZN(n436) );
  XNOR2_X1 U535 ( .A(n458), .B(n457), .ZN(n462) );
  XNOR2_X1 U536 ( .A(n647), .B(n646), .ZN(n686) );
  XNOR2_X1 U537 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U538 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U539 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U540 ( .A(n618), .B(KEYINPUT60), .ZN(n619) );
  XNOR2_X1 U541 ( .A(n620), .B(n619), .ZN(G60) );
  XOR2_X1 U542 ( .A(KEYINPUT125), .B(KEYINPUT54), .Z(n439) );
  XOR2_X2 U543 ( .A(G143), .B(G128), .Z(n448) );
  NAND2_X1 U544 ( .A1(G224), .A2(n720), .ZN(n426) );
  XNOR2_X1 U545 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U546 ( .A(n448), .B(n428), .ZN(n432) );
  XNOR2_X1 U547 ( .A(n487), .B(KEYINPUT16), .ZN(n431) );
  XOR2_X1 U548 ( .A(G116), .B(G107), .Z(n430) );
  XNOR2_X1 U549 ( .A(G122), .B(n430), .ZN(n497) );
  XNOR2_X1 U550 ( .A(n431), .B(n497), .ZN(n702) );
  XNOR2_X1 U551 ( .A(n432), .B(n702), .ZN(n437) );
  XNOR2_X1 U552 ( .A(G101), .B(n716), .ZN(n485) );
  XNOR2_X1 U553 ( .A(n485), .B(n700), .ZN(n450) );
  XNOR2_X2 U554 ( .A(G146), .B(G125), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n437), .B(n436), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n440), .B(KEYINPUT55), .ZN(n438) );
  NAND2_X1 U557 ( .A1(n440), .A2(n604), .ZN(n444) );
  XOR2_X1 U558 ( .A(KEYINPUT91), .B(KEYINPUT77), .Z(n442) );
  NAND2_X1 U559 ( .A1(G210), .A2(n517), .ZN(n441) );
  XNOR2_X1 U560 ( .A(n442), .B(n441), .ZN(n443) );
  NAND2_X1 U561 ( .A1(G227), .A2(n720), .ZN(n445) );
  XNOR2_X1 U562 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U563 ( .A(G137), .B(KEYINPUT68), .Z(n464) );
  XOR2_X1 U564 ( .A(G131), .B(G140), .Z(n505) );
  XOR2_X1 U565 ( .A(n447), .B(n714), .Z(n452) );
  XNOR2_X1 U566 ( .A(n488), .B(n450), .ZN(n451) );
  INV_X1 U567 ( .A(KEYINPUT25), .ZN(n469) );
  XNOR2_X2 U568 ( .A(n453), .B(KEYINPUT10), .ZN(n713) );
  NAND2_X1 U569 ( .A1(n713), .A2(KEYINPUT24), .ZN(n454) );
  NAND2_X1 U570 ( .A1(n455), .A2(n454), .ZN(n458) );
  NAND2_X1 U571 ( .A1(n720), .A2(G234), .ZN(n460) );
  XNOR2_X1 U572 ( .A(n460), .B(n459), .ZN(n494) );
  AND2_X1 U573 ( .A1(G221), .A2(n494), .ZN(n461) );
  NOR2_X1 U574 ( .A1(G902), .A2(n697), .ZN(n468) );
  NAND2_X1 U575 ( .A1(G234), .A2(n604), .ZN(n466) );
  XNOR2_X1 U576 ( .A(KEYINPUT20), .B(n466), .ZN(n470) );
  NAND2_X1 U577 ( .A1(n470), .A2(G217), .ZN(n467) );
  NAND2_X1 U578 ( .A1(G221), .A2(n470), .ZN(n471) );
  XNOR2_X1 U579 ( .A(n471), .B(KEYINPUT21), .ZN(n652) );
  NAND2_X1 U580 ( .A1(G234), .A2(G237), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n472), .B(KEYINPUT14), .ZN(n474) );
  NAND2_X1 U582 ( .A1(G952), .A2(n474), .ZN(n680) );
  NOR2_X1 U583 ( .A1(n680), .A2(G953), .ZN(n473) );
  XNOR2_X1 U584 ( .A(n473), .B(KEYINPUT92), .ZN(n560) );
  NAND2_X1 U585 ( .A1(G902), .A2(n474), .ZN(n558) );
  NOR2_X1 U586 ( .A1(G900), .A2(n558), .ZN(n475) );
  NAND2_X1 U587 ( .A1(G953), .A2(n475), .ZN(n476) );
  XNOR2_X1 U588 ( .A(KEYINPUT111), .B(n476), .ZN(n477) );
  NOR2_X1 U589 ( .A1(n560), .A2(n477), .ZN(n478) );
  NOR2_X1 U590 ( .A1(n652), .A2(n478), .ZN(n531) );
  XOR2_X1 U591 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n480) );
  NAND2_X1 U592 ( .A1(n502), .A2(G210), .ZN(n479) );
  XNOR2_X1 U593 ( .A(n480), .B(n479), .ZN(n484) );
  XOR2_X1 U594 ( .A(n486), .B(n485), .Z(n489) );
  XNOR2_X1 U595 ( .A(G472), .B(KEYINPUT96), .ZN(n490) );
  XNOR2_X1 U596 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U597 ( .A(n718), .B(n493), .Z(n496) );
  NAND2_X1 U598 ( .A1(G217), .A2(n494), .ZN(n495) );
  NOR2_X1 U599 ( .A1(G902), .A2(n693), .ZN(n498) );
  XNOR2_X1 U600 ( .A(G478), .B(n498), .ZN(n548) );
  XNOR2_X1 U601 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U602 ( .A(n713), .B(n501), .Z(n504) );
  NAND2_X1 U603 ( .A1(G214), .A2(n502), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n504), .B(n503), .ZN(n511) );
  XNOR2_X1 U605 ( .A(n505), .B(KEYINPUT100), .ZN(n509) );
  XNOR2_X1 U606 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U607 ( .A1(n614), .A2(G902), .ZN(n514) );
  XOR2_X1 U608 ( .A(KEYINPUT13), .B(KEYINPUT102), .Z(n513) );
  XNOR2_X1 U609 ( .A(KEYINPUT101), .B(G475), .ZN(n512) );
  INV_X1 U610 ( .A(n547), .ZN(n544) );
  NAND2_X1 U611 ( .A1(n548), .A2(n544), .ZN(n515) );
  NAND2_X1 U612 ( .A1(n346), .A2(n636), .ZN(n516) );
  NOR2_X1 U613 ( .A1(n521), .A2(n516), .ZN(n518) );
  NAND2_X1 U614 ( .A1(G214), .A2(n517), .ZN(n665) );
  NAND2_X1 U615 ( .A1(n518), .A2(n665), .ZN(n539) );
  NOR2_X1 U616 ( .A1(n586), .A2(n539), .ZN(n519) );
  XNOR2_X1 U617 ( .A(n519), .B(KEYINPUT43), .ZN(n520) );
  NOR2_X1 U618 ( .A1(n362), .A2(n520), .ZN(n645) );
  XNOR2_X1 U619 ( .A(KEYINPUT28), .B(KEYINPUT114), .ZN(n522) );
  XNOR2_X1 U620 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U621 ( .A1(n524), .A2(n591), .ZN(n543) );
  NAND2_X1 U622 ( .A1(n547), .A2(n548), .ZN(n525) );
  XNOR2_X1 U623 ( .A(n525), .B(KEYINPUT106), .ZN(n666) );
  XNOR2_X1 U624 ( .A(n362), .B(KEYINPUT38), .ZN(n668) );
  NOR2_X1 U625 ( .A1(n666), .A2(n668), .ZN(n673) );
  NOR2_X1 U626 ( .A1(n543), .A2(n681), .ZN(n527) );
  XNOR2_X1 U627 ( .A(KEYINPUT30), .B(KEYINPUT112), .ZN(n529) );
  XNOR2_X1 U628 ( .A(n529), .B(n528), .ZN(n530) );
  NOR2_X1 U629 ( .A1(n653), .A2(n530), .ZN(n533) );
  AND2_X1 U630 ( .A1(n531), .A2(n591), .ZN(n532) );
  NAND2_X1 U631 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U632 ( .A1(n549), .A2(n668), .ZN(n536) );
  XNOR2_X1 U633 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n536), .B(n535), .ZN(n554) );
  NAND2_X1 U635 ( .A1(n554), .A2(n545), .ZN(n537) );
  XNOR2_X1 U636 ( .A(n537), .B(KEYINPUT40), .ZN(n733) );
  XNOR2_X1 U637 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n538) );
  INV_X1 U638 ( .A(n362), .ZN(n540) );
  XNOR2_X1 U639 ( .A(KEYINPUT36), .B(n541), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n542), .A2(n586), .ZN(n642) );
  NOR2_X1 U641 ( .A1(n544), .A2(n548), .ZN(n638) );
  NOR2_X1 U642 ( .A1(n545), .A2(n638), .ZN(n667) );
  INV_X1 U643 ( .A(n667), .ZN(n546) );
  NAND2_X1 U644 ( .A1(n631), .A2(n546), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n553), .A2(KEYINPUT47), .ZN(n551) );
  OR2_X1 U646 ( .A1(n548), .A2(n547), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n551), .A2(n729), .ZN(n552) );
  NAND2_X1 U648 ( .A1(n554), .A2(n638), .ZN(n644) );
  NOR2_X1 U649 ( .A1(n652), .A2(n653), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n589), .A2(n586), .ZN(n556) );
  INV_X1 U651 ( .A(KEYINPUT73), .ZN(n555) );
  INV_X1 U652 ( .A(KEYINPUT33), .ZN(n557) );
  NOR2_X1 U653 ( .A1(G898), .A2(n720), .ZN(n703) );
  INV_X1 U654 ( .A(n558), .ZN(n559) );
  NAND2_X1 U655 ( .A1(n703), .A2(n559), .ZN(n562) );
  INV_X1 U656 ( .A(n560), .ZN(n561) );
  NAND2_X1 U657 ( .A1(n562), .A2(n561), .ZN(n565) );
  XNOR2_X1 U658 ( .A(n566), .B(KEYINPUT34), .ZN(n569) );
  XOR2_X1 U659 ( .A(n567), .B(KEYINPUT76), .Z(n568) );
  NAND2_X1 U660 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X2 U661 ( .A(n571), .B(n570), .ZN(n730) );
  INV_X1 U662 ( .A(n730), .ZN(n572) );
  INV_X1 U663 ( .A(KEYINPUT44), .ZN(n579) );
  NAND2_X1 U664 ( .A1(n572), .A2(n579), .ZN(n584) );
  NOR2_X1 U665 ( .A1(n652), .A2(n666), .ZN(n573) );
  XNOR2_X1 U666 ( .A(KEYINPUT22), .B(n574), .ZN(n577) );
  AND2_X1 U667 ( .A1(n586), .A2(n653), .ZN(n575) );
  NAND2_X1 U668 ( .A1(n653), .A2(n657), .ZN(n576) );
  NOR2_X1 U669 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U670 ( .A(KEYINPUT1), .B(n591), .Z(n648) );
  NAND2_X1 U671 ( .A1(n578), .A2(n648), .ZN(n630) );
  NAND2_X1 U672 ( .A1(n579), .A2(KEYINPUT86), .ZN(n580) );
  XNOR2_X1 U673 ( .A(n582), .B(n581), .ZN(n583) );
  NOR2_X1 U674 ( .A1(n586), .A2(n653), .ZN(n587) );
  NAND2_X1 U675 ( .A1(n585), .A2(n587), .ZN(n588) );
  XNOR2_X1 U676 ( .A(KEYINPUT107), .B(n588), .ZN(n727) );
  INV_X1 U677 ( .A(n589), .ZN(n649) );
  NOR2_X1 U678 ( .A1(n590), .A2(n649), .ZN(n593) );
  AND2_X1 U679 ( .A1(n657), .A2(n591), .ZN(n592) );
  NAND2_X1 U680 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U681 ( .A(KEYINPUT97), .B(n594), .ZN(n626) );
  NOR2_X1 U682 ( .A1(n657), .A2(n345), .ZN(n662) );
  NAND2_X1 U683 ( .A1(n596), .A2(n662), .ZN(n597) );
  XNOR2_X1 U684 ( .A(n597), .B(KEYINPUT31), .ZN(n639) );
  NOR2_X1 U685 ( .A1(n626), .A2(n639), .ZN(n598) );
  NOR2_X1 U686 ( .A1(n667), .A2(n598), .ZN(n599) );
  NOR2_X1 U687 ( .A1(n727), .A2(n599), .ZN(n600) );
  XNOR2_X1 U688 ( .A(KEYINPUT108), .B(n600), .ZN(n601) );
  NAND2_X1 U689 ( .A1(n609), .A2(n603), .ZN(n608) );
  XNOR2_X1 U690 ( .A(KEYINPUT83), .B(n604), .ZN(n605) );
  NAND2_X1 U691 ( .A1(n605), .A2(KEYINPUT2), .ZN(n606) );
  XNOR2_X1 U692 ( .A(KEYINPUT66), .B(n606), .ZN(n607) );
  NAND2_X1 U693 ( .A1(KEYINPUT2), .A2(n609), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n616) );
  INV_X1 U695 ( .A(KEYINPUT59), .ZN(n613) );
  INV_X1 U696 ( .A(KEYINPUT67), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT62), .ZN(n623) );
  XOR2_X1 U698 ( .A(KEYINPUT89), .B(KEYINPUT116), .Z(n622) );
  NAND2_X1 U699 ( .A1(n636), .A2(n626), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(G104), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n628) );
  NAND2_X1 U702 ( .A1(n626), .A2(n638), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U704 ( .A(G107), .B(n629), .ZN(G9) );
  XNOR2_X1 U705 ( .A(G110), .B(n630), .ZN(G12) );
  XOR2_X1 U706 ( .A(KEYINPUT118), .B(KEYINPUT29), .Z(n633) );
  NAND2_X1 U707 ( .A1(n631), .A2(n638), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U709 ( .A(G128), .B(n634), .ZN(G30) );
  NAND2_X1 U710 ( .A1(n636), .A2(n631), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(G146), .ZN(G48) );
  NAND2_X1 U712 ( .A1(n636), .A2(n639), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(G113), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(G116), .ZN(G18) );
  XOR2_X1 U716 ( .A(G125), .B(KEYINPUT37), .Z(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(G27) );
  XOR2_X1 U718 ( .A(G134), .B(KEYINPUT119), .Z(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(G36) );
  XOR2_X1 U720 ( .A(G140), .B(n645), .Z(G42) );
  XOR2_X1 U721 ( .A(KEYINPUT122), .B(KEYINPUT50), .Z(n651) );
  NAND2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(n660) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT121), .B(KEYINPUT49), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(KEYINPUT120), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U731 ( .A(KEYINPUT51), .B(n663), .Z(n664) );
  NOR2_X1 U732 ( .A1(n681), .A2(n664), .ZN(n676) );
  INV_X1 U733 ( .A(n666), .ZN(n670) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n389), .A2(n671), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n682), .A2(n674), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U740 ( .A(n677), .B(KEYINPUT123), .Z(n678) );
  XNOR2_X1 U741 ( .A(KEYINPUT52), .B(n678), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n687), .B(KEYINPUT124), .ZN(n688) );
  XNOR2_X1 U747 ( .A(n689), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U748 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n690) );
  NAND2_X1 U749 ( .A1(G478), .A2(n695), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U751 ( .A1(n699), .A2(n694), .ZN(G63) );
  NAND2_X1 U752 ( .A1(G217), .A2(n695), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U754 ( .A1(n699), .A2(n698), .ZN(G66) );
  XOR2_X1 U755 ( .A(G101), .B(n700), .Z(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n711) );
  NAND2_X1 U758 ( .A1(G953), .A2(G224), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n705), .B(KEYINPUT61), .ZN(n706) );
  NAND2_X1 U760 ( .A1(n706), .A2(G898), .ZN(n709) );
  OR2_X1 U761 ( .A1(G953), .A2(n707), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U764 ( .A(KEYINPUT126), .B(n712), .ZN(G69) );
  XNOR2_X1 U765 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(n722) );
  XNOR2_X1 U768 ( .A(n719), .B(n722), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n721), .A2(n720), .ZN(n726) );
  XNOR2_X1 U770 ( .A(G227), .B(n722), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(G953), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n726), .A2(n725), .ZN(G72) );
  XNOR2_X1 U774 ( .A(G101), .B(n727), .ZN(n728) );
  XNOR2_X1 U775 ( .A(n728), .B(KEYINPUT117), .ZN(G3) );
  XNOR2_X1 U776 ( .A(n729), .B(G143), .ZN(G45) );
  XNOR2_X1 U777 ( .A(G122), .B(n730), .ZN(G24) );
  XNOR2_X1 U778 ( .A(n731), .B(G119), .ZN(G21) );
  XNOR2_X1 U779 ( .A(G137), .B(n732), .ZN(G39) );
  XNOR2_X1 U780 ( .A(G131), .B(n733), .ZN(G33) );
endmodule

