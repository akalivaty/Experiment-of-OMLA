

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751;

  INV_X1 U372 ( .A(n726), .ZN(n352) );
  INV_X1 U373 ( .A(n726), .ZN(n356) );
  OR2_X1 U374 ( .A1(n563), .A2(KEYINPUT79), .ZN(n564) );
  XNOR2_X1 U375 ( .A(n613), .B(n572), .ZN(n686) );
  NAND2_X1 U376 ( .A1(n554), .A2(n555), .ZN(n482) );
  XNOR2_X1 U377 ( .A(n429), .B(n428), .ZN(n507) );
  XNOR2_X1 U378 ( .A(n427), .B(G101), .ZN(n429) );
  INV_X1 U379 ( .A(G104), .ZN(n427) );
  INV_X2 U380 ( .A(G953), .ZN(n517) );
  INV_X1 U381 ( .A(n351), .ZN(n370) );
  NAND2_X1 U382 ( .A1(n353), .A2(n352), .ZN(n351) );
  XNOR2_X1 U383 ( .A(n716), .B(n354), .ZN(n353) );
  INV_X1 U384 ( .A(n715), .ZN(n354) );
  INV_X1 U385 ( .A(n355), .ZN(n631) );
  NAND2_X1 U386 ( .A1(n357), .A2(n356), .ZN(n355) );
  XNOR2_X1 U387 ( .A(n627), .B(n358), .ZN(n357) );
  INV_X1 U388 ( .A(n626), .ZN(n358) );
  NAND2_X1 U389 ( .A1(n401), .A2(KEYINPUT65), .ZN(n382) );
  NAND2_X2 U390 ( .A1(n395), .A2(n624), .ZN(n401) );
  XNOR2_X2 U391 ( .A(n549), .B(KEYINPUT91), .ZN(n553) );
  XOR2_X1 U392 ( .A(G104), .B(KEYINPUT11), .Z(n462) );
  XNOR2_X1 U393 ( .A(KEYINPUT4), .B(G146), .ZN(n483) );
  INV_X1 U394 ( .A(KEYINPUT45), .ZN(n379) );
  AND2_X1 U395 ( .A1(n596), .A2(n595), .ZN(n655) );
  XNOR2_X1 U396 ( .A(KEYINPUT42), .B(n586), .ZN(n751) );
  NAND2_X2 U397 ( .A1(n366), .A2(n399), .ZN(n383) );
  AND2_X2 U398 ( .A1(n384), .A2(n400), .ZN(n366) );
  NAND2_X4 U399 ( .A1(n383), .A2(n380), .ZN(n721) );
  XNOR2_X2 U400 ( .A(n449), .B(KEYINPUT25), .ZN(n575) );
  XNOR2_X2 U401 ( .A(n525), .B(n524), .ZN(n549) );
  XNOR2_X1 U402 ( .A(n406), .B(n454), .ZN(n671) );
  XNOR2_X1 U403 ( .A(n432), .B(n431), .ZN(n496) );
  NAND2_X1 U404 ( .A1(n408), .A2(n419), .ZN(n738) );
  INV_X1 U405 ( .A(n546), .ZN(n368) );
  OR2_X1 U406 ( .A1(G237), .A2(G902), .ZN(n436) );
  XNOR2_X1 U407 ( .A(n415), .B(n365), .ZN(n408) );
  OR2_X1 U408 ( .A1(n639), .A2(G902), .ZN(n511) );
  NAND2_X1 U409 ( .A1(n359), .A2(n667), .ZN(n381) );
  NAND2_X1 U410 ( .A1(n667), .A2(n623), .ZN(n384) );
  NOR2_X1 U411 ( .A1(n608), .A2(n417), .ZN(n416) );
  AND2_X1 U412 ( .A1(n671), .A2(n363), .ZN(n577) );
  INV_X1 U413 ( .A(n702), .ZN(n405) );
  AND2_X1 U414 ( .A1(n367), .A2(n658), .ZN(n609) );
  NOR2_X1 U415 ( .A1(n368), .A2(n501), .ZN(n367) );
  INV_X1 U416 ( .A(n577), .ZN(n392) );
  INV_X1 U417 ( .A(KEYINPUT30), .ZN(n394) );
  XNOR2_X1 U418 ( .A(n677), .B(n500), .ZN(n546) );
  XNOR2_X1 U419 ( .A(n737), .B(n497), .ZN(n625) );
  OR2_X1 U420 ( .A1(n621), .A2(n620), .ZN(n624) );
  XOR2_X1 U421 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n425) );
  XOR2_X1 U422 ( .A(KEYINPUT86), .B(G125), .Z(n420) );
  XNOR2_X1 U423 ( .A(n422), .B(n421), .ZN(n387) );
  XNOR2_X1 U424 ( .A(KEYINPUT76), .B(G143), .ZN(n422) );
  INV_X1 U425 ( .A(n738), .ZN(n397) );
  NAND2_X1 U426 ( .A1(n414), .A2(n580), .ZN(n581) );
  INV_X1 U427 ( .A(KEYINPUT36), .ZN(n503) );
  NOR2_X1 U428 ( .A1(n536), .A2(n546), .ZN(n537) );
  AND2_X1 U429 ( .A1(n403), .A2(n585), .ZN(n596) );
  BUF_X1 U430 ( .A(n539), .Z(n677) );
  XNOR2_X1 U431 ( .A(n535), .B(KEYINPUT22), .ZN(n538) );
  XNOR2_X1 U432 ( .A(n373), .B(n413), .ZN(n728) );
  XNOR2_X1 U433 ( .A(n475), .B(KEYINPUT16), .ZN(n413) );
  XNOR2_X1 U434 ( .A(n507), .B(n496), .ZN(n373) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n488) );
  XNOR2_X1 U436 ( .A(n402), .B(KEYINPUT15), .ZN(n617) );
  XNOR2_X1 U437 ( .A(G902), .B(KEYINPUT84), .ZN(n402) );
  XNOR2_X1 U438 ( .A(G125), .B(KEYINPUT10), .ZN(n444) );
  XNOR2_X1 U439 ( .A(G143), .B(G122), .ZN(n463) );
  INV_X1 U440 ( .A(n617), .ZN(n620) );
  INV_X1 U441 ( .A(KEYINPUT78), .ZN(n407) );
  XNOR2_X1 U442 ( .A(n457), .B(KEYINPUT69), .ZN(n485) );
  XNOR2_X1 U443 ( .A(G131), .B(KEYINPUT70), .ZN(n457) );
  XNOR2_X1 U444 ( .A(n579), .B(KEYINPUT111), .ZN(n414) );
  INV_X1 U445 ( .A(KEYINPUT38), .ZN(n572) );
  XNOR2_X1 U446 ( .A(n481), .B(G478), .ZN(n532) );
  INV_X1 U447 ( .A(G902), .ZN(n498) );
  NAND2_X1 U448 ( .A1(n453), .A2(G221), .ZN(n406) );
  XNOR2_X1 U449 ( .A(G119), .B(KEYINPUT85), .ZN(n430) );
  XNOR2_X1 U450 ( .A(G119), .B(G137), .ZN(n438) );
  XOR2_X1 U451 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n440) );
  XOR2_X1 U452 ( .A(G116), .B(G122), .Z(n475) );
  XNOR2_X1 U453 ( .A(n387), .B(G134), .ZN(n487) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n450) );
  INV_X1 U455 ( .A(KEYINPUT34), .ZN(n385) );
  BUF_X1 U456 ( .A(n571), .Z(n613) );
  XNOR2_X1 U457 ( .A(n390), .B(n389), .ZN(n589) );
  INV_X1 U458 ( .A(KEYINPUT74), .ZN(n389) );
  NOR2_X1 U459 ( .A1(n576), .A2(n392), .ZN(n391) );
  INV_X1 U460 ( .A(n532), .ZN(n555) );
  XNOR2_X1 U461 ( .A(n632), .B(KEYINPUT59), .ZN(n633) );
  INV_X1 U462 ( .A(n401), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n728), .B(n372), .ZN(n714) );
  XNOR2_X1 U464 ( .A(n374), .B(n412), .ZN(n372) );
  AND2_X1 U465 ( .A1(n628), .A2(G953), .ZN(n726) );
  XNOR2_X1 U466 ( .A(n504), .B(n364), .ZN(n513) );
  INV_X1 U467 ( .A(KEYINPUT32), .ZN(n375) );
  OR2_X2 U468 ( .A1(n538), .A2(n377), .ZN(n376) );
  NAND2_X1 U469 ( .A1(n537), .A2(n378), .ZN(n377) );
  AND2_X1 U470 ( .A1(n410), .A2(n409), .ZN(n646) );
  INV_X1 U471 ( .A(n677), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n411), .B(KEYINPUT93), .ZN(n410) );
  AND2_X1 U473 ( .A1(n623), .A2(KEYINPUT65), .ZN(n359) );
  AND2_X1 U474 ( .A1(n419), .A2(n407), .ZN(n360) );
  INV_X1 U475 ( .A(n670), .ZN(n378) );
  XOR2_X1 U476 ( .A(n434), .B(n433), .Z(n361) );
  AND2_X1 U477 ( .A1(n673), .A2(n585), .ZN(n362) );
  AND2_X1 U478 ( .A1(n405), .A2(n455), .ZN(n363) );
  XOR2_X1 U479 ( .A(n503), .B(KEYINPUT80), .Z(n364) );
  XNOR2_X1 U480 ( .A(KEYINPUT48), .B(KEYINPUT71), .ZN(n365) );
  INV_X1 U481 ( .A(KEYINPUT65), .ZN(n400) );
  AND2_X2 U482 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U483 ( .A1(n589), .A2(n686), .ZN(n578) );
  INV_X1 U484 ( .A(n583), .ZN(n573) );
  NAND2_X1 U485 ( .A1(n583), .A2(n687), .ZN(n574) );
  XNOR2_X2 U486 ( .A(n539), .B(KEYINPUT106), .ZN(n583) );
  XNOR2_X1 U487 ( .A(n578), .B(KEYINPUT39), .ZN(n388) );
  XNOR2_X1 U488 ( .A(n369), .B(n478), .ZN(n480) );
  XNOR2_X1 U489 ( .A(n477), .B(n479), .ZN(n369) );
  XNOR2_X1 U490 ( .A(n574), .B(n394), .ZN(n393) );
  XNOR2_X1 U491 ( .A(n370), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X2 U492 ( .A(n371), .B(KEYINPUT40), .ZN(n749) );
  NAND2_X1 U493 ( .A1(n388), .A2(n658), .ZN(n371) );
  NAND2_X1 U494 ( .A1(n393), .A2(n391), .ZN(n390) );
  OR2_X2 U495 ( .A1(n714), .A2(n620), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n423), .B(n426), .ZN(n374) );
  XNOR2_X2 U497 ( .A(n376), .B(n375), .ZN(n748) );
  NAND2_X1 U498 ( .A1(n398), .A2(n517), .ZN(n733) );
  XNOR2_X2 U499 ( .A(n570), .B(n379), .ZN(n398) );
  XNOR2_X1 U500 ( .A(n386), .B(n385), .ZN(n529) );
  NAND2_X1 U501 ( .A1(n553), .A2(n706), .ZN(n386) );
  XNOR2_X2 U502 ( .A(n528), .B(n527), .ZN(n706) );
  XNOR2_X1 U503 ( .A(n737), .B(n508), .ZN(n639) );
  XNOR2_X2 U504 ( .A(n487), .B(n486), .ZN(n737) );
  XNOR2_X1 U505 ( .A(n387), .B(KEYINPUT18), .ZN(n412) );
  NAND2_X1 U506 ( .A1(n388), .A2(n661), .ZN(n664) );
  NAND2_X2 U507 ( .A1(n398), .A2(n397), .ZN(n667) );
  NAND2_X1 U508 ( .A1(n396), .A2(n398), .ZN(n395) );
  NOR2_X1 U509 ( .A1(n738), .A2(n619), .ZN(n396) );
  XNOR2_X2 U510 ( .A(n511), .B(n510), .ZN(n585) );
  NAND2_X1 U511 ( .A1(n617), .A2(G234), .ZN(n446) );
  NAND2_X1 U512 ( .A1(n655), .A2(n692), .ZN(n597) );
  XNOR2_X1 U513 ( .A(n584), .B(n404), .ZN(n403) );
  INV_X1 U514 ( .A(KEYINPUT28), .ZN(n404) );
  NAND2_X1 U515 ( .A1(n408), .A2(n360), .ZN(n622) );
  NAND2_X1 U516 ( .A1(n553), .A2(n362), .ZN(n411) );
  NAND2_X1 U517 ( .A1(n414), .A2(n692), .ZN(n693) );
  NAND2_X1 U518 ( .A1(n418), .A2(n416), .ZN(n415) );
  INV_X1 U519 ( .A(n750), .ZN(n417) );
  XNOR2_X1 U520 ( .A(n588), .B(n587), .ZN(n418) );
  XNOR2_X2 U521 ( .A(n531), .B(n530), .ZN(n563) );
  AND2_X1 U522 ( .A1(n664), .A2(n616), .ZN(n419) );
  INV_X1 U523 ( .A(n674), .ZN(n536) );
  XNOR2_X1 U524 ( .A(n485), .B(n458), .ZN(n459) );
  XNOR2_X1 U525 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U526 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U527 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U528 ( .A(n420), .B(n483), .ZN(n423) );
  INV_X1 U529 ( .A(G128), .ZN(n421) );
  NAND2_X1 U530 ( .A1(G224), .A2(n517), .ZN(n424) );
  XNOR2_X1 U531 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U532 ( .A(G110), .B(G107), .ZN(n428) );
  INV_X1 U533 ( .A(n430), .ZN(n432) );
  XNOR2_X1 U534 ( .A(G113), .B(KEYINPUT3), .ZN(n431) );
  XOR2_X1 U535 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n434) );
  NAND2_X1 U536 ( .A1(G210), .A2(n436), .ZN(n433) );
  XNOR2_X2 U537 ( .A(n435), .B(n361), .ZN(n571) );
  NAND2_X1 U538 ( .A1(G214), .A2(n436), .ZN(n687) );
  NAND2_X1 U539 ( .A1(n571), .A2(n687), .ZN(n516) );
  NAND2_X1 U540 ( .A1(G234), .A2(n517), .ZN(n437) );
  XOR2_X1 U541 ( .A(KEYINPUT8), .B(n437), .Z(n476) );
  NAND2_X1 U542 ( .A1(G221), .A2(n476), .ZN(n443) );
  XOR2_X1 U543 ( .A(G110), .B(G128), .Z(n439) );
  XNOR2_X1 U544 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U545 ( .A(n444), .B(G140), .ZN(n736) );
  XNOR2_X1 U546 ( .A(G146), .B(n736), .ZN(n460) );
  XNOR2_X1 U547 ( .A(n445), .B(n460), .ZN(n722) );
  NOR2_X1 U548 ( .A1(G902), .A2(n722), .ZN(n448) );
  XNOR2_X1 U549 ( .A(KEYINPUT20), .B(n446), .ZN(n453) );
  NAND2_X1 U550 ( .A1(n453), .A2(G217), .ZN(n447) );
  XNOR2_X1 U551 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U552 ( .A(KEYINPUT14), .B(n450), .Z(n702) );
  NOR2_X1 U553 ( .A1(G900), .A2(n517), .ZN(n451) );
  NAND2_X1 U554 ( .A1(n451), .A2(G902), .ZN(n452) );
  NAND2_X1 U555 ( .A1(G952), .A2(n517), .ZN(n518) );
  NAND2_X1 U556 ( .A1(n452), .A2(n518), .ZN(n455) );
  XOR2_X1 U557 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n454) );
  XOR2_X1 U558 ( .A(n577), .B(KEYINPUT72), .Z(n456) );
  NOR2_X1 U559 ( .A1(n575), .A2(n456), .ZN(n582) );
  INV_X1 U560 ( .A(n582), .ZN(n501) );
  NAND2_X1 U561 ( .A1(G214), .A2(n488), .ZN(n458) );
  XNOR2_X1 U562 ( .A(n460), .B(n459), .ZN(n468) );
  XNOR2_X1 U563 ( .A(G113), .B(KEYINPUT12), .ZN(n461) );
  XNOR2_X1 U564 ( .A(n462), .B(n461), .ZN(n466) );
  XOR2_X1 U565 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n464) );
  XNOR2_X1 U566 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U567 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U568 ( .A(n468), .B(n467), .ZN(n632) );
  NAND2_X1 U569 ( .A1(n632), .A2(n498), .ZN(n472) );
  XOR2_X1 U570 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n470) );
  XNOR2_X1 U571 ( .A(KEYINPUT13), .B(G475), .ZN(n469) );
  XOR2_X1 U572 ( .A(n470), .B(n469), .Z(n471) );
  XNOR2_X1 U573 ( .A(n472), .B(n471), .ZN(n554) );
  XOR2_X1 U574 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n474) );
  XNOR2_X1 U575 ( .A(G107), .B(KEYINPUT101), .ZN(n473) );
  XNOR2_X1 U576 ( .A(n474), .B(n473), .ZN(n479) );
  XOR2_X1 U577 ( .A(KEYINPUT7), .B(n475), .Z(n478) );
  NAND2_X1 U578 ( .A1(G217), .A2(n476), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n480), .B(n487), .ZN(n718) );
  NAND2_X1 U580 ( .A1(n718), .A2(n498), .ZN(n481) );
  XNOR2_X2 U581 ( .A(n482), .B(KEYINPUT103), .ZN(n658) );
  XNOR2_X1 U582 ( .A(n483), .B(G137), .ZN(n484) );
  XNOR2_X1 U583 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U584 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n490) );
  NAND2_X1 U585 ( .A1(n488), .A2(G210), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n490), .B(n489), .ZN(n494) );
  XOR2_X1 U587 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n492) );
  XNOR2_X1 U588 ( .A(G116), .B(G101), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U590 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U591 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U592 ( .A1(n625), .A2(n498), .ZN(n499) );
  XNOR2_X2 U593 ( .A(n499), .B(G472), .ZN(n539) );
  INV_X1 U594 ( .A(KEYINPUT6), .ZN(n500) );
  XOR2_X1 U595 ( .A(KEYINPUT112), .B(n609), .Z(n502) );
  NOR2_X1 U596 ( .A1(n516), .A2(n502), .ZN(n504) );
  NAND2_X1 U597 ( .A1(n517), .A2(G227), .ZN(n505) );
  XNOR2_X1 U598 ( .A(n505), .B(G140), .ZN(n506) );
  XNOR2_X1 U599 ( .A(n507), .B(n506), .ZN(n508) );
  INV_X1 U600 ( .A(KEYINPUT73), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n509), .B(G469), .ZN(n510) );
  XNOR2_X1 U602 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n512) );
  XNOR2_X2 U603 ( .A(n585), .B(n512), .ZN(n674) );
  NAND2_X1 U604 ( .A1(n513), .A2(n674), .ZN(n607) );
  XOR2_X1 U605 ( .A(G125), .B(KEYINPUT37), .Z(n514) );
  XNOR2_X1 U606 ( .A(n607), .B(n514), .ZN(G27) );
  XNOR2_X1 U607 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n515) );
  XNOR2_X2 U608 ( .A(n516), .B(n515), .ZN(n594) );
  XNOR2_X1 U609 ( .A(G898), .B(KEYINPUT90), .ZN(n730) );
  NOR2_X1 U610 ( .A1(n517), .A2(n730), .ZN(n727) );
  NAND2_X1 U611 ( .A1(n727), .A2(G902), .ZN(n519) );
  AND2_X1 U612 ( .A1(n519), .A2(n518), .ZN(n520) );
  OR2_X1 U613 ( .A1(n520), .A2(n702), .ZN(n521) );
  NOR2_X2 U614 ( .A1(n594), .A2(n521), .ZN(n525) );
  XNOR2_X1 U615 ( .A(KEYINPUT82), .B(KEYINPUT0), .ZN(n523) );
  INV_X1 U616 ( .A(KEYINPUT68), .ZN(n522) );
  AND2_X1 U617 ( .A1(n575), .A2(n671), .ZN(n673) );
  AND2_X1 U618 ( .A1(n674), .A2(n673), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n550), .A2(n546), .ZN(n528) );
  XNOR2_X1 U620 ( .A(KEYINPUT107), .B(KEYINPUT33), .ZN(n526) );
  XNOR2_X1 U621 ( .A(n526), .B(KEYINPUT83), .ZN(n527) );
  AND2_X1 U622 ( .A1(n532), .A2(n554), .ZN(n591) );
  NAND2_X1 U623 ( .A1(n529), .A2(n591), .ZN(n531) );
  INV_X1 U624 ( .A(KEYINPUT35), .ZN(n530) );
  XNOR2_X1 U625 ( .A(n563), .B(G122), .ZN(G24) );
  NOR2_X1 U626 ( .A1(n554), .A2(n532), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n533), .B(KEYINPUT104), .ZN(n580) );
  INV_X1 U628 ( .A(n580), .ZN(n690) );
  NOR2_X1 U629 ( .A1(n690), .A2(n549), .ZN(n534) );
  NAND2_X1 U630 ( .A1(n534), .A2(n671), .ZN(n535) );
  XOR2_X1 U631 ( .A(KEYINPUT105), .B(n575), .Z(n670) );
  NOR2_X1 U632 ( .A1(n748), .A2(KEYINPUT44), .ZN(n542) );
  NOR2_X1 U633 ( .A1(n674), .A2(n575), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n540), .A2(n573), .ZN(n541) );
  NOR2_X1 U635 ( .A1(n538), .A2(n541), .ZN(n651) );
  NAND2_X1 U636 ( .A1(n542), .A2(n561), .ZN(n544) );
  INV_X1 U637 ( .A(KEYINPUT79), .ZN(n543) );
  NAND2_X1 U638 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U639 ( .A1(n545), .A2(n563), .ZN(n560) );
  NOR2_X1 U640 ( .A1(n378), .A2(n674), .ZN(n547) );
  NAND2_X1 U641 ( .A1(n547), .A2(n368), .ZN(n548) );
  NOR2_X1 U642 ( .A1(n538), .A2(n548), .ZN(n643) );
  INV_X1 U643 ( .A(n643), .ZN(n558) );
  BUF_X1 U644 ( .A(n549), .Z(n551) );
  NAND2_X1 U645 ( .A1(n550), .A2(n677), .ZN(n680) );
  NOR2_X1 U646 ( .A1(n551), .A2(n680), .ZN(n552) );
  XOR2_X1 U647 ( .A(KEYINPUT31), .B(n552), .Z(n662) );
  NOR2_X1 U648 ( .A1(n662), .A2(n646), .ZN(n556) );
  NOR2_X1 U649 ( .A1(n555), .A2(n554), .ZN(n661) );
  NOR2_X1 U650 ( .A1(n658), .A2(n661), .ZN(n603) );
  OR2_X1 U651 ( .A1(n556), .A2(n603), .ZN(n557) );
  AND2_X1 U652 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U653 ( .A1(n560), .A2(n559), .ZN(n569) );
  INV_X1 U654 ( .A(n651), .ZN(n561) );
  NAND2_X1 U655 ( .A1(KEYINPUT44), .A2(n561), .ZN(n562) );
  NOR2_X1 U656 ( .A1(n748), .A2(n562), .ZN(n565) );
  NAND2_X1 U657 ( .A1(n565), .A2(n564), .ZN(n567) );
  OR2_X1 U658 ( .A1(KEYINPUT79), .A2(KEYINPUT44), .ZN(n566) );
  AND2_X2 U659 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X2 U660 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U661 ( .A1(n575), .A2(n585), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n686), .A2(n687), .ZN(n579) );
  XNOR2_X2 U663 ( .A(n581), .B(KEYINPUT41), .ZN(n707) );
  NAND2_X1 U664 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U665 ( .A1(n707), .A2(n596), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n749), .A2(n751), .ZN(n588) );
  XOR2_X1 U667 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n587) );
  NAND2_X1 U668 ( .A1(n613), .A2(n589), .ZN(n590) );
  XNOR2_X1 U669 ( .A(KEYINPUT109), .B(n590), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U671 ( .A(KEYINPUT110), .B(n593), .ZN(n750) );
  INV_X1 U672 ( .A(n603), .ZN(n692) );
  INV_X1 U673 ( .A(n594), .ZN(n595) );
  XNOR2_X1 U674 ( .A(n597), .B(KEYINPUT47), .ZN(n598) );
  INV_X1 U675 ( .A(KEYINPUT77), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n598), .A2(n602), .ZN(n601) );
  NAND2_X1 U677 ( .A1(KEYINPUT47), .A2(n655), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n599), .A2(KEYINPUT77), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  AND2_X1 U683 ( .A1(n609), .A2(n687), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n610), .A2(n536), .ZN(n612) );
  XNOR2_X1 U685 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n612), .B(n611), .ZN(n615) );
  INV_X1 U687 ( .A(n613), .ZN(n614) );
  AND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n665) );
  INV_X1 U689 ( .A(n665), .ZN(n616) );
  NOR2_X1 U690 ( .A1(n617), .A2(KEYINPUT78), .ZN(n618) );
  NOR2_X1 U691 ( .A1(n618), .A2(KEYINPUT2), .ZN(n619) );
  INV_X1 U692 ( .A(n622), .ZN(n621) );
  INV_X1 U693 ( .A(KEYINPUT2), .ZN(n666) );
  AND2_X1 U694 ( .A1(n666), .A2(n622), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n721), .A2(G472), .ZN(n627) );
  XOR2_X1 U696 ( .A(KEYINPUT62), .B(n625), .Z(n626) );
  INV_X1 U697 ( .A(G952), .ZN(n628) );
  XNOR2_X1 U698 ( .A(KEYINPUT81), .B(KEYINPUT63), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n631), .B(n630), .ZN(G57) );
  NAND2_X1 U700 ( .A1(n721), .A2(G475), .ZN(n634) );
  XNOR2_X1 U701 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X2 U702 ( .A1(n635), .A2(n726), .ZN(n637) );
  XOR2_X1 U703 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n636) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(G60) );
  NAND2_X1 U705 ( .A1(n721), .A2(G469), .ZN(n641) );
  XOR2_X1 U706 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U708 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U709 ( .A1(n642), .A2(n726), .ZN(G54) );
  XOR2_X1 U710 ( .A(G101), .B(n643), .Z(G3) );
  XOR2_X1 U711 ( .A(G104), .B(KEYINPUT113), .Z(n645) );
  NAND2_X1 U712 ( .A1(n646), .A2(n658), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n645), .B(n644), .ZN(G6) );
  XNOR2_X1 U714 ( .A(G107), .B(KEYINPUT114), .ZN(n650) );
  XOR2_X1 U715 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n648) );
  NAND2_X1 U716 ( .A1(n646), .A2(n661), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(G9) );
  XOR2_X1 U719 ( .A(G110), .B(n651), .Z(G12) );
  XOR2_X1 U720 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n653) );
  NAND2_X1 U721 ( .A1(n655), .A2(n661), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U723 ( .A(G128), .B(n654), .Z(G30) );
  NAND2_X1 U724 ( .A1(n655), .A2(n658), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n656), .B(KEYINPUT116), .ZN(n657) );
  XNOR2_X1 U726 ( .A(G146), .B(n657), .ZN(G48) );
  XOR2_X1 U727 ( .A(G113), .B(KEYINPUT117), .Z(n660) );
  NAND2_X1 U728 ( .A1(n662), .A2(n658), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(G116), .ZN(G18) );
  XNOR2_X1 U732 ( .A(G134), .B(n664), .ZN(G36) );
  XOR2_X1 U733 ( .A(G140), .B(n665), .Z(G42) );
  AND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n711) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT49), .ZN(n679) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n675), .B(KEYINPUT50), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U744 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n682) );
  XNOR2_X1 U745 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U746 ( .A1(n707), .A2(n684), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n685), .B(KEYINPUT119), .ZN(n699) );
  NOR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT120), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n691), .B(KEYINPUT121), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U753 ( .A(KEYINPUT122), .B(n695), .Z(n697) );
  INV_X1 U754 ( .A(n706), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n700), .B(KEYINPUT52), .ZN(n701) );
  NOR2_X1 U758 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U759 ( .A1(n703), .A2(G952), .ZN(n704) );
  XNOR2_X1 U760 ( .A(KEYINPUT123), .B(n704), .ZN(n705) );
  NOR2_X1 U761 ( .A1(G953), .A2(n705), .ZN(n709) );
  NAND2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U763 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U765 ( .A(KEYINPUT53), .B(n712), .ZN(G75) );
  NAND2_X1 U766 ( .A1(n721), .A2(G210), .ZN(n716) );
  XOR2_X1 U767 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n713) );
  XNOR2_X1 U768 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U769 ( .A1(n721), .A2(G478), .ZN(n719) );
  XOR2_X1 U770 ( .A(n719), .B(n718), .Z(n720) );
  NOR2_X1 U771 ( .A1(n726), .A2(n720), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n721), .A2(G217), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n722), .B(KEYINPUT124), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U775 ( .A1(n726), .A2(n725), .ZN(G66) );
  NOR2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n735) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U778 ( .A(KEYINPUT61), .B(n729), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U781 ( .A(n735), .B(n734), .ZN(G69) );
  XNOR2_X1 U782 ( .A(n737), .B(n736), .ZN(n741) );
  XNOR2_X1 U783 ( .A(n738), .B(n741), .ZN(n739) );
  NOR2_X1 U784 ( .A1(G953), .A2(n739), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n740), .B(KEYINPUT125), .ZN(n746) );
  XOR2_X1 U786 ( .A(G227), .B(n741), .Z(n742) );
  XNOR2_X1 U787 ( .A(n742), .B(KEYINPUT126), .ZN(n743) );
  NAND2_X1 U788 ( .A1(n743), .A2(G900), .ZN(n744) );
  NAND2_X1 U789 ( .A1(G953), .A2(n744), .ZN(n745) );
  NAND2_X1 U790 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U791 ( .A(KEYINPUT127), .B(n747), .Z(G72) );
  XOR2_X1 U792 ( .A(G119), .B(n748), .Z(G21) );
  XNOR2_X1 U793 ( .A(n749), .B(G131), .ZN(G33) );
  XNOR2_X1 U794 ( .A(G143), .B(n750), .ZN(G45) );
  XNOR2_X1 U795 ( .A(n751), .B(G137), .ZN(G39) );
endmodule

