

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U323 ( .A(n365), .B(KEYINPUT77), .Z(n291) );
  XNOR2_X1 U324 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n424) );
  XNOR2_X1 U325 ( .A(n425), .B(n424), .ZN(n448) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n421) );
  XNOR2_X1 U327 ( .A(n422), .B(n421), .ZN(n546) );
  XOR2_X1 U328 ( .A(KEYINPUT78), .B(n558), .Z(n539) );
  NOR2_X1 U329 ( .A1(n530), .A2(n450), .ZN(n564) );
  XOR2_X1 U330 ( .A(n329), .B(n328), .Z(n530) );
  XNOR2_X1 U331 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U332 ( .A(n454), .B(n453), .ZN(G1349GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n301) );
  INV_X1 U334 ( .A(KEYINPUT75), .ZN(n292) );
  NAND2_X1 U335 ( .A1(KEYINPUT73), .A2(n292), .ZN(n295) );
  INV_X1 U336 ( .A(KEYINPUT73), .ZN(n293) );
  NAND2_X1 U337 ( .A1(n293), .A2(KEYINPUT75), .ZN(n294) );
  NAND2_X1 U338 ( .A1(n295), .A2(n294), .ZN(n297) );
  XNOR2_X1 U339 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n299) );
  XNOR2_X1 U341 ( .A(G176GAT), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n298), .B(G64GAT), .ZN(n351) );
  XNOR2_X1 U343 ( .A(n299), .B(n351), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U345 ( .A(G148GAT), .B(G78GAT), .Z(n334) );
  XOR2_X1 U346 ( .A(KEYINPUT13), .B(G57GAT), .Z(n379) );
  XOR2_X1 U347 ( .A(n334), .B(n379), .Z(n303) );
  NAND2_X1 U348 ( .A1(G230GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U350 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U351 ( .A(G120GAT), .B(G71GAT), .Z(n321) );
  XOR2_X1 U352 ( .A(KEYINPUT74), .B(G85GAT), .Z(n307) );
  XNOR2_X1 U353 ( .A(G99GAT), .B(G92GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(G106GAT), .B(n308), .Z(n372) );
  XNOR2_X1 U356 ( .A(n321), .B(n372), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n577) );
  XOR2_X1 U358 ( .A(n577), .B(KEYINPUT41), .Z(n550) );
  XOR2_X1 U359 ( .A(n550), .B(KEYINPUT104), .Z(n533) );
  XOR2_X1 U360 ( .A(G176GAT), .B(KEYINPUT83), .Z(n312) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G113GAT), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n329) );
  XOR2_X1 U363 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n314) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U366 ( .A(n315), .B(KEYINPUT85), .Z(n320) );
  XNOR2_X1 U367 ( .A(KEYINPUT82), .B(KEYINPUT0), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n316), .B(KEYINPUT81), .ZN(n435) );
  XOR2_X1 U369 ( .A(G183GAT), .B(KEYINPUT17), .Z(n318) );
  XNOR2_X1 U370 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n347) );
  XNOR2_X1 U372 ( .A(n435), .B(n347), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U374 ( .A(G190GAT), .B(G134GAT), .Z(n323) );
  XOR2_X1 U375 ( .A(G15GAT), .B(G127GAT), .Z(n380) );
  XNOR2_X1 U376 ( .A(n380), .B(n321), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U378 ( .A(n325), .B(n324), .Z(n327) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(G99GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n331) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G162GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n345) );
  XOR2_X1 U384 ( .A(G211GAT), .B(KEYINPUT21), .Z(n333) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n352) );
  XOR2_X1 U387 ( .A(n352), .B(n334), .Z(n336) );
  NAND2_X1 U388 ( .A1(G228GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U390 ( .A(n337), .B(KEYINPUT22), .Z(n340) );
  XNOR2_X1 U391 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n338), .B(KEYINPUT2), .ZN(n434) );
  XNOR2_X1 U393 ( .A(n434), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U395 ( .A(n341), .B(G218GAT), .Z(n343) );
  XOR2_X1 U396 ( .A(G141GAT), .B(G22GAT), .Z(n402) );
  XNOR2_X1 U397 ( .A(G50GAT), .B(n402), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U399 ( .A(n345), .B(n344), .Z(n467) );
  XNOR2_X1 U400 ( .A(G36GAT), .B(G190GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n346), .B(G218GAT), .ZN(n365) );
  XNOR2_X1 U402 ( .A(n347), .B(n365), .ZN(n359) );
  XOR2_X1 U403 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n349) );
  NAND2_X1 U404 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U406 ( .A(n350), .B(KEYINPUT90), .Z(n354) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U409 ( .A(n355), .B(KEYINPUT92), .Z(n357) );
  XOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .Z(n399) );
  XNOR2_X1 U411 ( .A(n399), .B(G92GAT), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n359), .B(n358), .Z(n519) );
  XOR2_X1 U414 ( .A(KEYINPUT118), .B(n519), .Z(n423) );
  INV_X1 U415 ( .A(KEYINPUT36), .ZN(n376) );
  XOR2_X1 U416 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n361) );
  XNOR2_X1 U417 ( .A(KEYINPUT66), .B(KEYINPUT11), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U419 ( .A(n362), .B(KEYINPUT76), .Z(n364) );
  XOR2_X1 U420 ( .A(G134GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U421 ( .A(n439), .B(KEYINPUT10), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n368) );
  NAND2_X1 U423 ( .A1(G232GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n291), .B(n366), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n375) );
  XOR2_X1 U426 ( .A(KEYINPUT7), .B(G50GAT), .Z(n370) );
  XNOR2_X1 U427 ( .A(G43GAT), .B(G29GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U429 ( .A(KEYINPUT8), .B(n371), .Z(n411) );
  INV_X1 U430 ( .A(n411), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n558) );
  XNOR2_X1 U433 ( .A(n376), .B(n539), .ZN(n486) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n378) );
  XNOR2_X1 U435 ( .A(KEYINPUT15), .B(KEYINPUT79), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U437 ( .A(n379), .B(G71GAT), .Z(n382) );
  XNOR2_X1 U438 ( .A(G183GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U440 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U441 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n394) );
  XOR2_X1 U443 ( .A(G211GAT), .B(G78GAT), .Z(n388) );
  XNOR2_X1 U444 ( .A(G22GAT), .B(G155GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U446 ( .A(KEYINPUT80), .B(G64GAT), .Z(n390) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(G8GAT), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(n392), .B(n391), .Z(n393) );
  XOR2_X1 U450 ( .A(n394), .B(n393), .Z(n580) );
  NOR2_X1 U451 ( .A1(n486), .A2(n580), .ZN(n395) );
  XNOR2_X1 U452 ( .A(KEYINPUT45), .B(n395), .ZN(n396) );
  NAND2_X1 U453 ( .A1(n396), .A2(n577), .ZN(n413) );
  XOR2_X1 U454 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n398) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(KEYINPUT30), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n410) );
  XNOR2_X1 U457 ( .A(G15GAT), .B(G36GAT), .ZN(n401) );
  XOR2_X1 U458 ( .A(G113GAT), .B(G1GAT), .Z(n438) );
  XNOR2_X1 U459 ( .A(n438), .B(n399), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n405) );
  NAND2_X1 U463 ( .A1(G229GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U465 ( .A(KEYINPUT29), .B(n406), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n412) );
  XOR2_X1 U468 ( .A(n412), .B(n411), .Z(n572) );
  XNOR2_X1 U469 ( .A(KEYINPUT71), .B(n572), .ZN(n561) );
  NOR2_X1 U470 ( .A1(n413), .A2(n561), .ZN(n420) );
  OR2_X1 U471 ( .A1(n550), .A2(n572), .ZN(n415) );
  INV_X1 U472 ( .A(KEYINPUT46), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  INV_X1 U474 ( .A(n580), .ZN(n563) );
  NOR2_X1 U475 ( .A1(n416), .A2(n563), .ZN(n417) );
  NAND2_X1 U476 ( .A1(n558), .A2(n417), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n418), .B(KEYINPUT47), .ZN(n419) );
  NOR2_X1 U478 ( .A1(n420), .A2(n419), .ZN(n422) );
  INV_X1 U479 ( .A(n546), .ZN(n527) );
  NAND2_X1 U480 ( .A1(n423), .A2(n527), .ZN(n425) );
  XOR2_X1 U481 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n427) );
  XNOR2_X1 U482 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n447) );
  XOR2_X1 U484 ( .A(G148GAT), .B(G120GAT), .Z(n429) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(G127GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U487 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n431) );
  XNOR2_X1 U488 ( .A(G57GAT), .B(KEYINPUT88), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U490 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U493 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U496 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U497 ( .A(G29GAT), .B(G85GAT), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n516) );
  NAND2_X1 U500 ( .A1(n448), .A2(n516), .ZN(n570) );
  NOR2_X1 U501 ( .A1(n467), .A2(n570), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  NAND2_X1 U503 ( .A1(n533), .A2(n564), .ZN(n454) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT120), .Z(n452) );
  XNOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n451) );
  INV_X1 U506 ( .A(G190GAT), .ZN(n458) );
  NAND2_X1 U507 ( .A1(n564), .A2(n539), .ZN(n456) );
  XOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n460) );
  XNOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n480) );
  NAND2_X1 U514 ( .A1(n561), .A2(n577), .ZN(n490) );
  NOR2_X1 U515 ( .A1(n539), .A2(n580), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT16), .ZN(n477) );
  XNOR2_X1 U517 ( .A(n519), .B(KEYINPUT27), .ZN(n470) );
  NOR2_X1 U518 ( .A1(n470), .A2(n516), .ZN(n462) );
  XOR2_X1 U519 ( .A(KEYINPUT94), .B(n462), .Z(n545) );
  XOR2_X1 U520 ( .A(n467), .B(KEYINPUT28), .Z(n524) );
  INV_X1 U521 ( .A(n524), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n545), .A2(n463), .ZN(n528) );
  NAND2_X1 U523 ( .A1(n530), .A2(n528), .ZN(n476) );
  NOR2_X1 U524 ( .A1(n530), .A2(n519), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n467), .A2(n464), .ZN(n465) );
  XOR2_X1 U526 ( .A(n465), .B(KEYINPUT25), .Z(n466) );
  XNOR2_X1 U527 ( .A(KEYINPUT96), .B(n466), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT95), .B(KEYINPUT26), .Z(n469) );
  NAND2_X1 U529 ( .A1(n467), .A2(n530), .ZN(n468) );
  XOR2_X1 U530 ( .A(n469), .B(n468), .Z(n547) );
  INV_X1 U531 ( .A(n547), .ZN(n569) );
  NOR2_X1 U532 ( .A1(n569), .A2(n470), .ZN(n471) );
  NOR2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U534 ( .A(KEYINPUT97), .B(n473), .ZN(n474) );
  NAND2_X1 U535 ( .A1(n474), .A2(n516), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n488) );
  NAND2_X1 U537 ( .A1(n477), .A2(n488), .ZN(n502) );
  NOR2_X1 U538 ( .A1(n490), .A2(n502), .ZN(n478) );
  XOR2_X1 U539 ( .A(KEYINPUT98), .B(n478), .Z(n484) );
  NOR2_X1 U540 ( .A1(n484), .A2(n516), .ZN(n479) );
  XOR2_X1 U541 ( .A(n480), .B(n479), .Z(G1324GAT) );
  NOR2_X1 U542 ( .A1(n484), .A2(n519), .ZN(n481) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n483) );
  NOR2_X1 U545 ( .A1(n530), .A2(n484), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U547 ( .A1(n524), .A2(n484), .ZN(n485) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  NOR2_X1 U549 ( .A1(n563), .A2(n486), .ZN(n487) );
  AND2_X1 U550 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT37), .B(n489), .ZN(n515) );
  NOR2_X1 U552 ( .A1(n515), .A2(n490), .ZN(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(n491), .Z(n500) );
  NOR2_X1 U554 ( .A1(n500), .A2(n516), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n500), .A2(n519), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n497) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n499) );
  NOR2_X1 U563 ( .A1(n530), .A2(n500), .ZN(n498) );
  XOR2_X1 U564 ( .A(n499), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U565 ( .A1(n524), .A2(n500), .ZN(n501) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  NAND2_X1 U567 ( .A1(n533), .A2(n572), .ZN(n514) );
  OR2_X1 U568 ( .A1(n502), .A2(n514), .ZN(n510) );
  NOR2_X1 U569 ( .A1(n516), .A2(n510), .ZN(n504) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n519), .A2(n510), .ZN(n506) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(n506), .Z(n507) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NOR2_X1 U576 ( .A1(n530), .A2(n510), .ZN(n509) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U579 ( .A1(n524), .A2(n510), .ZN(n512) );
  XNOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U581 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  OR2_X1 U583 ( .A1(n515), .A2(n514), .ZN(n523) );
  NOR2_X1 U584 ( .A1(n516), .A2(n523), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n519), .A2(n523), .ZN(n520) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(n520), .Z(n521) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NOR2_X1 U590 ( .A1(n530), .A2(n523), .ZN(n522) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n525), .Z(n526) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT111), .B(n531), .Z(n540) );
  NAND2_X1 U598 ( .A1(n540), .A2(n561), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U601 ( .A1(n540), .A2(n533), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n563), .A2(n540), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT113), .Z(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n572), .A2(n557), .ZN(n549) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n557), .A2(n550), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT52), .B(KEYINPUT115), .Z(n552) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n580), .A2(n557), .ZN(n555) );
  XOR2_X1 U622 ( .A(KEYINPUT116), .B(n555), .Z(n556) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT121), .Z(n566) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n576) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT123), .ZN(n582) );
  NOR2_X1 U637 ( .A1(n572), .A2(n582), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n582), .ZN(n579) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n486), .A2(n582), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

