

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  INV_X1 U323 ( .A(n421), .ZN(n425) );
  INV_X1 U324 ( .A(KEYINPUT120), .ZN(n473) );
  XNOR2_X1 U325 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  XNOR2_X1 U326 ( .A(n421), .B(n335), .ZN(n336) );
  XNOR2_X1 U327 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U328 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U329 ( .A(n356), .B(n336), .ZN(n337) );
  INV_X1 U330 ( .A(KEYINPUT99), .ZN(n409) );
  XNOR2_X1 U331 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U332 ( .A(n410), .B(n409), .ZN(n491) );
  XNOR2_X1 U333 ( .A(KEYINPUT37), .B(n450), .ZN(n528) );
  INV_X1 U334 ( .A(G211GAT), .ZN(n479) );
  XOR2_X1 U335 ( .A(KEYINPUT81), .B(n465), .Z(n550) );
  XOR2_X1 U336 ( .A(KEYINPUT28), .B(n482), .Z(n536) );
  XNOR2_X1 U337 ( .A(n479), .B(KEYINPUT126), .ZN(n480) );
  XNOR2_X1 U338 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U339 ( .A(n481), .B(n480), .ZN(G1354GAT) );
  XNOR2_X1 U340 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT107), .B(KEYINPUT38), .Z(n453) );
  XOR2_X1 U342 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n292) );
  XNOR2_X1 U343 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U345 ( .A(G1GAT), .B(KEYINPUT71), .Z(n433) );
  XOR2_X1 U346 ( .A(G29GAT), .B(KEYINPUT8), .Z(n294) );
  XNOR2_X1 U347 ( .A(KEYINPUT70), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n418) );
  XOR2_X1 U349 ( .A(n433), .B(n418), .Z(n296) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G50GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n311) );
  XOR2_X1 U353 ( .A(G113GAT), .B(G15GAT), .Z(n300) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G36GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U356 ( .A(G8GAT), .B(G141GAT), .Z(n302) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(G197GAT), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U359 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U360 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n306) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT65), .B(n307), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U365 ( .A(n311), .B(n310), .Z(n513) );
  XOR2_X1 U366 ( .A(G64GAT), .B(KEYINPUT76), .Z(n313) );
  XNOR2_X1 U367 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(n314), .B(G92GAT), .Z(n316) );
  XOR2_X1 U370 ( .A(G120GAT), .B(G71GAT), .Z(n368) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(n368), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n329) );
  XNOR2_X1 U373 ( .A(G99GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n317), .B(G85GAT), .ZN(n417) );
  XOR2_X1 U375 ( .A(n417), .B(KEYINPUT74), .Z(n319) );
  NAND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U378 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n321) );
  XNOR2_X1 U379 ( .A(KEYINPUT32), .B(KEYINPUT77), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U381 ( .A(n323), .B(n322), .Z(n327) );
  XNOR2_X1 U382 ( .A(G78GAT), .B(KEYINPUT75), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n324), .B(G148GAT), .ZN(n349) );
  XNOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n325), .B(KEYINPUT13), .ZN(n436) );
  XNOR2_X1 U386 ( .A(n349), .B(n436), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n462) );
  NAND2_X1 U389 ( .A1(n513), .A2(n462), .ZN(n493) );
  INV_X1 U390 ( .A(n493), .ZN(n451) );
  XOR2_X1 U391 ( .A(G8GAT), .B(G64GAT), .Z(n431) );
  XOR2_X1 U392 ( .A(KEYINPUT87), .B(G211GAT), .Z(n331) );
  XNOR2_X1 U393 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U395 ( .A(G197GAT), .B(n332), .Z(n356) );
  XOR2_X1 U396 ( .A(G92GAT), .B(G218GAT), .Z(n334) );
  XNOR2_X1 U397 ( .A(G36GAT), .B(G190GAT), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n421) );
  XOR2_X1 U399 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n335) );
  XOR2_X1 U400 ( .A(n431), .B(n337), .Z(n339) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n345) );
  XNOR2_X1 U403 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n340), .B(KEYINPUT19), .ZN(n341) );
  XOR2_X1 U405 ( .A(n341), .B(KEYINPUT17), .Z(n343) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G176GAT), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n364) );
  INV_X1 U408 ( .A(n364), .ZN(n344) );
  XOR2_X1 U409 ( .A(n345), .B(n344), .Z(n532) );
  INV_X1 U410 ( .A(n532), .ZN(n520) );
  XNOR2_X1 U411 ( .A(n520), .B(KEYINPUT27), .ZN(n405) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n347) );
  XOR2_X1 U413 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XOR2_X1 U414 ( .A(G22GAT), .B(G155GAT), .Z(n430) );
  XNOR2_X1 U415 ( .A(n422), .B(n430), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U417 ( .A(n348), .B(G106GAT), .Z(n354) );
  XOR2_X1 U418 ( .A(n349), .B(KEYINPUT24), .Z(n351) );
  NAND2_X1 U419 ( .A1(G228GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n352), .B(G218GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT89), .B(KEYINPUT2), .Z(n358) );
  XNOR2_X1 U425 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U427 ( .A(G141GAT), .B(n359), .ZN(n398) );
  XNOR2_X1 U428 ( .A(n360), .B(n398), .ZN(n482) );
  XOR2_X1 U429 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n362) );
  XNOR2_X1 U430 ( .A(G99GAT), .B(G190GAT), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n364), .B(n363), .ZN(n372) );
  XOR2_X1 U433 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XOR2_X1 U434 ( .A(n432), .B(KEYINPUT84), .Z(n366) );
  NAND2_X1 U435 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U437 ( .A(G43GAT), .B(G134GAT), .Z(n423) );
  XOR2_X1 U438 ( .A(n367), .B(n423), .Z(n370) );
  XOR2_X1 U439 ( .A(G113GAT), .B(KEYINPUT0), .Z(n394) );
  XNOR2_X1 U440 ( .A(n368), .B(n394), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n372), .B(n371), .ZN(n534) );
  NOR2_X1 U443 ( .A1(n482), .A2(n534), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n373), .B(KEYINPUT26), .ZN(n555) );
  NAND2_X1 U445 ( .A1(n405), .A2(n555), .ZN(n378) );
  INV_X1 U446 ( .A(n534), .ZN(n374) );
  OR2_X1 U447 ( .A1(n374), .A2(n532), .ZN(n375) );
  NAND2_X1 U448 ( .A1(n482), .A2(n375), .ZN(n376) );
  XOR2_X1 U449 ( .A(KEYINPUT25), .B(n376), .Z(n377) );
  NAND2_X1 U450 ( .A1(n378), .A2(n377), .ZN(n403) );
  XOR2_X1 U451 ( .A(G57GAT), .B(KEYINPUT90), .Z(n380) );
  XNOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT95), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U454 ( .A(G155GAT), .B(G148GAT), .Z(n382) );
  XNOR2_X1 U455 ( .A(G120GAT), .B(G127GAT), .ZN(n381) );
  XNOR2_X1 U456 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U457 ( .A(n384), .B(n383), .ZN(n402) );
  XOR2_X1 U458 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n386) );
  XNOR2_X1 U459 ( .A(KEYINPUT1), .B(KEYINPUT91), .ZN(n385) );
  XNOR2_X1 U460 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n388) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n387) );
  XNOR2_X1 U463 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U464 ( .A(n390), .B(n389), .Z(n400) );
  XOR2_X1 U465 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(G134GAT), .ZN(n391) );
  XNOR2_X1 U467 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U468 ( .A(n394), .B(n393), .Z(n396) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U470 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U471 ( .A(n398), .B(n397), .Z(n399) );
  XNOR2_X1 U472 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n517) );
  INV_X1 U474 ( .A(n517), .ZN(n529) );
  NAND2_X1 U475 ( .A1(n403), .A2(n529), .ZN(n404) );
  XNOR2_X1 U476 ( .A(n404), .B(KEYINPUT98), .ZN(n408) );
  XOR2_X1 U477 ( .A(n534), .B(KEYINPUT86), .Z(n406) );
  NAND2_X1 U478 ( .A1(n517), .A2(n405), .ZN(n553) );
  NOR2_X1 U479 ( .A1(n553), .A2(n536), .ZN(n542) );
  NAND2_X1 U480 ( .A1(n406), .A2(n542), .ZN(n407) );
  NAND2_X1 U481 ( .A1(n408), .A2(n407), .ZN(n410) );
  XOR2_X1 U482 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n412) );
  XNOR2_X1 U483 ( .A(KEYINPUT10), .B(KEYINPUT78), .ZN(n411) );
  XNOR2_X1 U484 ( .A(n412), .B(n411), .ZN(n429) );
  XOR2_X1 U485 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n414) );
  NAND2_X1 U486 ( .A1(G232GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U487 ( .A(n414), .B(n413), .ZN(n416) );
  INV_X1 U488 ( .A(KEYINPUT9), .ZN(n415) );
  XNOR2_X1 U489 ( .A(n416), .B(n415), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n420), .B(n419), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n465) );
  XNOR2_X1 U494 ( .A(KEYINPUT36), .B(n550), .ZN(n457) );
  XOR2_X1 U495 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U498 ( .A(n436), .B(KEYINPUT83), .Z(n438) );
  NAND2_X1 U499 ( .A1(G231GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U501 ( .A(n440), .B(n439), .Z(n448) );
  XOR2_X1 U502 ( .A(G78GAT), .B(G211GAT), .Z(n442) );
  XNOR2_X1 U503 ( .A(G183GAT), .B(G71GAT), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U505 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n444) );
  XNOR2_X1 U506 ( .A(KEYINPUT12), .B(KEYINPUT82), .ZN(n443) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n489) );
  NOR2_X1 U510 ( .A1(n457), .A2(n489), .ZN(n449) );
  NAND2_X1 U511 ( .A1(n491), .A2(n449), .ZN(n450) );
  NAND2_X1 U512 ( .A1(n451), .A2(n528), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT106), .B(n454), .Z(n511) );
  NAND2_X1 U515 ( .A1(n511), .A2(n534), .ZN(n456) );
  INV_X1 U516 ( .A(KEYINPUT123), .ZN(n478) );
  INV_X1 U517 ( .A(n489), .ZN(n576) );
  NOR2_X1 U518 ( .A1(n457), .A2(n576), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT45), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n459), .A2(n462), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT113), .ZN(n461) );
  INV_X1 U522 ( .A(n513), .ZN(n580) );
  NAND2_X1 U523 ( .A1(n461), .A2(n580), .ZN(n470) );
  XOR2_X1 U524 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n468) );
  XOR2_X2 U525 ( .A(n462), .B(KEYINPUT41), .Z(n572) );
  NOR2_X1 U526 ( .A1(n580), .A2(n572), .ZN(n463) );
  XNOR2_X1 U527 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  NOR2_X1 U528 ( .A1(n489), .A2(n464), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT48), .B(n471), .Z(n554) );
  XNOR2_X1 U533 ( .A(n520), .B(KEYINPUT119), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n554), .A2(n472), .ZN(n475) );
  NOR2_X1 U535 ( .A1(n517), .A2(n476), .ZN(n483) );
  NAND2_X1 U536 ( .A1(n483), .A2(n555), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n586) );
  NOR2_X1 U538 ( .A1(n586), .A2(n576), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U540 ( .A(n484), .B(KEYINPUT55), .ZN(n485) );
  NAND2_X1 U541 ( .A1(n485), .A2(n534), .ZN(n575) );
  NOR2_X1 U542 ( .A1(n550), .A2(n575), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT58), .B(n486), .ZN(n488) );
  INV_X1 U544 ( .A(G190GAT), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  NAND2_X1 U546 ( .A1(n489), .A2(n550), .ZN(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n490), .Z(n492) );
  NAND2_X1 U548 ( .A1(n492), .A2(n491), .ZN(n514) );
  NOR2_X1 U549 ( .A1(n493), .A2(n514), .ZN(n504) );
  NAND2_X1 U550 ( .A1(n504), .A2(n517), .ZN(n497) );
  XOR2_X1 U551 ( .A(KEYINPUT101), .B(KEYINPUT34), .Z(n495) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n497), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n504), .A2(n520), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(KEYINPUT102), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G8GAT), .B(n499), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n501) );
  NAND2_X1 U559 ( .A1(n504), .A2(n534), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(n503) );
  XOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT103), .Z(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n536), .A2(n504), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n505), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT105), .B(KEYINPUT108), .Z(n507) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(n509) );
  NAND2_X1 U568 ( .A1(n511), .A2(n517), .ZN(n508) );
  XOR2_X1 U569 ( .A(n509), .B(n508), .Z(G1328GAT) );
  NAND2_X1 U570 ( .A1(n511), .A2(n520), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n536), .A2(n511), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U574 ( .A1(n513), .A2(n572), .ZN(n527) );
  INV_X1 U575 ( .A(n527), .ZN(n515) );
  NOR2_X1 U576 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U577 ( .A(KEYINPUT109), .B(n516), .Z(n524) );
  NAND2_X1 U578 ( .A1(n517), .A2(n524), .ZN(n518) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n518), .ZN(n519) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n524), .A2(n520), .ZN(n521) );
  XNOR2_X1 U582 ( .A(n521), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n524), .A2(n534), .ZN(n522) );
  XNOR2_X1 U584 ( .A(n522), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n523), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n526) );
  NAND2_X1 U587 ( .A1(n524), .A2(n536), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n537) );
  NOR2_X1 U590 ( .A1(n529), .A2(n537), .ZN(n531) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n531), .B(n530), .ZN(G1336GAT) );
  NOR2_X1 U593 ( .A1(n532), .A2(n537), .ZN(n533) );
  XOR2_X1 U594 ( .A(G92GAT), .B(n533), .Z(G1337GAT) );
  NOR2_X1 U595 ( .A1(n374), .A2(n537), .ZN(n535) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n535), .Z(G1338GAT) );
  INV_X1 U597 ( .A(n536), .ZN(n538) );
  NOR2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U599 ( .A(KEYINPUT44), .B(n539), .Z(n540) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U601 ( .A1(n374), .A2(n554), .ZN(n541) );
  NAND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n549) );
  NOR2_X1 U603 ( .A1(n580), .A2(n549), .ZN(n543) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n543), .Z(G1340GAT) );
  NOR2_X1 U605 ( .A1(n572), .A2(n549), .ZN(n545) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U608 ( .A1(n576), .A2(n549), .ZN(n547) );
  XNOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  NOR2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n566) );
  NOR2_X1 U617 ( .A1(n580), .A2(n566), .ZN(n558) );
  XNOR2_X1 U618 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U619 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  NOR2_X1 U621 ( .A1(n572), .A2(n566), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n561) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U625 ( .A(KEYINPUT117), .B(n562), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n576), .A2(n566), .ZN(n565) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n565), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n465), .A2(n566), .ZN(n567) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NOR2_X1 U631 ( .A1(n580), .A2(n575), .ZN(n569) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n571) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n574) );
  NOR2_X1 U637 ( .A1(n575), .A2(n572), .ZN(n573) );
  XOR2_X1 U638 ( .A(n574), .B(n573), .Z(G1349GAT) );
  NOR2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n577), .Z(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n582) );
  NOR2_X1 U644 ( .A1(n580), .A2(n586), .ZN(n581) );
  XOR2_X1 U645 ( .A(n582), .B(n581), .Z(G1352GAT) );
  NOR2_X1 U646 ( .A1(n586), .A2(n462), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NOR2_X1 U650 ( .A1(n457), .A2(n586), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

