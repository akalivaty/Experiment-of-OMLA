//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  INV_X1    g001(.A(G71gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT72), .ZN(new_n205));
  INV_X1    g004(.A(G99gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  INV_X1    g011(.A(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G127gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT68), .ZN(new_n215));
  INV_X1    g014(.A(G113gat), .ZN(new_n216));
  INV_X1    g015(.A(G120gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g018(.A1(G113gat), .A2(G120gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n213), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT69), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(G113gat), .A2(G120gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G113gat), .A2(G120gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(KEYINPUT23), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT64), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n235), .A2(new_n242), .A3(KEYINPUT23), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n236), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n242), .B1(new_n235), .B2(KEYINPUT23), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n240), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT65), .A3(new_n236), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  INV_X1    g050(.A(G183gat), .ZN(new_n252));
  INV_X1    g051(.A(G190gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT25), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n246), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n239), .A2(KEYINPUT26), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n234), .B1(new_n239), .B2(KEYINPUT26), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n258), .A2(new_n259), .B1(G183gat), .B2(G190gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n252), .A2(KEYINPUT27), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT27), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n261), .B2(new_n263), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(G190gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n265), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n261), .A2(new_n263), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n267), .B1(new_n271), .B2(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n260), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n251), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n253), .ZN(new_n278));
  NAND4_X1  g077(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(new_n249), .A3(new_n236), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT25), .ZN(new_n282));
  AND4_X1   g081(.A1(new_n233), .A2(new_n257), .A3(new_n274), .A4(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n262), .A2(G183gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n252), .A2(KEYINPUT27), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT67), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n268), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n272), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n289), .A2(new_n260), .B1(new_n281), .B2(KEYINPUT25), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n233), .B1(new_n290), .B2(new_n257), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G227gat), .ZN(new_n293));
  INV_X1    g092(.A(G233gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT70), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n257), .A2(new_n274), .A3(new_n282), .ZN(new_n297));
  INV_X1    g096(.A(new_n233), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n290), .A2(new_n233), .A3(new_n257), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n299), .A2(KEYINPUT70), .A3(new_n295), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT32), .B(new_n210), .C1(new_n296), .C2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n208), .A2(KEYINPUT32), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n296), .B2(new_n302), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n207), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n299), .A2(new_n295), .A3(new_n300), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n305), .B1(new_n312), .B2(new_n301), .ZN(new_n313));
  INV_X1    g112(.A(new_n207), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT73), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n304), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT34), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT74), .B(KEYINPUT34), .C1(new_n292), .C2(new_n295), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n319), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT75), .B1(new_n316), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n316), .A2(new_n324), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n316), .A2(KEYINPUT75), .A3(new_n324), .ZN(new_n328));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT0), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G57gat), .ZN(new_n331));
  INV_X1    g130(.A(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G141gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G148gat), .ZN(new_n335));
  INV_X1    g134(.A(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G141gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n335), .A2(new_n337), .B1(KEYINPUT2), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  NOR2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT78), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G155gat), .ZN(new_n343));
  INV_X1    g142(.A(G162gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n338), .ZN(new_n349));
  XNOR2_X1  g148(.A(G141gat), .B(G148gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(G155gat), .B2(G162gat), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n349), .B(KEYINPUT78), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n233), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n223), .A2(KEYINPUT79), .A3(new_n232), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(KEYINPUT3), .A3(new_n353), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n356), .A2(new_n358), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n348), .A2(KEYINPUT3), .A3(new_n353), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT3), .B1(new_n348), .B2(new_n353), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n223), .A2(KEYINPUT79), .A3(new_n232), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT79), .B1(new_n223), .B2(new_n232), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(KEYINPUT80), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n348), .A2(new_n353), .ZN(new_n373));
  OR3_X1    g172(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n298), .A2(new_n354), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AND4_X1   g176(.A1(KEYINPUT5), .A2(new_n371), .A3(new_n372), .A4(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n359), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n375), .B1(new_n380), .B2(new_n354), .ZN(new_n381));
  INV_X1    g180(.A(new_n372), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n363), .A2(new_n370), .B1(new_n376), .B2(new_n374), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(new_n372), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n333), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  INV_X1    g186(.A(new_n383), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n361), .A2(new_n362), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT80), .B1(new_n366), .B2(new_n369), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n377), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n388), .B1(new_n391), .B2(new_n382), .ZN(new_n392));
  INV_X1    g191(.A(new_n333), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n384), .A2(KEYINPUT5), .A3(new_n372), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT86), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n386), .A2(new_n395), .A3(new_n398), .A4(new_n387), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n392), .A2(KEYINPUT6), .A3(new_n393), .A4(new_n394), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT81), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G197gat), .B(G204gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT22), .ZN(new_n405));
  INV_X1    g204(.A(G211gat), .ZN(new_n406));
  INV_X1    g205(.A(G218gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n404), .A3(new_n408), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(KEYINPUT76), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n415), .A3(new_n411), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(KEYINPUT29), .B2(new_n365), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n422), .A3(new_n416), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n354), .B1(new_n423), .B2(new_n355), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT29), .B1(new_n412), .B2(new_n413), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n373), .B1(new_n426), .B2(KEYINPUT3), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n418), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(G22gat), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n428), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n423), .A2(new_n355), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n420), .B(new_n418), .C1(new_n432), .C2(new_n354), .ZN(new_n433));
  INV_X1    g232(.A(G22gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT31), .ZN(new_n438));
  INV_X1    g237(.A(G50gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n430), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n431), .A2(new_n433), .A3(KEYINPUT82), .A4(new_n434), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(new_n440), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n435), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n443), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n441), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT77), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n422), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n297), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n290), .A2(new_n257), .A3(new_n453), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n417), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n417), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G8gat), .B(G36gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(G64gat), .ZN(new_n463));
  INV_X1    g262(.A(G92gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n465), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n461), .A2(KEYINPUT30), .A3(new_n465), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT87), .B(KEYINPUT35), .Z(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n450), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n327), .A2(new_n328), .A3(new_n403), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n308), .B1(new_n307), .B2(new_n207), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n313), .A2(KEYINPUT73), .A3(new_n314), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n303), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n323), .ZN(new_n478));
  INV_X1    g277(.A(new_n441), .ZN(new_n479));
  INV_X1    g278(.A(new_n449), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n448), .B1(new_n443), .B2(new_n445), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n303), .B(new_n324), .C1(new_n475), .C2(new_n476), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n402), .A2(new_n396), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT35), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n482), .B1(new_n485), .B2(new_n487), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n378), .A2(new_n385), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n469), .A2(new_n470), .B1(new_n393), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT84), .B1(new_n384), .B2(new_n372), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n391), .A2(new_n496), .A3(new_n382), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT39), .ZN(new_n498));
  INV_X1    g297(.A(new_n381), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(new_n372), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n384), .A2(KEYINPUT84), .A3(new_n372), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n496), .B1(new_n391), .B2(new_n382), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n333), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT39), .B1(new_n495), .B2(new_n497), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT85), .B1(new_n508), .B2(new_n393), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n502), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n494), .B1(new_n510), .B2(KEYINPUT40), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT40), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n512), .B(new_n502), .C1(new_n507), .C2(new_n509), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n461), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT38), .ZN(new_n517));
  INV_X1    g316(.A(new_n465), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n459), .A2(KEYINPUT37), .A3(new_n460), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n468), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n465), .B1(new_n461), .B2(new_n515), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n517), .B1(new_n522), .B2(new_n519), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n400), .A2(new_n402), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n482), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n492), .B1(new_n514), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n478), .A2(KEYINPUT36), .A3(new_n483), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n483), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n328), .A3(new_n478), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n528), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n490), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G15gat), .B(G22gat), .Z(new_n535));
  INV_X1    g334(.A(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(G1gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n537), .A2(new_n540), .A3(new_n546), .A4(new_n541), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n549));
  XOR2_X1   g348(.A(G43gat), .B(G50gat), .Z(new_n550));
  INV_X1    g349(.A(KEYINPUT15), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G29gat), .A2(G36gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT88), .Z(new_n554));
  NOR2_X1   g353(.A1(G29gat), .A2(G36gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n550), .A2(new_n551), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT17), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n558), .A2(new_n559), .ZN(new_n564));
  AOI211_X1 g363(.A(new_n551), .B(new_n550), .C1(new_n554), .C2(new_n557), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n567), .A3(new_n547), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n549), .A2(new_n562), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT91), .Z(new_n571));
  OAI211_X1 g370(.A(new_n545), .B(new_n547), .C1(new_n564), .C2(new_n565), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n572), .A4(new_n571), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n548), .A2(new_n561), .A3(new_n560), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(new_n572), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n571), .B(KEYINPUT13), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT11), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n237), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT12), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n586), .A2(new_n576), .A3(new_n580), .A4(new_n575), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G78gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n203), .A2(new_n591), .A3(KEYINPUT9), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G57gat), .B(G64gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n203), .A3(new_n591), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n599), .A2(new_n600), .B1(G71gat), .B2(G78gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  OAI22_X1  g402(.A1(new_n601), .A2(new_n602), .B1(new_n595), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n593), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT93), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n597), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n406), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n595), .A2(new_n603), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n606), .B2(KEYINPUT93), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n601), .A2(new_n602), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n596), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n548), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(G183gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n252), .A3(new_n548), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  NOR2_X1   g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n622), .A2(new_n625), .ZN(new_n627));
  OR3_X1    g426(.A1(new_n613), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n613), .B1(new_n626), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT94), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n560), .A2(new_n561), .ZN(new_n640));
  OR2_X1    g439(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n464), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(G106gat), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT8), .B1(new_n206), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G99gat), .B(G106gat), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT7), .ZN(new_n649));
  OAI211_X1 g448(.A(KEYINPUT95), .B(new_n649), .C1(new_n332), .C2(new_n464), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(KEYINPUT95), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT7), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n651), .A2(new_n653), .A3(G85gat), .A4(G92gat), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n646), .A2(new_n648), .A3(new_n650), .A4(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n654), .A2(new_n643), .A3(new_n645), .A4(new_n650), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n647), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n640), .A2(new_n659), .B1(KEYINPUT41), .B2(new_n633), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n562), .A2(new_n566), .A3(new_n658), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n639), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n637), .B1(new_n662), .B2(KEYINPUT97), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n638), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n660), .A2(new_n661), .A3(new_n639), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n631), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n630), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n656), .B2(new_n647), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n657), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n656), .A2(new_n677), .A3(new_n647), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n617), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n658), .A2(new_n608), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n658), .B2(new_n608), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n676), .B(new_n681), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n659), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n675), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n692));
  INV_X1    g491(.A(new_n675), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G204gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT102), .B(G176gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n696), .B(new_n697), .Z(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n691), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n693), .B1(new_n685), .B2(new_n687), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n702), .B2(new_n694), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AND4_X1   g504(.A1(new_n590), .A2(new_n672), .A3(new_n674), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n534), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n485), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n536), .ZN(G1324gat));
  INV_X1    g508(.A(new_n707), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT16), .B(G8gat), .Z(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n486), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT42), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT42), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n710), .A2(new_n486), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n716), .A2(KEYINPUT104), .A3(G8gat), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT104), .B1(new_n716), .B2(G8gat), .ZN(new_n718));
  OAI22_X1  g517(.A1(new_n714), .A2(new_n715), .B1(new_n717), .B2(new_n718), .ZN(G1325gat));
  NAND2_X1  g518(.A1(new_n532), .A2(new_n529), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n478), .A2(KEYINPUT36), .A3(new_n483), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G15gat), .B1(new_n707), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n532), .A2(G15gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n707), .B2(new_n724), .ZN(G1326gat));
  NOR2_X1   g524(.A1(new_n707), .A2(new_n482), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT43), .B(G22gat), .Z(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  AOI21_X1  g527(.A(new_n506), .B1(new_n505), .B2(new_n333), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n508), .A2(KEYINPUT85), .A3(new_n393), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n501), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n512), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n510), .A2(KEYINPUT40), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n494), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n493), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n393), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT81), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n401), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n397), .B2(new_n399), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n450), .B1(new_n739), .B2(new_n524), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n491), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  AOI22_X1  g540(.A1(new_n741), .A2(new_n722), .B1(new_n489), .B2(new_n474), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n670), .ZN(new_n743));
  INV_X1    g542(.A(new_n590), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(new_n630), .A3(new_n704), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n746), .A2(G29gat), .A3(new_n485), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n745), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT44), .B1(new_n742), .B2(new_n670), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n534), .A2(new_n752), .A3(new_n671), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G29gat), .B1(new_n755), .B2(new_n485), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n749), .A2(new_n756), .ZN(G1328gat));
  INV_X1    g556(.A(G36gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n754), .B2(new_n486), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n487), .A2(G36gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n534), .A2(new_n671), .A3(new_n745), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT46), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT105), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT105), .B1(new_n759), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1329gat));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n766), .A2(KEYINPUT106), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(KEYINPUT106), .ZN(new_n768));
  INV_X1    g567(.A(G43gat), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n754), .B2(new_n533), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n746), .A2(G43gat), .A3(new_n532), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n767), .B(new_n768), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n742), .A2(KEYINPUT44), .A3(new_n670), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n752), .B1(new_n534), .B2(new_n671), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n533), .B(new_n745), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G43gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n534), .A2(new_n671), .ZN(new_n777));
  OR4_X1    g576(.A1(G43gat), .A2(new_n777), .A3(new_n532), .A4(new_n750), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n776), .A2(KEYINPUT106), .A3(new_n766), .A4(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n772), .A2(new_n779), .ZN(G1330gat));
  INV_X1    g579(.A(KEYINPUT48), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n777), .A2(KEYINPUT107), .A3(new_n750), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n482), .A2(G50gat), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n439), .B1(new_n754), .B2(new_n450), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n786), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(KEYINPUT48), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1331gat));
  NAND4_X1  g590(.A1(new_n672), .A2(new_n744), .A3(new_n674), .A4(new_n704), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n742), .A2(new_n485), .A3(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(G57gat), .Z(G1332gat));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n742), .B2(new_n792), .ZN(new_n796));
  INV_X1    g595(.A(new_n792), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n534), .A2(KEYINPUT108), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n487), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT109), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n800), .A2(KEYINPUT109), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(KEYINPUT109), .ZN(new_n804));
  NOR2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n806), .ZN(G1333gat));
  NOR2_X1   g606(.A1(new_n722), .A2(new_n203), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n796), .A2(new_n798), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n532), .B(KEYINPUT110), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n534), .A2(new_n797), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n203), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n809), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n814), .A2(KEYINPUT50), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT50), .B1(new_n814), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(G1334gat));
  NAND3_X1  g618(.A1(new_n796), .A2(new_n798), .A3(new_n450), .ZN(new_n820));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(G78gat), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n820), .B(new_n821), .ZN(G1335gat));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n630), .A2(new_n590), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n777), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n743), .A2(KEYINPUT51), .A3(new_n824), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT113), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT113), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n641), .A2(new_n642), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n402), .A2(new_n704), .A3(new_n396), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n825), .A2(new_n705), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n751), .B2(new_n753), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n485), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n830), .A2(new_n832), .B1(new_n831), .B2(new_n837), .ZN(G1336gat));
  NOR2_X1   g637(.A1(new_n487), .A2(G92gat), .ZN(new_n839));
  INV_X1    g638(.A(new_n826), .ZN(new_n840));
  INV_X1    g639(.A(new_n827), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n704), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n464), .B1(new_n835), .B2(new_n486), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n839), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n705), .B(new_n847), .C1(new_n826), .C2(new_n827), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT52), .B1(new_n848), .B2(new_n843), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(G1337gat));
  OAI21_X1  g649(.A(G99gat), .B1(new_n836), .B2(new_n722), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n327), .A2(new_n206), .A3(new_n328), .A4(new_n704), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n830), .B2(new_n852), .ZN(G1338gat));
  NOR2_X1   g652(.A1(new_n482), .A2(G106gat), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n704), .B(new_n854), .C1(new_n840), .C2(new_n841), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n644), .B1(new_n835), .B2(new_n450), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n854), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n705), .B(new_n860), .C1(new_n826), .C2(new_n827), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT53), .B1(new_n861), .B2(new_n856), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(G1339gat));
  NAND3_X1  g662(.A1(new_n577), .A2(new_n572), .A3(new_n579), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT114), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n571), .B1(new_n569), .B2(new_n572), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n585), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n704), .A2(new_n589), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n698), .B1(new_n702), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n685), .A2(new_n687), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT101), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n693), .B1(new_n872), .B2(new_n688), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n871), .B2(new_n675), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(KEYINPUT55), .B(new_n870), .C1(new_n873), .C2(new_n874), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n590), .A3(new_n701), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n868), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n670), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n589), .A2(new_n867), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n877), .A2(new_n671), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n879), .A2(new_n701), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n630), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n672), .A2(new_n744), .A3(new_n674), .A4(new_n705), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n450), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n532), .A2(new_n485), .A3(new_n486), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT115), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G113gat), .B1(new_n897), .B2(new_n744), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n890), .A2(new_n485), .A3(new_n486), .ZN(new_n899));
  INV_X1    g698(.A(new_n484), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n590), .A2(new_n216), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT116), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n898), .B1(new_n901), .B2(new_n903), .ZN(G1340gat));
  OAI21_X1  g703(.A(new_n217), .B1(new_n901), .B2(new_n705), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n704), .A2(G120gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n897), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n905), .B(KEYINPUT117), .C1(new_n897), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1341gat));
  OAI21_X1  g710(.A(G127gat), .B1(new_n897), .B2(new_n631), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n630), .A2(new_n211), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n901), .B2(new_n913), .ZN(G1342gat));
  OAI21_X1  g713(.A(G134gat), .B1(new_n897), .B2(new_n670), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n901), .A2(G134gat), .A3(new_n670), .ZN(new_n916));
  NAND2_X1  g715(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g717(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n919));
  OAI211_X1 g718(.A(new_n915), .B(new_n918), .C1(new_n916), .C2(new_n919), .ZN(G1343gat));
  NOR2_X1   g719(.A1(new_n485), .A2(new_n486), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n722), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n482), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT119), .B(new_n870), .C1(new_n873), .C2(new_n874), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT55), .B1(new_n875), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n880), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n868), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n670), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n630), .B1(new_n930), .B2(new_n886), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n888), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n875), .A2(new_n926), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n876), .A3(new_n925), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n879), .A2(new_n590), .A3(new_n701), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n671), .B1(new_n937), .B2(new_n868), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n884), .A2(new_n885), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n631), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(KEYINPUT120), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n924), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n923), .B1(new_n890), .B2(new_n482), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n922), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n334), .B1(new_n944), .B2(new_n590), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n533), .A2(new_n482), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT121), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n590), .A2(new_n334), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT122), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n899), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT58), .B1(new_n945), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n922), .ZN(new_n953));
  INV_X1    g752(.A(new_n924), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n889), .B1(new_n940), .B2(KEYINPUT120), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n931), .A2(new_n932), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n887), .A2(new_n889), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT57), .B1(new_n958), .B2(new_n450), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n953), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G141gat), .B1(new_n960), .B2(new_n744), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT58), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n962), .A3(new_n950), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n952), .A2(new_n963), .ZN(G1344gat));
  AND2_X1   g763(.A1(new_n947), .A2(new_n899), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n336), .A3(new_n704), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT59), .B(new_n336), .C1(new_n944), .C2(new_n704), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n958), .A2(KEYINPUT57), .A3(new_n450), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n888), .B(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n482), .B1(new_n971), .B2(new_n940), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n972), .B2(KEYINPUT57), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n704), .A3(new_n953), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n968), .B1(new_n974), .B2(G148gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n966), .B1(new_n967), .B2(new_n975), .ZN(G1345gat));
  NAND3_X1  g775(.A1(new_n947), .A2(new_n630), .A3(new_n899), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  AOI21_X1  g777(.A(G155gat), .B1(new_n977), .B2(KEYINPUT124), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n631), .A2(new_n343), .ZN(new_n980));
  AOI22_X1  g779(.A1(new_n978), .A2(new_n979), .B1(new_n944), .B2(new_n980), .ZN(G1346gat));
  OAI21_X1  g780(.A(G162gat), .B1(new_n960), .B2(new_n670), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n344), .A3(new_n671), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1347gat));
  AOI21_X1  g783(.A(new_n487), .B1(new_n402), .B2(new_n396), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n810), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n891), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n987), .A2(new_n237), .A3(new_n744), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n890), .B1(new_n402), .B2(new_n396), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(new_n486), .A3(new_n900), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n590), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n991), .B2(new_n237), .ZN(G1348gat));
  NAND3_X1  g791(.A1(new_n990), .A2(new_n238), .A3(new_n704), .ZN(new_n993));
  OAI21_X1  g792(.A(G176gat), .B1(new_n987), .B2(new_n705), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1349gat));
  NOR3_X1   g794(.A1(new_n631), .A2(new_n266), .A3(new_n265), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n990), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT60), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n998), .A2(KEYINPUT125), .ZN(new_n999));
  OAI21_X1  g798(.A(G183gat), .B1(new_n987), .B2(new_n631), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n999), .B1(new_n997), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1350gat));
  NAND3_X1  g802(.A1(new_n990), .A2(new_n253), .A3(new_n671), .ZN(new_n1004));
  OAI21_X1  g803(.A(G190gat), .B1(new_n987), .B2(new_n670), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n1005), .A2(KEYINPUT61), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n1005), .A2(KEYINPUT61), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1351gat));
  NOR3_X1   g807(.A1(new_n533), .A2(new_n487), .A3(new_n482), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g809(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g810(.A(G197gat), .B1(new_n1011), .B2(new_n590), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n1014));
  OAI211_X1 g813(.A(new_n969), .B(new_n1014), .C1(new_n972), .C2(KEYINPUT57), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n722), .A2(new_n985), .ZN(new_n1017));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  INV_X1    g818(.A(new_n1019), .ZN(new_n1020));
  AND3_X1   g819(.A1(new_n1020), .A2(G197gat), .A3(new_n590), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1012), .B1(new_n1016), .B2(new_n1021), .ZN(G1352gat));
  NOR2_X1   g821(.A1(new_n705), .A2(G204gat), .ZN(new_n1023));
  INV_X1    g822(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g823(.A(KEYINPUT62), .B1(new_n1010), .B2(new_n1024), .ZN(new_n1025));
  OR3_X1    g824(.A1(new_n1010), .A2(KEYINPUT62), .A3(new_n1024), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1020), .A2(new_n704), .ZN(new_n1027));
  AOI21_X1  g826(.A(new_n1027), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1028));
  INV_X1    g827(.A(G204gat), .ZN(new_n1029));
  OAI211_X1 g828(.A(new_n1025), .B(new_n1026), .C1(new_n1028), .C2(new_n1029), .ZN(G1353gat));
  NAND3_X1  g829(.A1(new_n1011), .A2(new_n406), .A3(new_n630), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n973), .A2(new_n630), .A3(new_n1020), .ZN(new_n1032));
  AND3_X1   g831(.A1(new_n1032), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1033));
  AOI21_X1  g832(.A(KEYINPUT63), .B1(new_n1032), .B2(G211gat), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(G1354gat));
  AOI21_X1  g834(.A(G218gat), .B1(new_n1011), .B2(new_n671), .ZN(new_n1036));
  NOR3_X1   g835(.A1(new_n1019), .A2(new_n407), .A3(new_n670), .ZN(new_n1037));
  AOI21_X1  g836(.A(new_n1036), .B1(new_n1016), .B2(new_n1037), .ZN(G1355gat));
endmodule


