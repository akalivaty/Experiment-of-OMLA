//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n202));
  NAND2_X1  g001(.A1(G15gat), .A2(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT87), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  INV_X1    g006(.A(G22gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT87), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(new_n203), .ZN(new_n211));
  INV_X1    g010(.A(G1gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT16), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n206), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(G1gat), .B1(new_n206), .B2(new_n211), .ZN(new_n215));
  OAI21_X1  g014(.A(G8gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n206), .A2(new_n211), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n212), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n206), .A2(new_n211), .A3(new_n213), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT21), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT91), .ZN(new_n225));
  INV_X1    g024(.A(G57gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G64gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(G64gat), .ZN(new_n228));
  INV_X1    g027(.A(G64gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G71gat), .A2(G78gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G71gat), .A2(G78gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT92), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT92), .ZN(new_n236));
  INV_X1    g035(.A(new_n234), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(new_n232), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT9), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n231), .A2(new_n235), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n234), .B(new_n233), .C1(new_n242), .C2(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n222), .B(new_n223), .C1(new_n224), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n216), .A2(new_n221), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n244), .A2(new_n224), .ZN(new_n247));
  OAI21_X1  g046(.A(G183gat), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G231gat), .A2(G233gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n202), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  INV_X1    g054(.A(new_n202), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n244), .A2(new_n224), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n258), .B(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G127gat), .B(G155gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n254), .A2(new_n257), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n254), .B2(new_n257), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT37), .ZN(new_n268));
  OR3_X1    g067(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n269), .A2(new_n270), .B1(G169gat), .B2(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n272), .A2(KEYINPUT25), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT24), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n223), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n271), .A2(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n276), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n223), .A2(new_n275), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(KEYINPUT24), .A3(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n280), .C1(new_n272), .C2(new_n271), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(KEYINPUT28), .A3(new_n275), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n284), .A2(new_n223), .A3(KEYINPUT27), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(KEYINPUT66), .B2(G183gat), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n285), .A2(new_n287), .A3(G190gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n283), .B1(new_n288), .B2(KEYINPUT28), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT26), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n290), .B2(new_n291), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT26), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n289), .A2(new_n278), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT24), .B1(new_n276), .B2(KEYINPUT65), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n279), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n276), .A2(KEYINPUT65), .A3(KEYINPUT24), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n271), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT25), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n305), .B2(new_n302), .ZN(new_n306));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT22), .ZN(new_n308));
  NAND2_X1  g107(.A1(G211gat), .A2(G218gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n260), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT22), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n307), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n303), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n302), .B1(new_n301), .B2(new_n304), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT72), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n316), .B(KEYINPUT71), .Z(new_n325));
  OAI211_X1 g124(.A(new_n268), .B(new_n318), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n323), .A3(new_n325), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n317), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT37), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT38), .ZN(new_n331));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(new_n229), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(G92gat), .Z(new_n334));
  NAND4_X1  g133(.A1(new_n326), .A2(new_n330), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n334), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n318), .B(new_n337), .C1(new_n324), .C2(new_n325), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  INV_X1    g139(.A(G155gat), .ZN(new_n341));
  INV_X1    g140(.A(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G141gat), .B(G148gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT73), .B(KEYINPUT2), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n340), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n344), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n343), .B2(KEYINPUT2), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352));
  INV_X1    g151(.A(G120gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT67), .B1(new_n353), .B2(G113gat), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n351), .B(new_n352), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G127gat), .B(G134gat), .Z(new_n360));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(KEYINPUT1), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n359), .B2(new_n362), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n339), .B(new_n350), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n349), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT4), .B1(new_n368), .B2(new_n363), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(KEYINPUT5), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n350), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n363), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(KEYINPUT74), .A3(new_n369), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n372), .A2(new_n374), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n368), .B(new_n363), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n373), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n363), .B(KEYINPUT68), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n363), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n373), .A2(new_n339), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n378), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT5), .B(new_n382), .C1(new_n385), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n380), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G57gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G85gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n389), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n390), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n338), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT79), .B1(new_n336), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n404), .A2(new_n335), .A3(new_n405), .A4(new_n338), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n326), .A2(new_n334), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n325), .B1(new_n321), .B2(new_n323), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n306), .A2(new_n317), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(new_n268), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT80), .B(KEYINPUT38), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT38), .B1(new_n407), .B2(new_n411), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n402), .A2(new_n406), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n396), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n372), .A2(new_n378), .A3(new_n379), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n373), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(KEYINPUT39), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n395), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(KEYINPUT39), .C1(new_n373), .C2(new_n381), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT40), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT78), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT40), .A4(new_n422), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n417), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n334), .B1(new_n408), .B2(new_n409), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n338), .A2(new_n428), .A3(KEYINPUT30), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n430), .A3(new_n337), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n421), .A2(new_n422), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n435), .A2(KEYINPUT40), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(KEYINPUT77), .A3(new_n431), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n427), .A2(new_n434), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G228gat), .ZN(new_n439));
  INV_X1    g238(.A(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT3), .B1(new_n316), .B2(new_n304), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT29), .B1(new_n350), .B2(new_n375), .ZN(new_n443));
  OAI221_X1 g242(.A(new_n441), .B1(new_n350), .B2(new_n442), .C1(new_n325), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT75), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n314), .A2(new_n445), .A3(new_n307), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(new_n304), .C1(new_n316), .C2(new_n445), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n350), .B1(new_n447), .B2(new_n375), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n443), .A2(new_n316), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n448), .A2(new_n449), .B1(new_n439), .B2(new_n440), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n208), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n208), .A3(new_n450), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT31), .B(G50gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n451), .B2(KEYINPUT76), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n452), .A2(KEYINPUT76), .A3(new_n453), .A4(new_n457), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n416), .A2(new_n438), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  AND2_X1   g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n301), .A2(new_n383), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n364), .A2(new_n366), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n466), .A2(new_n300), .A3(new_n295), .A4(new_n281), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n468), .A2(KEYINPUT34), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(KEYINPUT34), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n467), .A3(new_n464), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT69), .ZN(new_n475));
  XOR2_X1   g274(.A(G15gat), .B(G43gat), .Z(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n472), .B(KEYINPUT32), .C1(new_n473), .C2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n472), .B2(new_n473), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n471), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n478), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n469), .A2(new_n470), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n463), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(KEYINPUT70), .A3(new_n485), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT70), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT36), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n432), .A2(new_n403), .ZN(new_n490));
  INV_X1    g289(.A(new_n461), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n486), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT81), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT35), .ZN(new_n495));
  INV_X1    g294(.A(new_n437), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT77), .B1(new_n429), .B2(new_n431), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n487), .A2(new_n488), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n403), .A3(new_n461), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n499), .A2(new_n403), .A3(new_n461), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n434), .A2(new_n437), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT81), .A4(new_n495), .ZN(new_n504));
  INV_X1    g303(.A(new_n482), .ZN(new_n505));
  INV_X1    g304(.A(new_n485), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n491), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT35), .B1(new_n508), .B2(new_n490), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n501), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT96), .B(G134gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT41), .ZN(new_n514));
  NAND2_X1  g313(.A1(G232gat), .A2(G233gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT95), .ZN(new_n516));
  XOR2_X1   g315(.A(G99gat), .B(G106gat), .Z(new_n517));
  INV_X1    g316(.A(G99gat), .ZN(new_n518));
  INV_X1    g317(.A(G106gat), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT8), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT98), .B(G85gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n517), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n517), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n528), .A2(new_n532), .A3(KEYINPUT97), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n526), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(G85gat), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n536), .A2(KEYINPUT98), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(KEYINPUT98), .ZN(new_n538));
  OAI22_X1  g337(.A1(new_n537), .A2(new_n538), .B1(new_n522), .B2(new_n521), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n531), .A2(new_n535), .A3(new_n539), .A4(new_n520), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n530), .A2(KEYINPUT100), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n529), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT100), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n531), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT85), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n547), .A2(G29gat), .A3(G36gat), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  INV_X1    g348(.A(G36gat), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT14), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n546), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT14), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n547), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT85), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT83), .ZN(new_n557));
  INV_X1    g356(.A(G43gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(G50gat), .ZN(new_n559));
  INV_X1    g358(.A(G50gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(G43gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(G43gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(G50gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT83), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(KEYINPUT15), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G29gat), .A2(G36gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT15), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(KEYINPUT84), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n556), .A2(new_n566), .A3(new_n567), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n554), .A3(new_n567), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n562), .A2(new_n573), .A3(KEYINPUT15), .A4(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT17), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n545), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n545), .A2(new_n575), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n514), .B(new_n516), .C1(new_n581), .C2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G162gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT17), .B1(new_n575), .B2(new_n576), .ZN(new_n588));
  AOI211_X1 g387(.A(KEYINPUT86), .B(new_n578), .C1(new_n572), .C2(new_n574), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n544), .B(new_n541), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n516), .A2(new_n514), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n516), .A2(new_n514), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n582), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n584), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n587), .B1(new_n584), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n513), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n584), .A2(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n586), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n584), .A2(new_n587), .A3(new_n593), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n512), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n222), .B1(new_n588), .B2(new_n589), .ZN(new_n602));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT88), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n246), .A2(new_n575), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(KEYINPUT90), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n602), .A2(KEYINPUT18), .A3(new_n604), .A4(new_n605), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n572), .A2(new_n216), .A3(new_n221), .A4(new_n574), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n604), .B(KEYINPUT13), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT89), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT89), .ZN(new_n615));
  AOI211_X1 g414(.A(new_n615), .B(new_n612), .C1(new_n605), .C2(new_n610), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n608), .A2(new_n609), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G169gat), .B(G197gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n607), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT90), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n609), .A3(new_n617), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n618), .A2(new_n627), .B1(new_n628), .B2(new_n624), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n244), .B1(new_n540), .B2(new_n530), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n545), .B2(new_n244), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT101), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(KEYINPUT102), .A3(new_n633), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(KEYINPUT103), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT102), .B1(new_n631), .B2(new_n633), .ZN(new_n640));
  INV_X1    g439(.A(new_n244), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n541), .B2(new_n544), .ZN(new_n642));
  INV_X1    g441(.A(new_n633), .ZN(new_n643));
  NOR4_X1   g442(.A1(new_n642), .A2(new_n635), .A3(new_n630), .A4(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n639), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n642), .B2(new_n630), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n545), .A2(KEYINPUT10), .A3(new_n641), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n643), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n291), .ZN(new_n652));
  INV_X1    g451(.A(G204gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n638), .A2(new_n645), .A3(new_n650), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n636), .A2(new_n637), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n633), .B1(new_n647), .B2(new_n648), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n629), .A2(new_n660), .ZN(new_n661));
  AND4_X1   g460(.A1(new_n267), .A2(new_n511), .A3(new_n601), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n404), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n496), .A2(new_n497), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n666), .B2(new_n219), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT104), .B(G8gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  MUX2_X1   g469(.A(KEYINPUT42), .B(new_n667), .S(new_n670), .Z(G1325gat));
  AOI21_X1  g470(.A(G15gat), .B1(new_n662), .B2(new_n499), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n489), .A2(new_n486), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n207), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n672), .B1(new_n662), .B2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n491), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n678), .B(new_n680), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n596), .A2(new_n600), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n511), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n267), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n661), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n549), .A3(new_n404), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n601), .B1(new_n493), .B2(new_n510), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n685), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n403), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n688), .A2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n686), .A2(new_n550), .A3(new_n665), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n695), .B2(new_n503), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  OAI21_X1  g500(.A(G43gat), .B1(new_n695), .B2(new_n673), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n686), .A2(new_n558), .A3(new_n499), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n675), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n693), .A2(new_n706), .A3(new_n694), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n707), .B2(G43gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n705), .B1(KEYINPUT47), .B2(new_n708), .ZN(G1330gat));
  NAND4_X1  g508(.A1(new_n693), .A2(KEYINPUT108), .A3(new_n491), .A4(new_n694), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n690), .A2(new_n491), .A3(new_n694), .A4(new_n692), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n713), .A3(G50gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n461), .A2(G50gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n686), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(KEYINPUT48), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n711), .A2(G50gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n717), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n714), .A2(new_n724), .A3(KEYINPUT48), .A4(new_n717), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(new_n723), .A3(new_n725), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n601), .A2(new_n267), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n606), .A2(new_n607), .ZN(new_n728));
  INV_X1    g527(.A(new_n616), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n611), .A2(new_n613), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n615), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n609), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n624), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n625), .A2(new_n626), .ZN(new_n734));
  INV_X1    g533(.A(new_n624), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n608), .A2(new_n609), .A3(new_n617), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n727), .A2(new_n738), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n511), .A2(new_n660), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n404), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g541(.A(new_n503), .B(KEYINPUT110), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT111), .Z(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n740), .A2(new_n750), .A3(new_n499), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n740), .A2(new_n706), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n750), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g553(.A1(new_n740), .A2(new_n491), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n267), .A2(new_n738), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n693), .A2(new_n660), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n524), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n403), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  INV_X1    g560(.A(new_n660), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n511), .A2(new_n682), .A3(new_n757), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n691), .A2(KEYINPUT51), .A3(new_n757), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n524), .B1(new_n767), .B2(new_n404), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n760), .A2(new_n761), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n761), .B1(new_n760), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1336gat));
  NOR2_X1   g570(.A1(new_n744), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n765), .B2(new_n766), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT51), .B1(new_n691), .B2(new_n757), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(KEYINPUT113), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n660), .B(new_n772), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n691), .A2(KEYINPUT51), .A3(new_n757), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT113), .B1(new_n780), .B2(new_n775), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n773), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(KEYINPUT114), .A3(new_n660), .A4(new_n772), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n523), .B1(new_n758), .B2(new_n503), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n779), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n523), .B1(new_n758), .B2(new_n744), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(new_n767), .B2(new_n772), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n758), .B2(new_n675), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n767), .A2(new_n518), .A3(new_n499), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1338gat));
  OAI21_X1  g593(.A(G106gat), .B1(new_n758), .B2(new_n461), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n765), .A2(new_n766), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n461), .A2(new_n762), .A3(G106gat), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT53), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n797), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(G1339gat));
  AOI21_X1  g602(.A(new_n604), .B1(new_n602), .B2(new_n605), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n611), .A2(new_n613), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n623), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n736), .B2(new_n737), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n647), .A2(new_n633), .A3(new_n648), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT54), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n658), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n649), .A2(new_n813), .A3(new_n643), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n654), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n809), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n655), .B1(new_n658), .B2(new_n813), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n656), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n732), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n734), .A3(new_n735), .A4(new_n608), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n806), .ZN(new_n825));
  AND4_X1   g624(.A1(new_n682), .A2(new_n808), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n818), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT55), .B1(new_n817), .B2(new_n818), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n738), .A3(new_n656), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n823), .A2(new_n660), .A3(new_n806), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n682), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n684), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n739), .A2(new_n762), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n403), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n507), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n743), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n355), .A3(new_n738), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n743), .A2(new_n403), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(new_n499), .A3(new_n461), .A4(new_n835), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n629), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(G1340gat));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n353), .A3(new_n660), .ZN(new_n845));
  OAI21_X1  g644(.A(G120gat), .B1(new_n842), .B2(new_n762), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1341gat));
  INV_X1    g646(.A(G127gat), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n842), .A2(new_n848), .A3(new_n684), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n839), .A2(new_n267), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n848), .ZN(G1342gat));
  NOR2_X1   g650(.A1(new_n838), .A2(G134gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n665), .A2(new_n601), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT56), .Z(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n842), .B2(new_n601), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1343gat));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n836), .B2(new_n461), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n831), .B1(new_n629), .B2(new_n820), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n601), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n808), .A2(new_n821), .A3(new_n682), .A4(new_n825), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n267), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n727), .A2(new_n738), .A3(new_n660), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT57), .B(new_n491), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n841), .A2(new_n673), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n629), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n675), .A2(new_n491), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n837), .B1(new_n872), .B2(KEYINPUT116), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(KEYINPUT116), .B2(new_n872), .ZN(new_n874));
  INV_X1    g673(.A(G141gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n744), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n870), .B1(new_n629), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT58), .ZN(G1344gat));
  AND2_X1   g677(.A1(new_n874), .A2(new_n744), .ZN(new_n879));
  AOI21_X1  g678(.A(G148gat), .B1(new_n879), .B2(new_n660), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n869), .B2(new_n762), .ZN(new_n882));
  INV_X1    g681(.A(new_n867), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n883), .B2(KEYINPUT117), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT119), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n863), .B2(new_n864), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n887), .A3(new_n491), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n858), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n835), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n491), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n865), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n762), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n884), .B(new_n894), .C1(KEYINPUT117), .C2(new_n883), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n882), .A2(new_n895), .ZN(new_n896));
  AOI22_X1  g695(.A1(KEYINPUT59), .A2(new_n880), .B1(new_n896), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g696(.A(G155gat), .B1(new_n879), .B2(new_n267), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n684), .A2(new_n341), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n868), .B2(new_n899), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n869), .B2(new_n601), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n874), .A2(new_n342), .A3(new_n853), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n665), .A2(new_n403), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT120), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(KEYINPUT120), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n835), .A2(new_n499), .A3(new_n461), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT121), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT121), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n629), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n743), .A2(new_n835), .A3(new_n403), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n508), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n290), .A3(new_n738), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n915), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n914), .B2(new_n660), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n911), .A2(new_n762), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g718(.A(G183gat), .B1(new_n911), .B2(new_n684), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n267), .A3(new_n282), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n275), .A3(new_n682), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  INV_X1    g724(.A(new_n911), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n682), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n927), .B2(G190gat), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT61), .B(new_n275), .C1(new_n926), .C2(new_n682), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n932), .B(new_n924), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1351gat));
  NAND3_X1  g733(.A1(new_n905), .A2(new_n675), .A3(new_n906), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n935), .B1(new_n889), .B2(new_n893), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n629), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n913), .A2(new_n871), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n738), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1352gat));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n653), .A3(new_n660), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n945));
  INV_X1    g744(.A(new_n935), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n894), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n944), .B(new_n945), .C1(new_n947), .C2(new_n653), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT123), .Z(G1353gat));
  NAND2_X1  g748(.A1(new_n889), .A2(new_n893), .ZN(new_n950));
  AND4_X1   g749(.A1(KEYINPUT124), .A2(new_n950), .A3(new_n267), .A4(new_n946), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT124), .B1(new_n936), .B2(new_n267), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n953), .A2(G211gat), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n950), .A2(new_n267), .A3(new_n946), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n936), .A2(KEYINPUT124), .A3(new_n267), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n961), .A2(G211gat), .A3(new_n957), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n955), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n939), .A2(new_n260), .A3(new_n267), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n958), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n958), .A2(new_n964), .A3(new_n968), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n939), .B2(new_n682), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT127), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n937), .A2(new_n310), .A3(new_n601), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


