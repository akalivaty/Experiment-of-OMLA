//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n211), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n202), .A2(new_n203), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n223), .B(new_n230), .C1(KEYINPUT1), .C2(new_n218), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n220), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n201), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n203), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  AOI21_X1  g0051(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1698), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n256), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(G1698), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(KEYINPUT69), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n252), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G274), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT68), .B(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n276), .B1(G226), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n270), .A2(new_n271), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT75), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n205), .A2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n228), .A2(KEYINPUT72), .A3(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT72), .B1(new_n228), .B2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT74), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n205), .A2(new_n298), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT73), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n300), .B1(new_n293), .B2(new_n295), .C1(new_n291), .C2(new_n292), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n287), .A2(new_n297), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT71), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n304), .A2(KEYINPUT70), .A3(new_n227), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT70), .B1(new_n304), .B2(new_n227), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n227), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n304), .A2(KEYINPUT70), .A3(new_n227), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(KEYINPUT71), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n302), .A2(new_n314), .B1(new_n201), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n307), .B2(new_n312), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n272), .A2(G20), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(G50), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n270), .A2(new_n282), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n285), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n322), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT79), .B1(new_n327), .B2(G190), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(G200), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT9), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT10), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n302), .A2(new_n314), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n316), .A2(new_n201), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n334), .A2(KEYINPUT9), .A3(new_n320), .A4(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n330), .A2(new_n332), .A3(new_n333), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n328), .A3(new_n329), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT9), .B1(new_n317), .B2(new_n320), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT10), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n326), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n262), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G226), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G1698), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n343), .B(new_n345), .C1(new_n263), .C2(new_n264), .ZN(new_n346));
  INV_X1    g0146(.A(G87), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n254), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n276), .B1(new_n350), .B2(new_n252), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT84), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n278), .A2(G232), .A3(new_n279), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT82), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT82), .A4(G232), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n351), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n352), .B1(new_n351), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n323), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n351), .A2(KEYINPUT83), .A3(new_n271), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n350), .A2(new_n252), .ZN(new_n362));
  INV_X1    g0162(.A(G41), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT68), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G41), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n272), .B(G274), .C1(new_n367), .C2(G45), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n357), .A2(new_n362), .A3(new_n271), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT83), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n360), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n292), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n313), .A2(new_n315), .A3(new_n319), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n292), .A2(new_n316), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n255), .A2(new_n228), .A3(new_n256), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT7), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n255), .A2(new_n379), .A3(new_n228), .A4(new_n256), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(G68), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n378), .A2(KEYINPUT81), .A3(G68), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(G58), .B(G68), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(KEYINPUT16), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n310), .A2(new_n311), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n381), .A2(new_n387), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n376), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT18), .B1(new_n372), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  INV_X1    g0195(.A(new_n357), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G223), .A2(G1698), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n344), .B2(G1698), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n348), .B1(new_n398), .B2(new_n260), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n368), .B1(new_n399), .B2(new_n278), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n396), .A2(new_n400), .A3(G190), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT84), .B1(new_n396), .B2(new_n400), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n351), .A2(new_n352), .A3(new_n357), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G200), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n374), .A2(new_n375), .ZN(new_n407));
  INV_X1    g0207(.A(new_n387), .ZN(new_n408));
  AOI211_X1 g0208(.A(new_n391), .B(new_n408), .C1(new_n383), .C2(new_n384), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n390), .A2(new_n391), .ZN(new_n410));
  INV_X1    g0210(.A(new_n389), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n407), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n395), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(G169), .B1(new_n402), .B2(new_n403), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n371), .A2(new_n361), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n413), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n405), .B1(new_n358), .B2(new_n359), .ZN(new_n420));
  INV_X1    g0220(.A(new_n401), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(new_n393), .A3(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n394), .A2(new_n414), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT78), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n315), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n272), .A2(KEYINPUT78), .A3(G13), .A4(G20), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n389), .A2(new_n429), .A3(new_n319), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(new_n259), .ZN(new_n431));
  INV_X1    g0231(.A(new_n429), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n259), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n291), .A2(new_n434), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n292), .A2(new_n295), .B1(new_n228), .B2(new_n259), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n411), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(G232), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n260), .A2(KEYINPUT76), .A3(G232), .A4(new_n342), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n260), .A2(new_n208), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G238), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n267), .B2(new_n268), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n252), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n276), .B1(G244), .B2(new_n281), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n445), .B1(new_n442), .B2(new_n443), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT69), .B1(new_n260), .B2(G1698), .ZN(new_n455));
  INV_X1    g0255(.A(new_n268), .ZN(new_n456));
  OAI21_X1  g0256(.A(G238), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n278), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n452), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT77), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n439), .B1(new_n461), .B2(new_n271), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n453), .A2(new_n460), .A3(new_n323), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(G77), .B1(new_n289), .B2(new_n290), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n307), .A3(new_n312), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n307), .A3(new_n312), .A4(new_n469), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n203), .A2(KEYINPUT12), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n429), .A2(new_n474), .B1(KEYINPUT12), .B2(new_n316), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n430), .A2(KEYINPUT12), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(G68), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G226), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G97), .ZN(new_n480));
  INV_X1    g0280(.A(G232), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n479), .B(new_n480), .C1(new_n265), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n252), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n276), .B1(G238), .B2(new_n281), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT13), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT13), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(G179), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n323), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT14), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n488), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n487), .B1(new_n483), .B2(new_n484), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n491), .B(G169), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n478), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n464), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n453), .A2(new_n460), .A3(G200), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n439), .ZN(new_n501));
  INV_X1    g0301(.A(G190), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n453), .B2(new_n460), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n473), .A2(new_n477), .ZN(new_n505));
  OAI21_X1  g0305(.A(G200), .B1(new_n493), .B2(new_n494), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n486), .A2(G190), .A3(new_n488), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AND4_X1   g0309(.A1(new_n341), .A2(new_n425), .A3(new_n499), .A4(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT5), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G41), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n274), .B2(KEYINPUT5), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n272), .A2(G45), .A3(G274), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n278), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n515), .A2(KEYINPUT86), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT86), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n367), .B2(new_n512), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n516), .A2(new_n278), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G250), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n252), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n272), .A2(G45), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n514), .B(new_n530), .C1(new_n274), .C2(KEYINPUT5), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G264), .A3(new_n278), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(G169), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n528), .A2(new_n532), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT86), .B1(new_n515), .B2(new_n517), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n520), .A2(new_n519), .A3(new_n521), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(G179), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT91), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n228), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n260), .A2(new_n544), .A3(new_n228), .A4(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n228), .A2(G107), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n547), .A2(new_n548), .B1(G20), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT89), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(KEYINPUT89), .A3(new_n548), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n546), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n546), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n411), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  AOI21_X1  g0360(.A(G107), .B1(new_n560), .B2(KEYINPUT90), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n316), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n560), .A2(KEYINPUT90), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n254), .A2(G1), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n316), .B(new_n565), .C1(new_n307), .C2(new_n312), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n566), .B2(G107), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n540), .A2(new_n541), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n534), .A2(new_n539), .A3(KEYINPUT91), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n559), .A2(new_n567), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n523), .A2(new_n533), .A3(G190), .ZN(new_n572));
  AOI21_X1  g0372(.A(G200), .B1(new_n535), .B2(new_n538), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n568), .A2(new_n569), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n529), .A2(G250), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT87), .B1(new_n252), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT87), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n278), .A2(new_n578), .A3(G250), .A4(new_n529), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n516), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G238), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n549), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n252), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n405), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n580), .A2(new_n584), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(G190), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n565), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n318), .A2(G87), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n260), .A2(new_n228), .A3(G68), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n228), .B1(new_n480), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G87), .B2(new_n209), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT72), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n254), .B2(G20), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n207), .B1(new_n595), .B2(new_n288), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n590), .B(new_n593), .C1(KEYINPUT19), .C2(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n411), .B1(new_n432), .B2(new_n434), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n580), .A2(new_n584), .A3(new_n271), .ZN(new_n600));
  AOI21_X1  g0400(.A(G169), .B1(new_n580), .B2(new_n584), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n434), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n313), .A2(new_n315), .A3(new_n588), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n587), .A2(new_n599), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G97), .A2(G107), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT6), .B1(new_n209), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n208), .A2(KEYINPUT6), .A3(G97), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n610), .A2(new_n228), .B1(new_n259), .B2(new_n295), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n378), .A2(G107), .A3(new_n380), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n411), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n318), .A2(G97), .A3(new_n588), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n316), .A2(new_n207), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n252), .B1(new_n520), .B2(new_n530), .ZN(new_n617));
  AOI22_X1  g0417(.A1(G257), .A2(new_n617), .B1(new_n536), .B2(new_n537), .ZN(new_n618));
  OAI211_X1 g0418(.A(G244), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT4), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(KEYINPUT85), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n260), .A2(G244), .A3(new_n342), .A4(new_n621), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n620), .A2(KEYINPUT85), .B1(G33), .B2(G283), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n623), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n252), .ZN(new_n628));
  AOI21_X1  g0428(.A(G200), .B1(new_n618), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n531), .A2(G257), .A3(new_n278), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n502), .A2(new_n628), .A3(new_n538), .A4(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n616), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n628), .A2(new_n538), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n323), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n628), .A2(new_n538), .A3(new_n271), .A4(new_n630), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n606), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  OAI211_X1 g0439(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n640));
  OAI211_X1 g0440(.A(G257), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n255), .A2(G303), .A3(new_n256), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n252), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n531), .A2(G270), .A3(new_n278), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n639), .B1(new_n523), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n538), .A2(KEYINPUT88), .A3(new_n644), .A4(new_n645), .ZN(new_n648));
  AOI21_X1  g0448(.A(G20), .B1(G33), .B2(G283), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(G33), .B2(new_n207), .ZN(new_n650));
  INV_X1    g0450(.A(G116), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G20), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n308), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT20), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n650), .A2(new_n308), .A3(KEYINPUT20), .A4(new_n652), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n655), .A2(new_n656), .B1(new_n432), .B2(new_n651), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n389), .A2(G116), .A3(new_n429), .A4(new_n588), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n323), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n647), .A2(new_n648), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT21), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n647), .A2(new_n659), .A3(KEYINPUT21), .A4(new_n648), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n538), .A2(G179), .A3(new_n644), .A4(new_n645), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n658), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n662), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n647), .A2(new_n648), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G190), .ZN(new_n670));
  INV_X1    g0470(.A(new_n666), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n647), .A2(G200), .A3(new_n648), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n575), .A2(new_n638), .A3(new_n668), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n511), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT92), .ZN(G372));
  AND3_X1   g0476(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n393), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT17), .B1(new_n422), .B2(new_n393), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n498), .A2(new_n679), .A3(new_n508), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n372), .A2(new_n393), .A3(KEYINPUT18), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n418), .B1(new_n417), .B2(new_n413), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n337), .A2(new_n340), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n326), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n559), .B(new_n567), .C1(new_n572), .C2(new_n573), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n606), .A2(new_n632), .A3(new_n687), .A4(new_n637), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT93), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n570), .A2(new_n540), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n570), .B2(new_n540), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n688), .B1(new_n692), .B2(new_n668), .ZN(new_n693));
  INV_X1    g0493(.A(new_n601), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n580), .A2(new_n584), .A3(new_n271), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n605), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT26), .B1(new_n697), .B2(new_n606), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n580), .A2(new_n584), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G200), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n580), .A2(new_n584), .A3(G190), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n598), .A3(new_n589), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT26), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n703), .A2(new_n637), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n696), .B1(new_n698), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n693), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n686), .B1(new_n511), .B2(new_n707), .ZN(G369));
  AOI22_X1  g0508(.A1(new_n660), .A2(new_n661), .B1(new_n666), .B2(new_n665), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n673), .A2(new_n663), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n272), .A2(new_n228), .A3(G13), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n666), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n668), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n570), .A2(new_n716), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n575), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n568), .A2(new_n569), .A3(new_n716), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n662), .A2(new_n663), .A3(new_n667), .ZN(new_n728));
  INV_X1    g0528(.A(new_n716), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(new_n575), .A3(new_n722), .ZN(new_n732));
  INV_X1    g0532(.A(new_n691), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n570), .A2(new_n540), .A3(new_n689), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n729), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n727), .A2(new_n737), .ZN(G399));
  INV_X1    g0538(.A(new_n221), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n367), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(G1), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n225), .B2(new_n741), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  AND4_X1   g0546(.A1(new_n687), .A2(new_n606), .A3(new_n632), .A4(new_n637), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n523), .A2(new_n533), .A3(new_n271), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n323), .B1(new_n535), .B2(new_n538), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n541), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n569), .A3(new_n570), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n663), .A3(new_n709), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  OR4_X1    g0553(.A1(KEYINPUT96), .A2(new_n703), .A3(new_n637), .A4(new_n704), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n697), .A2(new_n606), .A3(KEYINPUT26), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n704), .B1(new_n703), .B2(new_n637), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT96), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n753), .A2(new_n696), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n746), .B1(new_n758), .B2(new_n729), .ZN(new_n759));
  INV_X1    g0559(.A(G330), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n618), .A2(new_n586), .A3(new_n535), .A4(new_n628), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n664), .ZN(new_n763));
  INV_X1    g0563(.A(new_n633), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n699), .A2(new_n533), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n764), .A2(new_n665), .A3(KEYINPUT30), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(G179), .B1(new_n535), .B2(new_n538), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n586), .A2(KEYINPUT95), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT95), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n699), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n767), .A2(new_n633), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n763), .B(new_n766), .C1(new_n669), .C2(new_n771), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n772), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n773));
  AOI21_X1  g0573(.A(KEYINPUT31), .B1(new_n772), .B2(new_n716), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n710), .A2(new_n575), .A3(new_n638), .A4(new_n729), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n760), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n747), .B1(new_n735), .B2(new_n728), .ZN(new_n778));
  INV_X1    g0578(.A(new_n696), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n755), .B2(new_n756), .ZN(new_n780));
  AOI211_X1 g0580(.A(KEYINPUT29), .B(new_n716), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n759), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n745), .B1(new_n782), .B2(G1), .ZN(G364));
  INV_X1    g0583(.A(new_n720), .ZN(new_n784));
  INV_X1    g0584(.A(G13), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n272), .B1(new_n786), .B2(G45), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n740), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G330), .B2(new_n719), .ZN(new_n791));
  INV_X1    g0591(.A(new_n789), .ZN(new_n792));
  INV_X1    g0592(.A(new_n260), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n739), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n651), .B2(new_n739), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n250), .A2(new_n275), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n739), .A2(new_n260), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G45), .B2(new_n225), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n227), .B1(G20), .B2(new_n323), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n792), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT97), .ZN(new_n806));
  INV_X1    g0606(.A(new_n803), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n228), .A2(G190), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G179), .A2(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT100), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT100), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n405), .A2(G179), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n808), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT99), .Z(new_n818));
  AOI22_X1  g0618(.A1(new_n815), .A2(G329), .B1(new_n818), .B2(G283), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT101), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n228), .A2(new_n502), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n271), .A2(G200), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n808), .A2(new_n822), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G322), .A2(new_n824), .B1(new_n826), .B2(G311), .ZN(new_n827));
  INV_X1    g0627(.A(G303), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n821), .A2(new_n816), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n271), .A2(new_n405), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n808), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT33), .B(G317), .Z(new_n832));
  OAI221_X1 g0632(.A(new_n827), .B1(new_n828), .B2(new_n829), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n228), .B1(new_n809), .B2(G190), .ZN(new_n834));
  INV_X1    g0634(.A(G294), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n821), .A2(new_n830), .ZN(new_n836));
  INV_X1    g0636(.A(G326), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n793), .B1(new_n834), .B2(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n820), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n823), .B(KEYINPUT98), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT32), .ZN(new_n842));
  INV_X1    g0642(.A(G159), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n810), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n811), .A2(KEYINPUT32), .A3(G159), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n841), .A2(G58), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n836), .A2(new_n201), .B1(new_n829), .B2(new_n347), .ZN(new_n847));
  INV_X1    g0647(.A(new_n831), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(G68), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n260), .B1(new_n825), .B2(new_n259), .ZN(new_n850));
  INV_X1    g0650(.A(new_n834), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(G97), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n818), .A2(G107), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n846), .A2(new_n849), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n839), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n802), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n806), .B1(new_n807), .B2(new_n855), .C1(new_n719), .C2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n791), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G396));
  OAI221_X1 g0659(.A(new_n260), .B1(new_n834), .B2(new_n202), .C1(new_n201), .C2(new_n829), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n818), .A2(G68), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(G132), .C2(new_n815), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n825), .A2(new_n843), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n836), .A2(new_n865), .B1(new_n831), .B2(new_n293), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(new_n841), .C2(G143), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n863), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(G283), .A2(new_n848), .B1(new_n826), .B2(G116), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n815), .A2(G311), .B1(KEYINPUT102), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n793), .B1(new_n836), .B2(new_n828), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n208), .A2(new_n829), .B1(new_n823), .B2(new_n835), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n873), .B(new_n874), .C1(G97), .C2(new_n851), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n871), .A2(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n818), .A2(G87), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n872), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n807), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n803), .A2(new_n800), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n792), .B(new_n879), .C1(new_n259), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n461), .A2(new_n271), .ZN(new_n882));
  AND4_X1   g0682(.A1(new_n463), .A2(new_n882), .A3(new_n438), .A4(new_n729), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n438), .A2(new_n716), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n501), .B2(new_n503), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n464), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n881), .B1(new_n801), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n729), .B1(new_n693), .B2(new_n706), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OR3_X1    g0689(.A1(new_n889), .A2(KEYINPUT103), .A3(new_n886), .ZN(new_n890));
  INV_X1    g0690(.A(new_n777), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n885), .A2(new_n464), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n462), .A2(new_n463), .A3(new_n729), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n886), .B(new_n729), .C1(new_n693), .C2(new_n706), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n792), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n891), .B1(new_n890), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n887), .B1(new_n899), .B2(new_n900), .ZN(G384));
  NOR2_X1   g0701(.A1(new_n786), .A2(new_n272), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n772), .A2(new_n716), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT31), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n772), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(new_n674), .C2(new_n716), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n510), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT106), .Z(new_n909));
  NAND2_X1  g0709(.A1(new_n385), .A2(new_n387), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n391), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n408), .B1(new_n383), .B2(new_n384), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n313), .B1(new_n912), .B2(KEYINPUT16), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n376), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n914), .A2(new_n714), .B1(new_n413), .B2(new_n406), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n372), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n417), .A2(new_n413), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n422), .A2(new_n393), .ZN(new_n919));
  INV_X1    g0719(.A(new_n714), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n413), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n918), .A2(new_n919), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n914), .A2(new_n714), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n424), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n924), .A2(KEYINPUT38), .A3(new_n926), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n478), .A2(new_n716), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n508), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n497), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n478), .B(new_n729), .C1(new_n492), .C2(new_n496), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n892), .A2(new_n893), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n907), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n907), .A2(new_n938), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT104), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n922), .B1(new_n921), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n944), .A2(new_n918), .A3(new_n919), .A4(new_n921), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n393), .A2(new_n714), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT37), .B1(new_n947), .B2(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n921), .B1(new_n683), .B2(new_n679), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n928), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n942), .A2(KEYINPUT105), .B1(new_n931), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n941), .B1(new_n953), .B2(new_n930), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n760), .B1(new_n909), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n909), .B2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n946), .B(new_n944), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n424), .A2(new_n947), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT38), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n924), .A2(KEYINPUT38), .A3(new_n926), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n936), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n931), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n683), .A2(new_n920), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n935), .A2(new_n936), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n896), .B2(new_n893), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n929), .A2(new_n931), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n510), .B1(new_n759), .B2(new_n781), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n686), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n971), .B(new_n973), .Z(new_n974));
  AOI21_X1  g0774(.A(new_n902), .B1(new_n956), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n956), .ZN(new_n976));
  INV_X1    g0776(.A(new_n610), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT35), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT35), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n978), .A2(G116), .A3(new_n229), .A4(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT36), .ZN(new_n981));
  OAI21_X1  g0781(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n246), .B1(new_n225), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(G1), .A3(new_n785), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n976), .A2(new_n981), .A3(new_n984), .ZN(G367));
  OAI211_X1 g0785(.A(new_n632), .B(new_n637), .C1(new_n616), .C2(new_n729), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n697), .A2(new_n716), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT42), .B1(new_n732), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n637), .B1(new_n986), .B2(new_n751), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT107), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n729), .A3(new_n994), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n989), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n990), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT108), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(KEYINPUT108), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n599), .A2(new_n729), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n779), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n703), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n998), .B(new_n999), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n727), .A2(new_n988), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1003), .B1(new_n998), .B2(new_n999), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1006), .ZN(new_n1010));
  OR3_X1    g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n740), .B(KEYINPUT41), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n737), .A2(new_n989), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT44), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n732), .A2(new_n736), .A3(new_n988), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT45), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n727), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1022), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n727), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1024), .A2(new_n1016), .A3(new_n1025), .A4(new_n1020), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n723), .A2(new_n730), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n726), .B2(new_n730), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(new_n720), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1023), .A2(new_n782), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1013), .B1(new_n1030), .B2(new_n782), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1011), .B(new_n1012), .C1(new_n788), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n241), .A2(new_n797), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n803), .B(new_n802), .C1(new_n739), .C2(new_n603), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n792), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n836), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(G143), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n834), .A2(new_n203), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G150), .B2(new_n824), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1037), .B1(new_n1040), .B2(KEYINPUT113), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(KEYINPUT113), .B2(new_n1040), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT114), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n817), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G77), .A2(new_n1045), .B1(new_n811), .B2(G137), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n202), .B2(new_n829), .C1(new_n843), .C2(new_n831), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n793), .B(new_n1047), .C1(G50), .C2(new_n826), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1043), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT115), .Z(new_n1050));
  INV_X1    g0850(.A(new_n829), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT46), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n829), .B2(new_n651), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(new_n835), .C2(new_n831), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT111), .ZN(new_n1056));
  INV_X1    g0856(.A(G317), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n793), .B1(new_n810), .B2(new_n1057), .C1(new_n207), .C2(new_n817), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1060));
  INV_X1    g0860(.A(G311), .ZN(new_n1061));
  INV_X1    g0861(.A(G283), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n836), .A2(new_n1061), .B1(new_n825), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G107), .B2(new_n851), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1060), .B(new_n1064), .C1(new_n828), .C2(new_n840), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1056), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1050), .A2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(KEYINPUT47), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n803), .B1(new_n1067), .B2(KEYINPUT47), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1035), .B1(new_n856), .B2(new_n1002), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1032), .A2(new_n1070), .ZN(G387));
  NAND2_X1  g0871(.A1(new_n1029), .A2(new_n788), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n742), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n794), .A2(new_n1073), .B1(new_n208), .B2(new_n739), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n238), .A2(new_n275), .ZN(new_n1075));
  AOI21_X1  g0875(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n373), .A2(new_n201), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n742), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n797), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1074), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n792), .B1(new_n1082), .B2(new_n804), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n793), .B1(new_n811), .B2(G150), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n848), .A2(new_n373), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n851), .A2(new_n603), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n826), .A2(G68), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n829), .A2(new_n259), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G159), .B2(new_n1036), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n201), .B2(new_n823), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1088), .B(new_n1091), .C1(G97), .C2(new_n818), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G311), .A2(new_n848), .B1(new_n826), .B2(G303), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1036), .A2(G322), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n840), .C2(new_n1057), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1096), .A2(KEYINPUT48), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(KEYINPUT48), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1051), .A2(G294), .B1(new_n851), .B2(G283), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT49), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n793), .B1(new_n810), .B2(new_n837), .C1(new_n651), .C2(new_n817), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1101), .B2(KEYINPUT49), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1092), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1083), .B1(new_n1105), .B2(new_n807), .C1(new_n725), .C2(new_n856), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1029), .A2(new_n782), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n740), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1029), .A2(new_n782), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1072), .B(new_n1106), .C1(new_n1108), .C2(new_n1109), .ZN(G393));
  NAND2_X1  g0910(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n787), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1112), .B2(new_n1111), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n1107), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n740), .A3(new_n1030), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n797), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n804), .B1(new_n207), .B2(new_n221), .C1(new_n245), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n789), .ZN(new_n1119));
  INV_X1    g0919(.A(G143), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n825), .A2(new_n292), .B1(new_n810), .B2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n260), .B1(new_n834), .B2(new_n259), .C1(new_n203), .C2(new_n829), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(G50), .C2(new_n848), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G150), .A2(new_n1036), .B1(new_n824), .B2(G159), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n818), .A2(G87), .B1(new_n1124), .B2(KEYINPUT51), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(KEYINPUT51), .C2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n793), .B1(new_n829), .B2(new_n1062), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G322), .B2(new_n811), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n853), .A2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT118), .Z(new_n1130));
  OAI22_X1  g0930(.A1(new_n836), .A2(new_n1057), .B1(new_n823), .B2(new_n1061), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT52), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n848), .A2(G303), .B1(new_n851), .B2(G116), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(new_n1134), .B1(G294), .B2(new_n826), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n1135), .C1(new_n1134), .C2(new_n1133), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1126), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1119), .B1(new_n1137), .B2(new_n803), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n988), .B2(new_n856), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1114), .A2(new_n1116), .A3(new_n1139), .ZN(G390));
  OAI21_X1  g0940(.A(new_n893), .B1(new_n888), .B2(new_n894), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n967), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n962), .A2(new_n964), .B1(new_n1143), .B2(new_n936), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n967), .B(KEYINPUT120), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n758), .A2(new_n729), .A3(new_n892), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n893), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n936), .B1(new_n960), .B2(new_n961), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n907), .A2(G330), .A3(new_n886), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1150), .A2(new_n967), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1144), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n777), .A2(new_n886), .A3(new_n1142), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n931), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT39), .B1(new_n952), .B2(new_n931), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1154), .A2(new_n1155), .B1(new_n968), .B2(new_n963), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n963), .B1(new_n952), .B2(new_n931), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1146), .A2(new_n893), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n1145), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1153), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1150), .A2(new_n1145), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1161), .A2(new_n1158), .A3(new_n1153), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1150), .A2(new_n967), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n1153), .B1(new_n893), .B2(new_n896), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n510), .A2(new_n777), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n972), .A2(new_n1166), .A3(new_n686), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1152), .A2(new_n1160), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1151), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1156), .A2(new_n1159), .A3(new_n1153), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1142), .B1(new_n777), .B2(new_n886), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1141), .B1(new_n1151), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1161), .A2(new_n1158), .A3(new_n1153), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1167), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1169), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1168), .A2(new_n740), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n880), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n789), .B1(new_n373), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n801), .B1(new_n962), .B2(new_n964), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT54), .B(G143), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n260), .B1(new_n834), .B2(new_n843), .C1(new_n825), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(G132), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n823), .A2(new_n1182), .B1(new_n817), .B2(new_n201), .ZN(new_n1183));
  INV_X1    g0983(.A(G128), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n836), .A2(new_n1184), .B1(new_n831), .B2(new_n865), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1181), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n829), .A2(new_n293), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT53), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1186), .B(new_n1188), .C1(new_n1189), .C2(new_n814), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n862), .B1(G294), .B2(new_n815), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n260), .B1(new_n1051), .B2(G87), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n831), .A2(new_n208), .B1(new_n825), .B2(new_n207), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G283), .B2(new_n1036), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n823), .A2(new_n651), .B1(new_n834), .B2(new_n259), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT121), .Z(new_n1197));
  OAI21_X1  g0997(.A(new_n1190), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1178), .B(new_n1179), .C1(new_n803), .C2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1152), .A2(new_n1160), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1200), .B2(new_n788), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1176), .A2(new_n1201), .ZN(G378));
  NAND2_X1  g1002(.A1(new_n321), .A2(new_n920), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n341), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n341), .A2(new_n1203), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1204), .A2(new_n1205), .A3(KEYINPUT123), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT123), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n971), .A2(G330), .A3(new_n954), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n952), .A2(new_n931), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT105), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n907), .B2(new_n938), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT40), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n760), .B1(new_n1217), .B2(new_n941), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(new_n971), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1212), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n937), .B1(new_n776), .B2(new_n775), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1215), .A2(new_n1221), .B1(new_n960), .B2(new_n961), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1222), .A2(KEYINPUT40), .B1(new_n932), .B2(new_n940), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n965), .B(new_n970), .C1(new_n1223), .C2(new_n760), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n971), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n1211), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1220), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1211), .A2(new_n800), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n789), .B1(G50), .B2(new_n1177), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n836), .A2(new_n651), .B1(new_n831), .B2(new_n207), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n793), .A2(new_n274), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1089), .A4(new_n1038), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n823), .A2(new_n208), .B1(new_n825), .B2(new_n434), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G58), .B2(new_n1045), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(new_n1062), .C2(new_n814), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT58), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G50), .B1(new_n254), .B2(new_n363), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1235), .A2(new_n1236), .B1(new_n1231), .B2(new_n1237), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n811), .C2(G124), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n836), .A2(new_n1189), .B1(new_n834), .B2(new_n293), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT122), .Z(new_n1241));
  OAI22_X1  g1041(.A1(new_n1184), .A2(new_n823), .B1(new_n829), .B2(new_n1180), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n831), .A2(new_n1182), .B1(new_n825), .B2(new_n865), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT59), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1239), .B1(new_n843), .B2(new_n817), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1238), .B1(new_n1236), .B2(new_n1235), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1229), .B1(new_n1248), .B2(new_n803), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1227), .A2(new_n788), .B1(new_n1228), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1167), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1175), .A2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1224), .A2(new_n1225), .A3(new_n1211), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1211), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1254));
  OAI211_X1 g1054(.A(KEYINPUT57), .B(new_n1252), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n740), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1252), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1256), .B2(new_n1257), .ZN(G375));
  NOR2_X1   g1058(.A1(new_n1174), .A2(new_n1013), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n788), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1145), .A2(new_n800), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n792), .B1(new_n203), .B2(new_n880), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n260), .B1(new_n834), .B2(new_n201), .C1(new_n202), .C2(new_n817), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n829), .A2(new_n843), .B1(new_n825), .B2(new_n293), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n836), .A2(new_n1182), .B1(new_n831), .B2(new_n1180), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n815), .A2(G128), .B1(G137), .B2(new_n841), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n815), .A2(G303), .B1(new_n818), .B2(G77), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1086), .B(new_n793), .C1(new_n207), .C2(new_n829), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n651), .A2(new_n831), .B1(new_n823), .B2(new_n1062), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n836), .A2(new_n835), .B1(new_n825), .B2(new_n208), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1268), .A2(new_n1269), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1263), .B(new_n1264), .C1(new_n807), .C2(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1262), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1261), .A2(new_n1277), .ZN(G381));
  NAND3_X1  g1078(.A1(new_n1176), .A2(new_n1201), .A3(KEYINPUT124), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT124), .B1(new_n1176), .B2(new_n1201), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n1250), .C1(new_n1257), .C2(new_n1256), .ZN(new_n1283));
  INV_X1    g1083(.A(G390), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OR3_X1    g1086(.A1(new_n1283), .A2(G387), .A3(new_n1286), .ZN(G407));
  OAI211_X1 g1087(.A(G407), .B(G213), .C1(G343), .C2(new_n1283), .ZN(G409));
  XNOR2_X1  g1088(.A(G393), .B(new_n858), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(G387), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1289), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1032), .B2(new_n1070), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1284), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1293), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT126), .B1(new_n1032), .B2(new_n1070), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1295), .B(G390), .C1(new_n1289), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G378), .B(new_n1250), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1013), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1300), .B(new_n1252), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n788), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1228), .A2(new_n1249), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G378), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1306), .A3(new_n1279), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1299), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n715), .A2(G213), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT60), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1260), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1165), .A2(KEYINPUT60), .A3(new_n1167), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(new_n740), .A3(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(KEYINPUT125), .B(new_n887), .C1(new_n899), .C2(new_n900), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1277), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G384), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1314), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1322));
  INV_X1    g1122(.A(G2897), .ZN(new_n1323));
  OAI22_X1  g1123(.A1(new_n1321), .A2(new_n1322), .B1(new_n1323), .B2(new_n1309), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1322), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1309), .A2(new_n1323), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1320), .A3(new_n1326), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1310), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1330), .B1(new_n1310), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1309), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1333), .B1(new_n1299), .B2(new_n1307), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1331), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1298), .A2(new_n1329), .A3(new_n1332), .A4(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1334), .A2(new_n1338), .A3(new_n1335), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT61), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1340), .B1(new_n1334), .B2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1338), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1339), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1337), .B1(new_n1344), .B2(new_n1298), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1282), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1346), .A2(new_n1347), .A3(new_n1299), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1347), .B1(new_n1346), .B2(new_n1299), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1348), .A2(new_n1349), .A3(new_n1335), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1346), .A2(new_n1299), .ZN(new_n1351));
  NOR3_X1   g1151(.A1(new_n1351), .A2(new_n1331), .A3(KEYINPUT127), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1298), .B1(new_n1350), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1351), .A2(KEYINPUT127), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1346), .A2(new_n1347), .A3(new_n1299), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1354), .A2(new_n1331), .A3(new_n1355), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1348), .B1(new_n1349), .B2(new_n1335), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1356), .A2(new_n1357), .A3(new_n1294), .A4(new_n1297), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1353), .A2(new_n1358), .ZN(G402));
endmodule


