

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717;

  AND2_X1 U368 ( .A1(n384), .A2(n383), .ZN(n382) );
  INV_X2 U369 ( .A(G953), .ZN(n707) );
  AND2_X1 U370 ( .A1(n588), .A2(n618), .ZN(n556) );
  XNOR2_X1 U371 ( .A(n556), .B(n555), .ZN(n714) );
  NAND2_X2 U372 ( .A1(n373), .A2(n354), .ZN(n415) );
  NAND2_X1 U373 ( .A1(n361), .A2(n646), .ZN(n573) );
  XNOR2_X1 U374 ( .A(n526), .B(KEYINPUT31), .ZN(n622) );
  XNOR2_X1 U375 ( .A(n513), .B(n514), .ZN(n712) );
  NOR2_X1 U376 ( .A1(n622), .A2(n609), .ZN(n532) );
  NOR2_X1 U377 ( .A1(n523), .A2(n516), .ZN(n508) );
  NOR2_X1 U378 ( .A1(n648), .A2(n634), .ZN(n420) );
  XNOR2_X1 U379 ( .A(KEYINPUT64), .B(KEYINPUT22), .ZN(n499) );
  XNOR2_X1 U380 ( .A(KEYINPUT85), .B(KEYINPUT33), .ZN(n507) );
  NOR2_X2 U381 ( .A1(n549), .A2(n558), .ZN(n568) );
  XNOR2_X2 U382 ( .A(n702), .B(G146), .ZN(n460) );
  XNOR2_X2 U383 ( .A(G119), .B(KEYINPUT3), .ZN(n449) );
  XNOR2_X2 U384 ( .A(n688), .B(n355), .ZN(n669) );
  XNOR2_X2 U385 ( .A(n357), .B(n358), .ZN(n688) );
  XNOR2_X2 U386 ( .A(n371), .B(KEYINPUT103), .ZN(n711) );
  INV_X1 U387 ( .A(n627), .ZN(n589) );
  NOR2_X1 U388 ( .A1(n672), .A2(G902), .ZN(n416) );
  NAND2_X1 U389 ( .A1(G237), .A2(G234), .ZN(n494) );
  XNOR2_X1 U390 ( .A(n560), .B(KEYINPUT6), .ZN(n572) );
  XNOR2_X1 U391 ( .A(n460), .B(n459), .ZN(n597) );
  XNOR2_X1 U392 ( .A(n431), .B(n368), .ZN(n435) );
  XNOR2_X1 U393 ( .A(n466), .B(KEYINPUT65), .ZN(n467) );
  INV_X1 U394 ( .A(KEYINPUT1), .ZN(n466) );
  XNOR2_X1 U395 ( .A(n553), .B(n552), .ZN(n588) );
  XNOR2_X1 U396 ( .A(n551), .B(KEYINPUT69), .ZN(n552) );
  XNOR2_X1 U397 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U398 ( .A(n413), .B(n412), .ZN(n679) );
  XNOR2_X1 U399 ( .A(n477), .B(n474), .ZN(n412) );
  XNOR2_X1 U400 ( .A(n414), .B(n470), .ZN(n413) );
  INV_X1 U401 ( .A(G475), .ZN(n421) );
  AND2_X2 U402 ( .A1(n423), .A2(n415), .ZN(n362) );
  XNOR2_X1 U403 ( .A(G116), .B(G137), .ZN(n452) );
  XNOR2_X1 U404 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n582) );
  XNOR2_X1 U405 ( .A(n537), .B(KEYINPUT84), .ZN(n380) );
  INV_X1 U406 ( .A(KEYINPUT44), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n432), .B(n349), .ZN(n368) );
  XNOR2_X1 U408 ( .A(KEYINPUT98), .B(G134), .ZN(n427) );
  INV_X1 U409 ( .A(n463), .ZN(n403) );
  XNOR2_X1 U410 ( .A(G107), .B(G110), .ZN(n461) );
  XOR2_X1 U411 ( .A(G101), .B(G104), .Z(n462) );
  XNOR2_X1 U412 ( .A(n367), .B(G478), .ZN(n522) );
  OR2_X1 U413 ( .A1(n595), .A2(G902), .ZN(n367) );
  XNOR2_X1 U414 ( .A(n451), .B(n450), .ZN(n483) );
  XNOR2_X1 U415 ( .A(G101), .B(KEYINPUT68), .ZN(n450) );
  XNOR2_X1 U416 ( .A(n429), .B(G116), .ZN(n484) );
  XNOR2_X1 U417 ( .A(G107), .B(G122), .ZN(n429) );
  XNOR2_X1 U418 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n437) );
  XNOR2_X1 U419 ( .A(n473), .B(n476), .ZN(n414) );
  XNOR2_X1 U420 ( .A(G140), .B(KEYINPUT96), .ZN(n471) );
  XNOR2_X1 U421 ( .A(G122), .B(G143), .ZN(n469) );
  XNOR2_X1 U422 ( .A(n364), .B(G113), .ZN(n482) );
  INV_X1 U423 ( .A(G104), .ZN(n364) );
  NOR2_X1 U424 ( .A1(n593), .A2(n628), .ZN(n594) );
  XNOR2_X1 U425 ( .A(n460), .B(n400), .ZN(n672) );
  XNOR2_X1 U426 ( .A(n402), .B(n401), .ZN(n400) );
  XNOR2_X1 U427 ( .A(n426), .B(n465), .ZN(n401) );
  XNOR2_X1 U428 ( .A(n464), .B(n403), .ZN(n402) );
  XNOR2_X1 U429 ( .A(n356), .B(n489), .ZN(n355) );
  XNOR2_X1 U430 ( .A(n360), .B(n487), .ZN(n356) );
  OR2_X2 U431 ( .A1(n631), .A2(n347), .ZN(n523) );
  NAND2_X1 U432 ( .A1(n511), .A2(n510), .ZN(n648) );
  XNOR2_X1 U433 ( .A(n557), .B(KEYINPUT106), .ZN(n649) );
  INV_X1 U434 ( .A(n584), .ZN(n411) );
  INV_X1 U435 ( .A(n370), .ZN(n410) );
  BUF_X1 U436 ( .A(n573), .Z(n370) );
  XNOR2_X1 U437 ( .A(n572), .B(KEYINPUT76), .ZN(n501) );
  INV_X1 U438 ( .A(n572), .ZN(n516) );
  NAND2_X1 U439 ( .A1(n362), .A2(G472), .ZN(n599) );
  XNOR2_X1 U440 ( .A(n597), .B(KEYINPUT62), .ZN(n598) );
  INV_X1 U441 ( .A(n706), .ZN(n405) );
  XNOR2_X1 U442 ( .A(n482), .B(n359), .ZN(n358) );
  XNOR2_X1 U443 ( .A(n483), .B(n484), .ZN(n357) );
  XNOR2_X1 U444 ( .A(KEYINPUT16), .B(G110), .ZN(n359) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n644) );
  XNOR2_X1 U446 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n388) );
  NOR2_X1 U447 ( .A1(n649), .A2(n648), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n554), .B(KEYINPUT40), .ZN(n555) );
  INV_X1 U449 ( .A(KEYINPUT105), .ZN(n554) );
  NAND2_X1 U450 ( .A1(n407), .A2(n399), .ZN(n624) );
  XNOR2_X1 U451 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X1 U452 ( .A(KEYINPUT109), .B(KEYINPUT36), .ZN(n408) );
  NAND2_X1 U453 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U454 ( .A(KEYINPUT120), .ZN(n374) );
  XNOR2_X1 U455 ( .A(n378), .B(n377), .ZN(n376) );
  NOR2_X1 U456 ( .A1(n687), .A2(n682), .ZN(n683) );
  INV_X1 U457 ( .A(KEYINPUT56), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n395) );
  OR2_X2 U459 ( .A1(n633), .A2(n634), .ZN(n347) );
  AND2_X1 U460 ( .A1(n581), .A2(n381), .ZN(n348) );
  XNOR2_X1 U461 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n349) );
  NOR2_X1 U462 ( .A1(n586), .A2(n361), .ZN(n350) );
  XOR2_X1 U463 ( .A(G128), .B(G110), .Z(n351) );
  OR2_X1 U464 ( .A1(n631), .A2(n398), .ZN(n352) );
  AND2_X1 U465 ( .A1(n712), .A2(n379), .ZN(n353) );
  OR2_X1 U466 ( .A1(n592), .A2(n593), .ZN(n354) );
  XNOR2_X1 U467 ( .A(G902), .B(KEYINPUT15), .ZN(n592) );
  XNOR2_X1 U468 ( .A(KEYINPUT86), .B(n596), .ZN(n687) );
  INV_X1 U469 ( .A(n687), .ZN(n394) );
  XNOR2_X2 U470 ( .A(n457), .B(KEYINPUT4), .ZN(n487) );
  XNOR2_X1 U471 ( .A(n486), .B(n485), .ZN(n360) );
  XNOR2_X1 U472 ( .A(n361), .B(n550), .ZN(n645) );
  AND2_X1 U473 ( .A1(n566), .A2(n361), .ZN(n567) );
  XNOR2_X2 U474 ( .A(n492), .B(n491), .ZN(n361) );
  NAND2_X1 U475 ( .A1(n362), .A2(G478), .ZN(n378) );
  NAND2_X1 U476 ( .A1(n362), .A2(G210), .ZN(n397) );
  NAND2_X1 U477 ( .A1(n362), .A2(G469), .ZN(n675) );
  NAND2_X1 U478 ( .A1(n362), .A2(G217), .ZN(n685) );
  NAND2_X1 U479 ( .A1(n695), .A2(n417), .ZN(n369) );
  XNOR2_X2 U480 ( .A(n540), .B(KEYINPUT45), .ZN(n695) );
  XNOR2_X2 U481 ( .A(n458), .B(n487), .ZN(n702) );
  NOR2_X2 U482 ( .A1(n560), .A2(n523), .ZN(n524) );
  NAND2_X1 U483 ( .A1(n568), .A2(n645), .ZN(n553) );
  XNOR2_X1 U484 ( .A(n436), .B(n351), .ZN(n366) );
  XNOR2_X1 U485 ( .A(n363), .B(n499), .ZN(n503) );
  NAND2_X1 U486 ( .A1(n418), .A2(n420), .ZN(n363) );
  XNOR2_X1 U487 ( .A(n369), .B(KEYINPUT78), .ZN(n373) );
  XNOR2_X1 U488 ( .A(n372), .B(n509), .ZN(n512) );
  NOR2_X1 U489 ( .A1(n365), .A2(n603), .ZN(n533) );
  NOR2_X1 U490 ( .A1(n532), .A2(n650), .ZN(n365) );
  NAND2_X1 U491 ( .A1(n517), .A2(n500), .ZN(n371) );
  XNOR2_X1 U492 ( .A(n366), .B(n439), .ZN(n442) );
  NOR2_X2 U493 ( .A1(n600), .A2(n687), .ZN(n602) );
  NAND2_X1 U494 ( .A1(n654), .A2(n525), .ZN(n372) );
  NAND2_X1 U495 ( .A1(n537), .A2(n712), .ZN(n515) );
  XNOR2_X1 U496 ( .A(n375), .B(n374), .ZN(G63) );
  NAND2_X1 U497 ( .A1(n376), .A2(n394), .ZN(n375) );
  INV_X1 U498 ( .A(n595), .ZN(n377) );
  NAND2_X1 U499 ( .A1(n575), .A2(n498), .ZN(n419) );
  XNOR2_X2 U500 ( .A(n573), .B(KEYINPUT19), .ZN(n575) );
  NOR2_X2 U501 ( .A1(n711), .A2(n390), .ZN(n537) );
  NAND2_X1 U502 ( .A1(n380), .A2(n353), .ZN(n538) );
  NAND2_X2 U503 ( .A1(n382), .A2(n348), .ZN(n387) );
  NAND2_X1 U504 ( .A1(n714), .A2(n425), .ZN(n381) );
  NAND2_X1 U505 ( .A1(n716), .A2(n425), .ZN(n383) );
  NAND2_X1 U506 ( .A1(n386), .A2(n385), .ZN(n384) );
  NOR2_X1 U507 ( .A1(n714), .A2(n425), .ZN(n385) );
  INV_X1 U508 ( .A(n716), .ZN(n386) );
  XNOR2_X2 U509 ( .A(n387), .B(n582), .ZN(n591) );
  XNOR2_X1 U510 ( .A(n390), .B(n713), .ZN(G21) );
  XNOR2_X1 U511 ( .A(n506), .B(n505), .ZN(n390) );
  XNOR2_X2 U512 ( .A(n528), .B(G472), .ZN(n560) );
  NAND2_X1 U513 ( .A1(n391), .A2(n525), .ZN(n526) );
  XNOR2_X1 U514 ( .A(n524), .B(KEYINPUT94), .ZN(n391) );
  NOR2_X1 U515 ( .A1(n641), .A2(n391), .ZN(n642) );
  XNOR2_X1 U516 ( .A(n393), .B(n392), .ZN(G51) );
  NAND2_X1 U517 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U518 ( .A(n671), .ZN(n396) );
  INV_X1 U519 ( .A(n633), .ZN(n398) );
  NOR2_X2 U520 ( .A1(n503), .A2(n399), .ZN(n517) );
  INV_X1 U521 ( .A(n631), .ZN(n399) );
  NOR2_X2 U522 ( .A1(n406), .A2(n592), .ZN(n417) );
  NAND2_X1 U523 ( .A1(n695), .A2(n404), .ZN(n628) );
  INV_X1 U524 ( .A(n406), .ZN(n404) );
  XNOR2_X1 U525 ( .A(n406), .B(n405), .ZN(n708) );
  NAND2_X2 U526 ( .A1(n591), .A2(n590), .ZN(n406) );
  NAND2_X1 U527 ( .A1(n422), .A2(n415), .ZN(n681) );
  XNOR2_X2 U528 ( .A(n416), .B(G469), .ZN(n563) );
  INV_X1 U529 ( .A(n529), .ZN(n418) );
  XNOR2_X2 U530 ( .A(n419), .B(KEYINPUT0), .ZN(n529) );
  NOR2_X1 U531 ( .A1(n594), .A2(n421), .ZN(n422) );
  INV_X1 U532 ( .A(n594), .ZN(n423) );
  XNOR2_X2 U533 ( .A(n563), .B(n467), .ZN(n631) );
  NOR2_X2 U534 ( .A1(n490), .A2(n669), .ZN(n492) );
  INV_X1 U535 ( .A(n457), .ZN(n430) );
  XOR2_X2 U536 ( .A(KEYINPUT66), .B(G131), .Z(n468) );
  AND2_X1 U537 ( .A1(G224), .A2(n707), .ZN(n424) );
  XOR2_X1 U538 ( .A(KEYINPUT46), .B(KEYINPUT81), .Z(n425) );
  AND2_X1 U539 ( .A1(G227), .A2(n707), .ZN(n426) );
  XNOR2_X1 U540 ( .A(n488), .B(n424), .ZN(n489) );
  INV_X1 U541 ( .A(G472), .ZN(n527) );
  NOR2_X1 U542 ( .A1(n350), .A2(n589), .ZN(n590) );
  XNOR2_X1 U543 ( .A(n669), .B(n670), .ZN(n671) );
  XNOR2_X1 U544 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U545 ( .A(n504), .B(KEYINPUT75), .ZN(n505) );
  INV_X1 U546 ( .A(KEYINPUT63), .ZN(n601) );
  XOR2_X1 U547 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n428) );
  XNOR2_X1 U548 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X2 U549 ( .A(G143), .B(G128), .ZN(n457) );
  XNOR2_X1 U550 ( .A(n484), .B(n430), .ZN(n431) );
  NAND2_X1 U551 ( .A1(G234), .A2(n707), .ZN(n433) );
  XOR2_X1 U552 ( .A(KEYINPUT8), .B(n433), .Z(n440) );
  NAND2_X1 U553 ( .A1(G217), .A2(n440), .ZN(n434) );
  XOR2_X1 U554 ( .A(n435), .B(n434), .Z(n595) );
  XOR2_X1 U555 ( .A(G137), .B(G140), .Z(n463) );
  XOR2_X1 U556 ( .A(G146), .B(G125), .Z(n488) );
  XNOR2_X1 U557 ( .A(n488), .B(KEYINPUT10), .ZN(n470) );
  XNOR2_X1 U558 ( .A(n463), .B(n470), .ZN(n701) );
  XOR2_X1 U559 ( .A(KEYINPUT23), .B(G119), .Z(n436) );
  XOR2_X1 U560 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n438) );
  XNOR2_X1 U561 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U562 ( .A1(G221), .A2(n440), .ZN(n441) );
  XNOR2_X1 U563 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U564 ( .A(n701), .B(n443), .ZN(n684) );
  NOR2_X1 U565 ( .A1(n684), .A2(G902), .ZN(n448) );
  NAND2_X1 U566 ( .A1(n592), .A2(G234), .ZN(n444) );
  XNOR2_X1 U567 ( .A(n444), .B(KEYINPUT20), .ZN(n480) );
  NAND2_X1 U568 ( .A1(G217), .A2(n480), .ZN(n446) );
  INV_X1 U569 ( .A(KEYINPUT25), .ZN(n445) );
  XNOR2_X2 U570 ( .A(n448), .B(n447), .ZN(n633) );
  INV_X1 U571 ( .A(n449), .ZN(n451) );
  XOR2_X1 U572 ( .A(KEYINPUT5), .B(G113), .Z(n453) );
  XNOR2_X1 U573 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U574 ( .A(n483), .B(n454), .Z(n456) );
  NOR2_X1 U575 ( .A1(G953), .A2(G237), .ZN(n475) );
  NAND2_X1 U576 ( .A1(n475), .A2(G210), .ZN(n455) );
  XNOR2_X1 U577 ( .A(n456), .B(n455), .ZN(n459) );
  XNOR2_X2 U578 ( .A(n468), .B(G134), .ZN(n458) );
  NOR2_X2 U579 ( .A1(n597), .A2(G902), .ZN(n528) );
  AND2_X1 U580 ( .A1(n633), .A2(n560), .ZN(n500) );
  XNOR2_X1 U581 ( .A(KEYINPUT71), .B(KEYINPUT89), .ZN(n465) );
  XNOR2_X1 U582 ( .A(n462), .B(n461), .ZN(n464) );
  INV_X1 U583 ( .A(n522), .ZN(n511) );
  XNOR2_X1 U584 ( .A(n469), .B(n468), .ZN(n477) );
  XNOR2_X1 U585 ( .A(n482), .B(KEYINPUT95), .ZN(n474) );
  XOR2_X1 U586 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n472) );
  XNOR2_X1 U587 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U588 ( .A1(G214), .A2(n475), .ZN(n476) );
  NOR2_X1 U589 ( .A1(G902), .A2(n679), .ZN(n479) );
  XNOR2_X1 U590 ( .A(KEYINPUT13), .B(G475), .ZN(n478) );
  XNOR2_X1 U591 ( .A(n479), .B(n478), .ZN(n519) );
  INV_X1 U592 ( .A(n519), .ZN(n510) );
  NAND2_X1 U593 ( .A1(G221), .A2(n480), .ZN(n481) );
  XNOR2_X1 U594 ( .A(KEYINPUT21), .B(n481), .ZN(n634) );
  INV_X1 U595 ( .A(n592), .ZN(n490) );
  XOR2_X1 U596 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n486) );
  XNOR2_X1 U597 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n485) );
  OR2_X1 U598 ( .A1(G902), .A2(G237), .ZN(n493) );
  NAND2_X1 U599 ( .A1(G210), .A2(n493), .ZN(n491) );
  NAND2_X1 U600 ( .A1(G214), .A2(n493), .ZN(n646) );
  XNOR2_X1 U601 ( .A(n494), .B(KEYINPUT14), .ZN(n630) );
  XNOR2_X1 U602 ( .A(KEYINPUT87), .B(G898), .ZN(n693) );
  NAND2_X1 U603 ( .A1(n693), .A2(G953), .ZN(n495) );
  XOR2_X1 U604 ( .A(KEYINPUT88), .B(n495), .Z(n690) );
  NAND2_X1 U605 ( .A1(n690), .A2(G902), .ZN(n496) );
  NAND2_X1 U606 ( .A1(G952), .A2(n707), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n496), .A2(n542), .ZN(n497) );
  AND2_X1 U608 ( .A1(n630), .A2(n497), .ZN(n498) );
  OR2_X1 U609 ( .A1(n501), .A2(n352), .ZN(n502) );
  NOR2_X1 U610 ( .A1(n503), .A2(n502), .ZN(n506) );
  INV_X1 U611 ( .A(KEYINPUT32), .ZN(n504) );
  XOR2_X1 U612 ( .A(KEYINPUT80), .B(KEYINPUT35), .Z(n514) );
  XOR2_X1 U613 ( .A(KEYINPUT34), .B(KEYINPUT74), .Z(n509) );
  XNOR2_X1 U614 ( .A(n508), .B(n507), .ZN(n654) );
  INV_X1 U615 ( .A(n529), .ZN(n525) );
  NOR2_X1 U616 ( .A1(n511), .A2(n510), .ZN(n566) );
  NAND2_X1 U617 ( .A1(n512), .A2(n566), .ZN(n513) );
  NAND2_X1 U618 ( .A1(n515), .A2(KEYINPUT44), .ZN(n535) );
  NAND2_X1 U619 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U620 ( .A1(n633), .A2(n518), .ZN(n603) );
  XNOR2_X1 U621 ( .A(n519), .B(KEYINPUT97), .ZN(n521) );
  NOR2_X1 U622 ( .A1(n521), .A2(n522), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n520), .B(KEYINPUT101), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n522), .A2(n521), .ZN(n587) );
  NAND2_X1 U625 ( .A1(n569), .A2(n587), .ZN(n577) );
  INV_X1 U626 ( .A(n577), .ZN(n650) );
  NOR2_X2 U627 ( .A1(n563), .A2(n347), .ZN(n545) );
  XNOR2_X1 U628 ( .A(n528), .B(n527), .ZN(n640) );
  NOR2_X1 U629 ( .A1(n529), .A2(n640), .ZN(n530) );
  NAND2_X1 U630 ( .A1(n545), .A2(n530), .ZN(n531) );
  XNOR2_X1 U631 ( .A(KEYINPUT93), .B(n531), .ZN(n609) );
  XNOR2_X1 U632 ( .A(KEYINPUT102), .B(n533), .ZN(n534) );
  NAND2_X1 U633 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U634 ( .A(n536), .B(KEYINPUT83), .ZN(n539) );
  NAND2_X1 U635 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U636 ( .A1(G900), .A2(n707), .ZN(n541) );
  NAND2_X1 U637 ( .A1(n541), .A2(G902), .ZN(n543) );
  NAND2_X1 U638 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U639 ( .A1(n544), .A2(n630), .ZN(n558) );
  XNOR2_X1 U640 ( .A(n545), .B(KEYINPUT104), .ZN(n548) );
  NAND2_X1 U641 ( .A1(n640), .A2(n646), .ZN(n546) );
  XOR2_X1 U642 ( .A(KEYINPUT30), .B(n546), .Z(n547) );
  NAND2_X1 U643 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U644 ( .A(KEYINPUT38), .B(KEYINPUT70), .Z(n550) );
  XOR2_X1 U645 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n551) );
  INV_X1 U646 ( .A(n569), .ZN(n618) );
  XOR2_X1 U647 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n565) );
  NAND2_X1 U648 ( .A1(n646), .A2(n645), .ZN(n557) );
  NOR2_X1 U649 ( .A1(n634), .A2(n558), .ZN(n559) );
  NAND2_X1 U650 ( .A1(n633), .A2(n559), .ZN(n570) );
  NOR2_X1 U651 ( .A1(n560), .A2(n570), .ZN(n561) );
  XOR2_X1 U652 ( .A(KEYINPUT28), .B(n561), .Z(n562) );
  NOR2_X1 U653 ( .A1(n563), .A2(n562), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n644), .A2(n574), .ZN(n564) );
  XNOR2_X1 U655 ( .A(n565), .B(n564), .ZN(n716) );
  NAND2_X1 U656 ( .A1(n568), .A2(n567), .ZN(n615) );
  NOR2_X1 U657 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U658 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n615), .A2(n624), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U661 ( .A(n576), .B(KEYINPUT77), .ZN(n616) );
  NAND2_X1 U662 ( .A1(n577), .A2(n616), .ZN(n578) );
  XNOR2_X1 U663 ( .A(n578), .B(KEYINPUT47), .ZN(n579) );
  NOR2_X1 U664 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U665 ( .A1(n631), .A2(n646), .ZN(n583) );
  NOR2_X1 U666 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U667 ( .A(n585), .B(KEYINPUT43), .ZN(n586) );
  INV_X1 U668 ( .A(n587), .ZN(n621) );
  NAND2_X1 U669 ( .A1(n588), .A2(n621), .ZN(n627) );
  INV_X1 U670 ( .A(KEYINPUT2), .ZN(n593) );
  NOR2_X1 U671 ( .A1(G952), .A2(n707), .ZN(n596) );
  XNOR2_X1 U672 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U673 ( .A(n602), .B(n601), .ZN(G57) );
  XOR2_X1 U674 ( .A(G101), .B(n603), .Z(G3) );
  NAND2_X1 U675 ( .A1(n609), .A2(n618), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT110), .ZN(n605) );
  XNOR2_X1 U677 ( .A(G104), .B(n605), .ZN(G6) );
  XOR2_X1 U678 ( .A(KEYINPUT112), .B(KEYINPUT27), .Z(n607) );
  XNOR2_X1 U679 ( .A(G107), .B(KEYINPUT26), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n607), .B(n606), .ZN(n608) );
  XOR2_X1 U681 ( .A(KEYINPUT111), .B(n608), .Z(n611) );
  NAND2_X1 U682 ( .A1(n609), .A2(n621), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n611), .B(n610), .ZN(G9) );
  XOR2_X1 U684 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n613) );
  NAND2_X1 U685 ( .A1(n621), .A2(n616), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n614) );
  XOR2_X1 U687 ( .A(G128), .B(n614), .Z(G30) );
  XNOR2_X1 U688 ( .A(G143), .B(n615), .ZN(G45) );
  NAND2_X1 U689 ( .A1(n618), .A2(n616), .ZN(n617) );
  XNOR2_X1 U690 ( .A(n617), .B(G146), .ZN(G48) );
  NAND2_X1 U691 ( .A1(n622), .A2(n618), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n619), .B(KEYINPUT114), .ZN(n620) );
  XNOR2_X1 U693 ( .A(G113), .B(n620), .ZN(G15) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n623), .B(G116), .ZN(G18) );
  XNOR2_X1 U696 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(G125), .B(n626), .ZN(G27) );
  XNOR2_X1 U699 ( .A(G134), .B(n627), .ZN(G36) );
  XOR2_X1 U700 ( .A(G140), .B(n350), .Z(G42) );
  NAND2_X1 U701 ( .A1(n654), .A2(n644), .ZN(n666) );
  XNOR2_X1 U702 ( .A(KEYINPUT2), .B(KEYINPUT79), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(n663) );
  INV_X1 U704 ( .A(n630), .ZN(n660) );
  NAND2_X1 U705 ( .A1(n631), .A2(n347), .ZN(n632) );
  XNOR2_X1 U706 ( .A(KEYINPUT50), .B(n632), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n636) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n636), .B(n635), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U712 ( .A(KEYINPUT51), .B(n642), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n656) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n652) );
  NOR2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n651) );
  OR2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U718 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U719 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U720 ( .A(KEYINPUT52), .B(n657), .ZN(n658) );
  NAND2_X1 U721 ( .A1(n658), .A2(G952), .ZN(n659) );
  NOR2_X1 U722 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U723 ( .A(n661), .B(KEYINPUT117), .ZN(n662) );
  NAND2_X1 U724 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U725 ( .A1(G953), .A2(n664), .ZN(n665) );
  NAND2_X1 U726 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U727 ( .A(n667), .B(KEYINPUT53), .ZN(n668) );
  XOR2_X1 U728 ( .A(KEYINPUT118), .B(n668), .Z(G75) );
  XOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n670) );
  XNOR2_X1 U730 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n672), .B(KEYINPUT57), .ZN(n673) );
  XNOR2_X1 U732 ( .A(n674), .B(n673), .ZN(n676) );
  XNOR2_X1 U733 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U734 ( .A1(n687), .A2(n677), .ZN(G54) );
  INV_X1 U735 ( .A(KEYINPUT59), .ZN(n678) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U737 ( .A(KEYINPUT60), .B(n683), .ZN(G60) );
  XNOR2_X1 U738 ( .A(n684), .B(n685), .ZN(n686) );
  NOR2_X1 U739 ( .A1(n687), .A2(n686), .ZN(G66) );
  XOR2_X1 U740 ( .A(n688), .B(KEYINPUT123), .Z(n689) );
  NOR2_X1 U741 ( .A1(n690), .A2(n689), .ZN(n700) );
  NAND2_X1 U742 ( .A1(G953), .A2(G224), .ZN(n691) );
  XOR2_X1 U743 ( .A(KEYINPUT61), .B(n691), .Z(n692) );
  NOR2_X1 U744 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U745 ( .A(KEYINPUT121), .B(n694), .ZN(n698) );
  NAND2_X1 U746 ( .A1(n695), .A2(n707), .ZN(n696) );
  XNOR2_X1 U747 ( .A(KEYINPUT122), .B(n696), .ZN(n697) );
  NAND2_X1 U748 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U749 ( .A(n700), .B(n699), .ZN(G69) );
  XOR2_X1 U750 ( .A(n702), .B(n701), .Z(n706) );
  XOR2_X1 U751 ( .A(G227), .B(n706), .Z(n703) );
  NAND2_X1 U752 ( .A1(n703), .A2(G900), .ZN(n704) );
  NAND2_X1 U753 ( .A1(G953), .A2(n704), .ZN(n705) );
  XNOR2_X1 U754 ( .A(n705), .B(KEYINPUT124), .ZN(n710) );
  NAND2_X1 U755 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U756 ( .A1(n710), .A2(n709), .ZN(G72) );
  XOR2_X1 U757 ( .A(n711), .B(G110), .Z(G12) );
  XNOR2_X1 U758 ( .A(n712), .B(G122), .ZN(G24) );
  XNOR2_X1 U759 ( .A(G119), .B(KEYINPUT125), .ZN(n713) );
  XNOR2_X1 U760 ( .A(G131), .B(KEYINPUT127), .ZN(n715) );
  XNOR2_X1 U761 ( .A(n715), .B(n714), .ZN(G33) );
  XOR2_X1 U762 ( .A(G137), .B(n716), .Z(n717) );
  XNOR2_X1 U763 ( .A(KEYINPUT126), .B(n717), .ZN(G39) );
endmodule

