//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n203), .A2(new_n206), .A3(new_n204), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT14), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT15), .A4(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n214), .A2(new_n217), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT15), .B1(new_n221), .B2(new_n216), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n219), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n211), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT87), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n227), .A3(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n220), .B(new_n232), .C1(new_n222), .C2(new_n223), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n208), .B(new_n210), .C1(new_n231), .C2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n230), .A4(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n211), .A2(new_n224), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n211), .A2(new_n227), .A3(new_n224), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n227), .B1(new_n211), .B2(new_n224), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n230), .B(KEYINPUT13), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n242), .A3(KEYINPUT88), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n230), .A3(new_n235), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n250), .A2(new_n242), .A3(new_n236), .A4(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n242), .A3(new_n236), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n243), .A3(new_n249), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT36), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT26), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT26), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(G190gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT27), .B(G183gat), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n274), .A2(KEYINPUT28), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT28), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n270), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT25), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n267), .B2(new_n268), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT23), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n288), .A3(new_n264), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n280), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n267), .A3(new_n273), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n283), .A2(KEYINPUT64), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n293), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n291), .A2(new_n282), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  AND4_X1   g095(.A1(KEYINPUT25), .A2(new_n286), .A3(new_n288), .A4(new_n264), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n290), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n290), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n279), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  INV_X1    g104(.A(G120gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT1), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n307), .B(new_n309), .C1(new_n314), .C2(new_n306), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  AOI211_X1 g117(.A(new_n318), .B(new_n279), .C1(new_n301), .C2(new_n303), .ZN(new_n319));
  INV_X1    g118(.A(G227gat), .ZN(new_n320));
  INV_X1    g119(.A(G233gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n317), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n260), .B1(new_n324), .B2(KEYINPUT33), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n295), .A2(new_n297), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT66), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n295), .A2(new_n297), .A3(new_n296), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n302), .B1(new_n329), .B2(new_n290), .ZN(new_n330));
  INV_X1    g129(.A(new_n303), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n278), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n318), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n304), .A2(new_n316), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n322), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT33), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(KEYINPUT69), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G15gat), .B(G43gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n335), .B2(KEYINPUT32), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n323), .B1(new_n317), .B2(new_n319), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n343), .A2(KEYINPUT34), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(KEYINPUT34), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n335), .B(KEYINPUT32), .C1(new_n336), .C2(new_n340), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n342), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n259), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n341), .A2(new_n337), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT69), .B1(new_n335), .B2(new_n336), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n346), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT36), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G1gat), .B(G29gat), .Z(new_n358));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G141gat), .ZN(new_n367));
  INV_X1    g166(.A(G141gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G148gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n365), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(G155gat), .ZN(new_n372));
  INV_X1    g171(.A(G162gat), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT2), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n370), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n371), .B1(new_n370), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n364), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(new_n369), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(KEYINPUT73), .A3(new_n374), .ZN(new_n379));
  INV_X1    g178(.A(new_n371), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n370), .A2(new_n371), .A3(new_n374), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(KEYINPUT74), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n377), .A2(new_n383), .A3(new_n316), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n311), .A4(new_n315), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n385), .B2(KEYINPUT4), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n385), .A2(new_n391), .A3(KEYINPUT4), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n387), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n375), .A2(new_n376), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n316), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n377), .A2(KEYINPUT3), .A3(new_n383), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT75), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT75), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n377), .A2(new_n383), .A3(new_n404), .A4(KEYINPUT3), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT77), .B1(new_n397), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n405), .ZN(new_n408));
  INV_X1    g207(.A(new_n401), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT77), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n388), .B1(new_n394), .B2(new_n395), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n390), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n393), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n385), .A2(KEYINPUT4), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n385), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n410), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n423), .A2(KEYINPUT5), .A3(new_n388), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n363), .B1(new_n414), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n390), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n397), .A2(KEYINPUT77), .A3(new_n406), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n411), .B1(new_n410), .B2(new_n412), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n423), .A2(KEYINPUT5), .A3(new_n388), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n362), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(KEYINPUT6), .B(new_n363), .C1(new_n414), .C2(new_n424), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G197gat), .B(G204gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT22), .ZN(new_n437));
  INV_X1    g236(.A(G211gat), .ZN(new_n438));
  INV_X1    g237(.A(G218gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G211gat), .B(G218gat), .Z(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT70), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT70), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n445), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G226gat), .A2(G233gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n332), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n300), .A2(new_n278), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT72), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT72), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n455), .A3(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n447), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n449), .B(new_n278), .C1(new_n330), .C2(new_n331), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n452), .A2(new_n460), .A3(new_n448), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n447), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G8gat), .B(G36gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G64gat), .B(G92gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  NAND3_X1  g265(.A1(new_n458), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  INV_X1    g267(.A(new_n447), .ZN(new_n469));
  INV_X1    g268(.A(new_n450), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n448), .B1(new_n304), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n455), .B1(new_n452), .B2(new_n449), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT72), .B(new_n448), .C1(new_n300), .C2(new_n278), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n468), .B1(new_n475), .B2(new_n462), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n467), .A2(new_n476), .A3(KEYINPUT30), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n474), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n462), .B1(new_n478), .B2(new_n447), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n466), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n435), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n444), .A2(new_n460), .A3(new_n446), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n399), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n377), .A2(new_n383), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n400), .A2(new_n450), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n447), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(KEYINPUT80), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n447), .A2(new_n496), .A3(new_n489), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n399), .B1(new_n443), .B2(new_n470), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n381), .A2(new_n382), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G50gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n501), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n492), .B1(new_n488), .B2(new_n490), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G22gat), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n504), .B2(new_n507), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n484), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n509), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n505), .A2(new_n506), .A3(new_n502), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n503), .B1(new_n494), .B2(new_n501), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT81), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n350), .A2(new_n357), .B1(new_n483), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT39), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n423), .B2(new_n388), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT79), .B1(new_n385), .B2(KEYINPUT4), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(new_n417), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(new_n420), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n522), .B(new_n388), .C1(new_n526), .C2(new_n406), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n521), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n408), .A2(new_n409), .B1(new_n419), .B2(new_n421), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT82), .B1(new_n530), .B2(new_n387), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT39), .B1(new_n386), .B2(new_n388), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT83), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n534), .A3(new_n527), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n529), .A2(KEYINPUT40), .A3(new_n362), .A4(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n536), .A2(new_n425), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n477), .A2(new_n481), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n529), .A2(new_n362), .A3(new_n535), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT40), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n510), .A2(new_n511), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n478), .A2(new_n469), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n459), .A2(new_n461), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(new_n447), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT38), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT84), .B1(new_n479), .B2(new_n545), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n550));
  NOR4_X1   g349(.A1(new_n475), .A2(new_n462), .A3(new_n550), .A4(KEYINPUT37), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n468), .B(new_n548), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(new_n434), .A3(new_n433), .A4(new_n467), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT38), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n458), .A2(new_n545), .A3(new_n463), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n550), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n479), .A2(KEYINPUT84), .A3(new_n545), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n466), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT37), .B1(new_n475), .B2(new_n462), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n542), .B(new_n543), .C1(new_n553), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n520), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT85), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n348), .B2(new_n349), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n355), .A2(KEYINPUT85), .A3(new_n356), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n516), .A2(new_n517), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n433), .A2(new_n434), .B1(new_n481), .B2(new_n477), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n355), .A2(new_n543), .A3(new_n356), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT35), .B1(new_n570), .B2(new_n483), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n258), .B1(new_n562), .B2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT90), .B(G64gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(KEYINPUT89), .A2(G57gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  OR2_X1    g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n584));
  AND2_X1   g383(.A1(G57gat), .A2(G64gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n579), .B(new_n580), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(G127gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n588), .B(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G127gat), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n575), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n575), .A3(new_n594), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n211), .B1(new_n587), .B2(KEYINPUT21), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT91), .Z(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G155gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n599), .B(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n596), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n596), .B2(new_n597), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n611), .A2(new_n612), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  INV_X1    g414(.A(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(KEYINPUT8), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(KEYINPUT92), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT94), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n619), .B(new_n623), .C1(new_n620), .C2(KEYINPUT92), .ZN(new_n624));
  OAI211_X1 g423(.A(G85gat), .B(G92gat), .C1(new_n619), .C2(new_n620), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n622), .B2(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n618), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G99gat), .B(G106gat), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n631), .B(new_n618), .C1(new_n626), .C2(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n614), .B1(new_n634), .B2(new_n224), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n611), .A2(new_n612), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n633), .B1(new_n231), .B2(new_n234), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n635), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n610), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(new_n609), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n583), .A2(new_n586), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n633), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n587), .A2(new_n632), .A3(new_n630), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n633), .A2(KEYINPUT96), .A3(new_n646), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(KEYINPUT10), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n652), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n605), .A2(new_n645), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n573), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n435), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n482), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n209), .B2(new_n671), .ZN(new_n674));
  MUX2_X1   g473(.A(new_n673), .B(new_n674), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g474(.A1(new_n350), .A2(new_n357), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n668), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n564), .A2(new_n565), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(G15gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n677), .B1(new_n668), .B2(new_n680), .ZN(G1326gat));
  INV_X1    g480(.A(new_n519), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n668), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  AOI21_X1  g484(.A(new_n645), .B1(new_n562), .B2(new_n572), .ZN(new_n686));
  INV_X1    g485(.A(new_n605), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n665), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n258), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(G29gat), .A3(new_n435), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT97), .B(KEYINPUT45), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n562), .A2(new_n572), .ZN(new_n694));
  INV_X1    g493(.A(new_n645), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(KEYINPUT98), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n686), .A2(KEYINPUT98), .A3(KEYINPUT44), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n435), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n700), .A2(new_n701), .A3(new_n689), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n693), .B1(new_n702), .B2(new_n212), .ZN(G1328gat));
  NOR3_X1   g502(.A1(new_n690), .A2(G36gat), .A3(new_n482), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n700), .A2(new_n538), .A3(new_n689), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n213), .ZN(G1329gat));
  INV_X1    g506(.A(new_n676), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n698), .A2(new_n708), .A3(new_n699), .A4(new_n689), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(KEYINPUT47), .ZN(new_n712));
  NOR4_X1   g511(.A1(new_n679), .A2(G43gat), .A3(new_n645), .A4(new_n688), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(new_n573), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(KEYINPUT47), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT100), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n715), .B(new_n717), .ZN(G1330gat));
  NAND3_X1  g517(.A1(new_n700), .A2(new_n566), .A3(new_n689), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(G50gat), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n690), .A2(G50gat), .A3(new_n682), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n700), .A2(new_n519), .A3(new_n689), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n724), .B2(G50gat), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n720), .A2(new_n723), .B1(new_n725), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g525(.A1(new_n694), .A2(new_n258), .A3(new_n605), .A4(new_n645), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n664), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n435), .B(KEYINPUT101), .Z(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT102), .B(G57gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1332gat));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n733));
  INV_X1    g532(.A(G64gat), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n733), .B(new_n734), .C1(new_n728), .C2(new_n482), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n482), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n727), .A2(new_n664), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n728), .B2(new_n676), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n679), .A2(G71gat), .A3(new_n665), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n727), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g545(.A1(new_n728), .A2(new_n682), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g547(.A1(new_n605), .A2(new_n257), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n694), .A2(new_n695), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(KEYINPUT105), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n665), .A2(new_n435), .A3(G85gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n751), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n752), .B(new_n753), .C1(new_n756), .C2(KEYINPUT105), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n605), .A2(new_n665), .A3(new_n257), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n700), .A2(new_n701), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n759), .B2(new_n616), .ZN(G1336gat));
  NOR3_X1   g559(.A1(new_n665), .A2(new_n482), .A3(G92gat), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n752), .B(new_n761), .C1(new_n756), .C2(KEYINPUT105), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n698), .A2(new_n538), .A3(new_n699), .A4(new_n758), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G92gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n756), .A2(new_n761), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT106), .B1(new_n768), .B2(KEYINPUT52), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n764), .A2(G92gat), .B1(new_n756), .B2(new_n761), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n770), .A2(new_n771), .A3(new_n763), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n766), .B1(new_n769), .B2(new_n772), .ZN(G1337gat));
  NOR3_X1   g572(.A1(new_n679), .A2(G99gat), .A3(new_n665), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n752), .B(new_n774), .C1(new_n756), .C2(KEYINPUT105), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n700), .A2(new_n708), .A3(new_n758), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT107), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G99gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n776), .A2(KEYINPUT107), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(G1338gat));
  NOR3_X1   g579(.A1(new_n665), .A2(new_n543), .A3(G106gat), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n752), .B(new_n781), .C1(new_n756), .C2(KEYINPUT105), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n698), .A2(new_n566), .A3(new_n699), .A4(new_n758), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n698), .A2(new_n519), .A3(new_n699), .A4(new_n758), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n781), .B(KEYINPUT108), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n756), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT109), .B1(new_n791), .B2(KEYINPUT53), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n787), .A2(G106gat), .B1(new_n756), .B2(new_n789), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n794), .A3(new_n783), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n786), .B1(new_n792), .B2(new_n795), .ZN(G1339gat));
  XOR2_X1   g595(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n797));
  NAND4_X1  g596(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n656), .A2(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n661), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n662), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n798), .A2(new_n661), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(KEYINPUT55), .C1(new_n800), .C2(new_n799), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n253), .A2(new_n242), .A3(new_n236), .A4(new_n248), .ZN(new_n807));
  INV_X1    g606(.A(new_n241), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n229), .A2(new_n237), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n230), .B1(new_n229), .B2(new_n235), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n247), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND4_X1   g611(.A1(new_n644), .A2(new_n807), .A3(new_n642), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT111), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n658), .A2(new_n661), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n801), .B2(new_n802), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n806), .A4(new_n813), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n661), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n656), .A2(KEYINPUT54), .ZN(new_n821));
  INV_X1    g620(.A(new_n800), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n823), .A2(KEYINPUT55), .B1(new_n254), .B2(new_n256), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n807), .A2(new_n812), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n824), .A2(new_n817), .B1(new_n664), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n815), .B(new_n819), .C1(new_n826), .C2(new_n695), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n827), .A2(new_n687), .B1(new_n258), .B2(new_n667), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n729), .ZN(new_n829));
  INV_X1    g628(.A(new_n570), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n482), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n314), .A3(new_n257), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n819), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n803), .A2(new_n257), .A3(new_n662), .A4(new_n806), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n664), .A2(new_n825), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n695), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n687), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n667), .A2(new_n258), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n682), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n701), .A2(new_n482), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n841), .A2(new_n679), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n258), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n833), .A2(new_n844), .ZN(G1340gat));
  NAND2_X1  g644(.A1(new_n664), .A2(new_n306), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT113), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G120gat), .B1(new_n843), .B2(new_n665), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1341gat));
  NOR3_X1   g649(.A1(new_n843), .A2(new_n591), .A3(new_n687), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n687), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(G127gat), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT114), .B1(new_n831), .B2(new_n687), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(G1342gat));
  OR3_X1    g654(.A1(new_n831), .A2(G134gat), .A3(new_n645), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n843), .B2(new_n645), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(G1343gat));
  NOR3_X1   g659(.A1(new_n708), .A2(new_n543), .A3(new_n538), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n829), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n258), .A2(G141gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT58), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(KEYINPUT116), .A3(new_n864), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT57), .B1(new_n828), .B2(new_n682), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n840), .A2(new_n870), .A3(new_n566), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n708), .A2(new_n842), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT117), .B1(new_n873), .B2(new_n258), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G141gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n873), .A2(KEYINPUT117), .A3(new_n258), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n867), .B(new_n868), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G141gat), .B1(new_n873), .B2(new_n258), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n865), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(KEYINPUT115), .A3(KEYINPUT58), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT115), .B1(new_n879), .B2(KEYINPUT58), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(G1344gat));
  NOR3_X1   g681(.A1(new_n862), .A2(G148gat), .A3(new_n665), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT118), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n870), .B1(new_n840), .B2(new_n566), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n519), .A2(new_n870), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n817), .A2(new_n806), .A3(new_n813), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT119), .B1(new_n837), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n888), .C1(new_n826), .C2(new_n695), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n892), .A3(new_n687), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n887), .B1(new_n893), .B2(new_n839), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n664), .A3(new_n872), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n885), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n873), .A2(new_n665), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(KEYINPUT59), .A3(new_n366), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n884), .B1(new_n897), .B2(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(G155gat), .B1(new_n873), .B2(new_n687), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n863), .A2(new_n372), .A3(new_n605), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n863), .B2(new_n695), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n873), .A2(new_n373), .A3(new_n645), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1347gat));
  INV_X1    g705(.A(new_n841), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n907), .A2(new_n538), .A3(new_n678), .A4(new_n729), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n261), .A3(new_n258), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n828), .B2(new_n701), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n840), .A2(KEYINPUT120), .A3(new_n435), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n570), .A2(new_n482), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n257), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n909), .B1(new_n919), .B2(new_n261), .ZN(G1348gat));
  NOR3_X1   g719(.A1(new_n908), .A2(new_n262), .A3(new_n665), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n915), .A2(new_n665), .A3(new_n917), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n924), .A3(new_n262), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n922), .B2(G176gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(G1349gat));
  OAI21_X1  g726(.A(G183gat), .B1(new_n908), .B2(new_n687), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n929), .A2(new_n275), .A3(new_n605), .A4(new_n916), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT123), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n928), .A2(new_n930), .A3(new_n934), .A4(new_n931), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n928), .A2(new_n930), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n933), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n908), .B2(new_n645), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n918), .A2(new_n274), .A3(new_n695), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1351gat));
  NAND3_X1  g741(.A1(new_n676), .A2(new_n566), .A3(new_n538), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n911), .B2(new_n913), .ZN(new_n944));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n257), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n729), .A2(new_n676), .A3(new_n538), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n886), .A2(new_n894), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n257), .A2(G197gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n665), .A2(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT124), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n944), .A2(new_n951), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n893), .A2(new_n839), .ZN(new_n956));
  INV_X1    g755(.A(new_n887), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT57), .B1(new_n828), .B2(new_n543), .ZN(new_n959));
  INV_X1    g758(.A(new_n946), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n958), .A2(new_n664), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n944), .A2(new_n963), .A3(new_n950), .A4(new_n951), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n953), .A2(new_n955), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI22_X1  g766(.A1(new_n954), .A2(KEYINPUT62), .B1(G204gat), .B2(new_n961), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n968), .A2(KEYINPUT125), .A3(new_n953), .A4(new_n964), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n944), .A2(new_n438), .A3(new_n605), .ZN(new_n971));
  OR2_X1    g770(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n958), .A2(new_n605), .A3(new_n959), .A4(new_n960), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n975), .A2(new_n438), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n895), .A2(KEYINPUT126), .A3(new_n605), .A4(new_n960), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n977), .A2(new_n979), .A3(G211gat), .A4(new_n972), .ZN(new_n980));
  NAND2_X1  g779(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n971), .B1(new_n978), .B2(new_n982), .ZN(G1354gat));
  NAND3_X1  g782(.A1(new_n944), .A2(new_n439), .A3(new_n695), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n947), .A2(new_n695), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n985), .B2(new_n439), .ZN(G1355gat));
endmodule


