

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769;

  OR2_X1 U370 ( .A1(n680), .A2(n640), .ZN(n355) );
  NOR2_X1 U371 ( .A1(n572), .A2(n689), .ZN(n590) );
  XNOR2_X1 U372 ( .A(n575), .B(n574), .ZN(n713) );
  XNOR2_X1 U373 ( .A(n580), .B(KEYINPUT35), .ZN(n767) );
  XNOR2_X2 U374 ( .A(n469), .B(n468), .ZN(n554) );
  NOR2_X2 U375 ( .A1(n396), .A2(n395), .ZN(n424) );
  NOR2_X1 U376 ( .A1(n713), .A2(n591), .ZN(n576) );
  XNOR2_X2 U377 ( .A(n399), .B(G134), .ZN(n522) );
  NAND2_X1 U378 ( .A1(n384), .A2(n380), .ZN(n687) );
  NOR2_X1 U379 ( .A1(n700), .A2(n376), .ZN(n698) );
  NOR2_X1 U380 ( .A1(n725), .A2(n738), .ZN(n726) );
  NOR2_X1 U381 ( .A1(n649), .A2(n738), .ZN(n650) );
  AND2_X1 U382 ( .A1(n632), .A2(n631), .ZN(n758) );
  NOR2_X1 U383 ( .A1(n387), .A2(n620), .ZN(n676) );
  NAND2_X1 U384 ( .A1(n431), .A2(n430), .ZN(n621) );
  AND2_X1 U385 ( .A1(n435), .A2(n434), .ZN(n431) );
  NAND2_X1 U386 ( .A1(n411), .A2(n409), .ZN(n683) );
  AND2_X1 U387 ( .A1(n389), .A2(n429), .ZN(n428) );
  XNOR2_X1 U388 ( .A(n720), .B(n722), .ZN(n723) );
  XNOR2_X1 U389 ( .A(n687), .B(n545), .ZN(n573) );
  XOR2_X1 U390 ( .A(KEYINPUT123), .B(n646), .Z(n647) );
  XNOR2_X1 U391 ( .A(n391), .B(n390), .ZN(n728) );
  AND2_X1 U392 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U393 ( .A(n747), .B(n464), .ZN(n475) );
  XNOR2_X1 U394 ( .A(n463), .B(KEYINPUT87), .ZN(n747) );
  XNOR2_X1 U395 ( .A(n757), .B(G146), .ZN(n505) );
  XNOR2_X1 U396 ( .A(n522), .B(n470), .ZN(n757) );
  XNOR2_X1 U397 ( .A(n438), .B(KEYINPUT4), .ZN(n470) );
  XOR2_X1 U398 ( .A(G131), .B(G140), .Z(n529) );
  XNOR2_X1 U399 ( .A(G146), .B(G125), .ZN(n476) );
  XNOR2_X1 U400 ( .A(KEYINPUT65), .B(KEYINPUT69), .ZN(n438) );
  NAND2_X1 U401 ( .A1(n680), .A2(KEYINPUT81), .ZN(n442) );
  NOR2_X1 U402 ( .A1(n633), .A2(n349), .ZN(n347) );
  NOR2_X1 U403 ( .A1(n347), .A2(n348), .ZN(n443) );
  AND2_X1 U404 ( .A1(n361), .A2(n636), .ZN(n348) );
  OR2_X1 U405 ( .A1(KEYINPUT81), .A2(n350), .ZN(n349) );
  INV_X1 U406 ( .A(n361), .ZN(n350) );
  AND2_X2 U407 ( .A1(n444), .A2(n355), .ZN(n351) );
  AND2_X1 U408 ( .A1(n444), .A2(n355), .ZN(n727) );
  XNOR2_X1 U409 ( .A(n572), .B(n440), .ZN(n620) );
  INV_X1 U410 ( .A(KEYINPUT1), .ZN(n548) );
  NOR2_X1 U411 ( .A1(n405), .A2(n676), .ZN(n404) );
  AND2_X1 U412 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U413 ( .A(n415), .ZN(n414) );
  OR2_X1 U414 ( .A1(n735), .A2(n410), .ZN(n409) );
  NAND2_X1 U415 ( .A1(n415), .A2(n382), .ZN(n410) );
  XNOR2_X1 U416 ( .A(n436), .B(KEYINPUT70), .ZN(n478) );
  INV_X1 U417 ( .A(G137), .ZN(n436) );
  NAND2_X1 U418 ( .A1(n621), .A2(n560), .ZN(n562) );
  INV_X1 U419 ( .A(KEYINPUT85), .ZN(n440) );
  OR2_X1 U420 ( .A1(n641), .A2(n381), .ZN(n380) );
  NAND2_X1 U421 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U422 ( .A(G472), .ZN(n383) );
  INV_X1 U423 ( .A(KEYINPUT71), .ZN(n402) );
  NOR2_X1 U424 ( .A1(n769), .A2(n768), .ZN(n617) );
  NAND2_X1 U425 ( .A1(G902), .A2(G472), .ZN(n385) );
  NAND2_X1 U426 ( .A1(n641), .A2(G472), .ZN(n386) );
  NOR2_X1 U427 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U428 ( .A1(n377), .A2(n375), .ZN(n374) );
  NOR2_X1 U429 ( .A1(n384), .A2(n378), .ZN(n373) );
  NAND2_X1 U430 ( .A1(n376), .A2(n509), .ZN(n375) );
  NAND2_X1 U431 ( .A1(n427), .A2(n382), .ZN(n426) );
  XNOR2_X1 U432 ( .A(G107), .B(G104), .ZN(n462) );
  XNOR2_X1 U433 ( .A(n401), .B(KEYINPUT24), .ZN(n483) );
  INV_X1 U434 ( .A(KEYINPUT94), .ZN(n401) );
  XNOR2_X1 U435 ( .A(n480), .B(n479), .ZN(n519) );
  XNOR2_X1 U436 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U437 ( .A(n478), .ZN(n471) );
  XNOR2_X1 U438 ( .A(n608), .B(n369), .ZN(n712) );
  INV_X1 U439 ( .A(KEYINPUT41), .ZN(n369) );
  INV_X1 U440 ( .A(KEYINPUT40), .ZN(n370) );
  NAND2_X1 U441 ( .A1(n671), .A2(n370), .ZN(n366) );
  INV_X1 U442 ( .A(n554), .ZN(n433) );
  NAND2_X1 U443 ( .A1(n394), .A2(n393), .ZN(n396) );
  NOR2_X1 U444 ( .A1(n573), .A2(n352), .ZN(n393) );
  OR2_X1 U445 ( .A1(n620), .A2(n397), .ZN(n394) );
  AND2_X1 U446 ( .A1(n620), .A2(KEYINPUT102), .ZN(n395) );
  NOR2_X1 U447 ( .A1(n594), .A2(n683), .ZN(n570) );
  INV_X1 U448 ( .A(KEYINPUT22), .ZN(n441) );
  XNOR2_X1 U449 ( .A(n490), .B(n416), .ZN(n415) );
  XNOR2_X1 U450 ( .A(n491), .B(KEYINPUT25), .ZN(n416) );
  NAND2_X1 U451 ( .A1(n547), .A2(n379), .ZN(n378) );
  INV_X1 U452 ( .A(n509), .ZN(n379) );
  OR2_X1 U453 ( .A1(n380), .A2(n378), .ZN(n377) );
  NAND2_X1 U454 ( .A1(n354), .A2(n659), .ZN(n597) );
  XNOR2_X1 U455 ( .A(n466), .B(G902), .ZN(n639) );
  XNOR2_X1 U456 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n466) );
  XOR2_X1 U457 ( .A(KEYINPUT68), .B(G101), .Z(n495) );
  NOR2_X1 U458 ( .A1(n408), .A2(n407), .ZN(n610) );
  INV_X1 U459 ( .A(n411), .ZN(n408) );
  NAND2_X1 U460 ( .A1(n409), .A2(n353), .ZN(n407) );
  NAND2_X1 U461 ( .A1(n398), .A2(n439), .ZN(n397) );
  XNOR2_X1 U462 ( .A(G131), .B(G113), .ZN(n498) );
  XOR2_X1 U463 ( .A(KEYINPUT96), .B(G137), .Z(n499) );
  NOR2_X1 U464 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U465 ( .A(G122), .B(G113), .ZN(n536) );
  XNOR2_X1 U466 ( .A(KEYINPUT3), .B(G119), .ZN(n454) );
  XOR2_X1 U467 ( .A(KEYINPUT9), .B(G122), .Z(n524) );
  XNOR2_X1 U468 ( .A(G116), .B(G107), .ZN(n523) );
  NAND2_X1 U469 ( .A1(n372), .A2(n371), .ZN(n517) );
  NAND2_X1 U470 ( .A1(n356), .A2(n384), .ZN(n371) );
  NAND2_X1 U471 ( .A1(n433), .A2(n358), .ZN(n430) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n589) );
  INV_X1 U473 ( .A(KEYINPUT97), .ZN(n417) );
  NAND2_X1 U474 ( .A1(n420), .A2(n419), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n421), .B(KEYINPUT95), .ZN(n420) );
  INV_X1 U476 ( .A(KEYINPUT64), .ZN(n447) );
  XNOR2_X1 U477 ( .A(n488), .B(n754), .ZN(n735) );
  OR2_X1 U478 ( .A1(n759), .A2(G952), .ZN(n655) );
  XNOR2_X1 U479 ( .A(n475), .B(KEYINPUT79), .ZN(n390) );
  XNOR2_X1 U480 ( .A(n505), .B(n474), .ZN(n391) );
  XNOR2_X1 U481 ( .A(n473), .B(n755), .ZN(n474) );
  XNOR2_X1 U482 ( .A(n368), .B(KEYINPUT42), .ZN(n768) );
  NOR2_X1 U483 ( .A1(n712), .A2(n615), .ZN(n368) );
  NAND2_X1 U484 ( .A1(n365), .A2(n363), .ZN(n769) );
  AND2_X1 U485 ( .A1(n367), .A2(n366), .ZN(n365) );
  XNOR2_X1 U486 ( .A(n619), .B(KEYINPUT36), .ZN(n387) );
  NAND2_X1 U487 ( .A1(n568), .A2(n424), .ZN(n423) );
  INV_X1 U488 ( .A(KEYINPUT103), .ZN(n400) );
  AND2_X1 U489 ( .A1(n683), .A2(KEYINPUT102), .ZN(n352) );
  AND2_X1 U490 ( .A1(n682), .A2(n544), .ZN(n353) );
  OR2_X1 U491 ( .A1(n673), .A2(n623), .ZN(n354) );
  NAND2_X2 U492 ( .A1(n428), .A2(n425), .ZN(n609) );
  AND2_X1 U493 ( .A1(n380), .A2(n509), .ZN(n356) );
  AND2_X1 U494 ( .A1(n433), .A2(n547), .ZN(n357) );
  INV_X1 U495 ( .A(n683), .ZN(n398) );
  INV_X1 U496 ( .A(n687), .ZN(n419) );
  AND2_X1 U497 ( .A1(n547), .A2(n432), .ZN(n358) );
  AND2_X1 U498 ( .A1(n419), .A2(n570), .ZN(n359) );
  AND2_X1 U499 ( .A1(n596), .A2(n595), .ZN(n360) );
  INV_X1 U500 ( .A(G902), .ZN(n382) );
  INV_X1 U501 ( .A(n547), .ZN(n376) );
  INV_X1 U502 ( .A(KEYINPUT102), .ZN(n439) );
  NAND2_X1 U503 ( .A1(n639), .A2(n638), .ZN(n361) );
  XNOR2_X1 U504 ( .A(n362), .B(n583), .ZN(n600) );
  NAND2_X1 U505 ( .A1(n581), .A2(n582), .ZN(n362) );
  NAND2_X1 U506 ( .A1(n629), .A2(n370), .ZN(n367) );
  XNOR2_X1 U507 ( .A(n607), .B(KEYINPUT39), .ZN(n629) );
  OR2_X1 U508 ( .A1(n629), .A2(n364), .ZN(n363) );
  OR2_X1 U509 ( .A1(n671), .A2(n370), .ZN(n364) );
  NAND2_X1 U510 ( .A1(n610), .A2(n573), .ZN(n546) );
  NAND2_X1 U511 ( .A1(n392), .A2(n388), .ZN(n437) );
  XNOR2_X1 U512 ( .A(n388), .B(G110), .ZN(G12) );
  XNOR2_X2 U513 ( .A(n422), .B(n400), .ZN(n388) );
  NAND2_X1 U514 ( .A1(n728), .A2(n445), .ZN(n389) );
  XNOR2_X2 U515 ( .A(G143), .B(G128), .ZN(n399) );
  XNOR2_X1 U516 ( .A(n392), .B(G119), .ZN(G21) );
  XNOR2_X2 U517 ( .A(n423), .B(n569), .ZN(n392) );
  XNOR2_X1 U518 ( .A(n399), .B(n476), .ZN(n446) );
  NAND2_X1 U519 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X1 U520 ( .A1(n739), .A2(n758), .ZN(n633) );
  XNOR2_X1 U521 ( .A(n603), .B(n602), .ZN(n739) );
  XNOR2_X1 U522 ( .A(n403), .B(n402), .ZN(n626) );
  NAND2_X1 U523 ( .A1(n406), .A2(n404), .ZN(n403) );
  INV_X1 U524 ( .A(n625), .ZN(n405) );
  XNOR2_X1 U525 ( .A(n624), .B(KEYINPUT47), .ZN(n406) );
  NAND2_X1 U526 ( .A1(n414), .A2(G902), .ZN(n412) );
  NAND2_X1 U527 ( .A1(n735), .A2(n414), .ZN(n413) );
  NAND2_X1 U528 ( .A1(n587), .A2(n588), .ZN(n421) );
  NAND2_X1 U529 ( .A1(n568), .A2(n359), .ZN(n422) );
  XNOR2_X2 U530 ( .A(n609), .B(n548), .ZN(n572) );
  OR2_X1 U531 ( .A1(n728), .A2(n426), .ZN(n425) );
  INV_X1 U532 ( .A(n445), .ZN(n427) );
  NAND2_X1 U533 ( .A1(n445), .A2(G902), .ZN(n429) );
  XNOR2_X2 U534 ( .A(n567), .B(n441), .ZN(n568) );
  INV_X1 U535 ( .A(n555), .ZN(n432) );
  NAND2_X1 U536 ( .A1(n376), .A2(n555), .ZN(n434) );
  NAND2_X1 U537 ( .A1(n554), .A2(n555), .ZN(n435) );
  XNOR2_X1 U538 ( .A(n437), .B(n571), .ZN(n582) );
  NAND2_X1 U539 ( .A1(n568), .A2(n360), .ZN(n659) );
  BUF_X1 U540 ( .A(n554), .Z(n605) );
  XNOR2_X1 U541 ( .A(KEYINPUT72), .B(G469), .ZN(n445) );
  INV_X1 U542 ( .A(KEYINPUT84), .ZN(n571) );
  INV_X1 U543 ( .A(KEYINPUT46), .ZN(n616) );
  XNOR2_X1 U544 ( .A(n617), .B(n616), .ZN(n627) );
  INV_X1 U545 ( .A(KEYINPUT8), .ZN(n479) );
  NOR2_X1 U546 ( .A1(n494), .A2(n689), .ZN(n588) );
  XNOR2_X1 U547 ( .A(n446), .B(n470), .ZN(n453) );
  XNOR2_X2 U548 ( .A(n447), .B(G953), .ZN(n759) );
  NAND2_X1 U549 ( .A1(n759), .A2(G224), .ZN(n451) );
  XNOR2_X1 U550 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n449) );
  XNOR2_X1 U551 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n448) );
  XNOR2_X1 U552 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U553 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U554 ( .A(n453), .B(n452), .ZN(n456) );
  XNOR2_X1 U555 ( .A(n454), .B(G116), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n536), .B(KEYINPUT16), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n496), .B(n455), .ZN(n749) );
  XNOR2_X1 U558 ( .A(n456), .B(n749), .ZN(n465) );
  INV_X1 U559 ( .A(G110), .ZN(n457) );
  NAND2_X1 U560 ( .A1(n457), .A2(KEYINPUT75), .ZN(n460) );
  INV_X1 U561 ( .A(KEYINPUT75), .ZN(n458) );
  NAND2_X1 U562 ( .A1(n458), .A2(G110), .ZN(n459) );
  NAND2_X1 U563 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U564 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U565 ( .A(n495), .B(KEYINPUT73), .ZN(n464) );
  XNOR2_X1 U566 ( .A(n465), .B(n475), .ZN(n720) );
  NAND2_X1 U567 ( .A1(n720), .A2(n639), .ZN(n469) );
  INV_X1 U568 ( .A(G237), .ZN(n467) );
  NAND2_X1 U569 ( .A1(n382), .A2(n467), .ZN(n506) );
  NAND2_X1 U570 ( .A1(n506), .A2(G210), .ZN(n468) );
  NAND2_X1 U571 ( .A1(n759), .A2(G227), .ZN(n472) );
  XOR2_X1 U572 ( .A(KEYINPUT93), .B(n529), .Z(n755) );
  INV_X1 U573 ( .A(n609), .ZN(n494) );
  XOR2_X1 U574 ( .A(KEYINPUT10), .B(n476), .Z(n530) );
  INV_X1 U575 ( .A(n530), .ZN(n477) );
  XOR2_X1 U576 ( .A(n478), .B(n477), .Z(n754) );
  NAND2_X1 U577 ( .A1(n759), .A2(G234), .ZN(n480) );
  NAND2_X1 U578 ( .A1(n519), .A2(G221), .ZN(n487) );
  XNOR2_X1 U579 ( .A(G119), .B(G110), .ZN(n481) );
  XNOR2_X1 U580 ( .A(n481), .B(KEYINPUT23), .ZN(n485) );
  XNOR2_X1 U581 ( .A(G128), .B(G140), .ZN(n482) );
  XNOR2_X1 U582 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U583 ( .A(n485), .B(n484), .Z(n486) );
  XNOR2_X1 U584 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U585 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n491) );
  NAND2_X1 U586 ( .A1(G234), .A2(n639), .ZN(n489) );
  XNOR2_X1 U587 ( .A(n489), .B(KEYINPUT20), .ZN(n492) );
  NAND2_X1 U588 ( .A1(n492), .A2(G217), .ZN(n490) );
  NAND2_X1 U589 ( .A1(G221), .A2(n492), .ZN(n493) );
  XOR2_X1 U590 ( .A(KEYINPUT21), .B(n493), .Z(n682) );
  NAND2_X1 U591 ( .A1(n683), .A2(n682), .ZN(n689) );
  XNOR2_X1 U592 ( .A(n495), .B(KEYINPUT5), .ZN(n497) );
  XNOR2_X1 U593 ( .A(n497), .B(n496), .ZN(n503) );
  XNOR2_X1 U594 ( .A(n499), .B(n498), .ZN(n501) );
  NOR2_X1 U595 ( .A1(G953), .A2(G237), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n533), .A2(G210), .ZN(n500) );
  XNOR2_X1 U597 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U598 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U599 ( .A(n505), .B(n504), .ZN(n641) );
  NAND2_X1 U600 ( .A1(n506), .A2(G214), .ZN(n508) );
  INV_X1 U601 ( .A(KEYINPUT89), .ZN(n507) );
  XNOR2_X1 U602 ( .A(n508), .B(n507), .ZN(n547) );
  XNOR2_X1 U603 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n509) );
  NAND2_X1 U604 ( .A1(G234), .A2(G237), .ZN(n510) );
  XNOR2_X1 U605 ( .A(n510), .B(KEYINPUT14), .ZN(n513) );
  NAND2_X1 U606 ( .A1(G952), .A2(n513), .ZN(n711) );
  NOR2_X1 U607 ( .A1(G953), .A2(n711), .ZN(n512) );
  INV_X1 U608 ( .A(KEYINPUT90), .ZN(n511) );
  XNOR2_X1 U609 ( .A(n512), .B(n511), .ZN(n559) );
  NAND2_X1 U610 ( .A1(n513), .A2(G902), .ZN(n514) );
  XNOR2_X1 U611 ( .A(n514), .B(KEYINPUT91), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n759), .A2(G900), .ZN(n515) );
  NAND2_X1 U613 ( .A1(n556), .A2(n515), .ZN(n516) );
  NAND2_X1 U614 ( .A1(n559), .A2(n516), .ZN(n544) );
  AND2_X1 U615 ( .A1(n517), .A2(n544), .ZN(n518) );
  NAND2_X1 U616 ( .A1(n588), .A2(n518), .ZN(n606) );
  XOR2_X1 U617 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n521) );
  NAND2_X1 U618 ( .A1(G217), .A2(n519), .ZN(n520) );
  XNOR2_X1 U619 ( .A(n521), .B(n520), .ZN(n527) );
  XNOR2_X1 U620 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U621 ( .A(n522), .B(n525), .Z(n526) );
  XNOR2_X1 U622 ( .A(n527), .B(n526), .ZN(n646) );
  NOR2_X1 U623 ( .A1(n646), .A2(G902), .ZN(n528) );
  XOR2_X1 U624 ( .A(n528), .B(G478), .Z(n563) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(G475), .ZN(n542) );
  XNOR2_X1 U626 ( .A(n530), .B(n529), .ZN(n532) );
  XNOR2_X1 U627 ( .A(G143), .B(G104), .ZN(n531) );
  XNOR2_X1 U628 ( .A(n532), .B(n531), .ZN(n540) );
  XOR2_X1 U629 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n535) );
  NAND2_X1 U630 ( .A1(G214), .A2(n533), .ZN(n534) );
  XNOR2_X1 U631 ( .A(n535), .B(n534), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n536), .B(KEYINPUT98), .ZN(n537) );
  XNOR2_X1 U633 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U634 ( .A(n540), .B(n539), .ZN(n652) );
  NOR2_X1 U635 ( .A1(G902), .A2(n652), .ZN(n541) );
  XNOR2_X1 U636 ( .A(n542), .B(n541), .ZN(n585) );
  NAND2_X1 U637 ( .A1(n563), .A2(n585), .ZN(n577) );
  NOR2_X1 U638 ( .A1(n606), .A2(n577), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n433), .A2(n543), .ZN(n625) );
  XNOR2_X1 U640 ( .A(n625), .B(G143), .ZN(G45) );
  INV_X1 U641 ( .A(n563), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n585), .A2(n584), .ZN(n671) );
  INV_X1 U643 ( .A(KEYINPUT6), .ZN(n545) );
  NOR2_X1 U644 ( .A1(n671), .A2(n546), .ZN(n618) );
  INV_X1 U645 ( .A(n572), .ZN(n594) );
  NOR2_X1 U646 ( .A1(n376), .A2(n594), .ZN(n549) );
  NAND2_X1 U647 ( .A1(n618), .A2(n549), .ZN(n550) );
  XNOR2_X1 U648 ( .A(KEYINPUT106), .B(n550), .ZN(n552) );
  XNOR2_X1 U649 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n551) );
  XOR2_X1 U650 ( .A(n552), .B(n551), .Z(n553) );
  NAND2_X1 U651 ( .A1(n553), .A2(n605), .ZN(n630) );
  XNOR2_X1 U652 ( .A(n630), .B(G140), .ZN(G42) );
  INV_X1 U653 ( .A(n573), .ZN(n595) );
  XNOR2_X1 U654 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n555) );
  INV_X1 U655 ( .A(G953), .ZN(n740) );
  NOR2_X1 U656 ( .A1(G898), .A2(n740), .ZN(n751) );
  NAND2_X1 U657 ( .A1(n556), .A2(n751), .ZN(n557) );
  XNOR2_X1 U658 ( .A(n557), .B(KEYINPUT92), .ZN(n558) );
  NAND2_X1 U659 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U660 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n561) );
  XNOR2_X2 U661 ( .A(n562), .B(n561), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n563), .A2(n585), .ZN(n701) );
  AND2_X1 U663 ( .A1(n701), .A2(n682), .ZN(n565) );
  INV_X1 U664 ( .A(KEYINPUT101), .ZN(n564) );
  XNOR2_X1 U665 ( .A(n565), .B(n564), .ZN(n566) );
  NAND2_X1 U666 ( .A1(n587), .A2(n566), .ZN(n567) );
  XNOR2_X1 U667 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n569) );
  NAND2_X1 U668 ( .A1(n573), .A2(n590), .ZN(n575) );
  XOR2_X1 U669 ( .A(KEYINPUT104), .B(KEYINPUT33), .Z(n574) );
  INV_X1 U670 ( .A(n587), .ZN(n591) );
  XNOR2_X1 U671 ( .A(n576), .B(KEYINPUT34), .ZN(n579) );
  INV_X1 U672 ( .A(n577), .ZN(n578) );
  NAND2_X1 U673 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U674 ( .A(n767), .ZN(n581) );
  INV_X1 U675 ( .A(KEYINPUT44), .ZN(n583) );
  NOR2_X1 U676 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U677 ( .A(KEYINPUT100), .B(n586), .Z(n674) );
  NOR2_X1 U678 ( .A1(n674), .A2(n589), .ZN(n662) );
  NOR2_X1 U679 ( .A1(n671), .A2(n589), .ZN(n661) );
  OR2_X1 U680 ( .A1(n662), .A2(n661), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n590), .A2(n687), .ZN(n693) );
  OR2_X1 U682 ( .A1(n693), .A2(n591), .ZN(n593) );
  INV_X1 U683 ( .A(KEYINPUT31), .ZN(n592) );
  XNOR2_X1 U684 ( .A(n593), .B(n592), .ZN(n673) );
  NAND2_X1 U685 ( .A1(n671), .A2(n674), .ZN(n699) );
  INV_X1 U686 ( .A(n699), .ZN(n623) );
  NOR2_X1 U687 ( .A1(n594), .A2(n398), .ZN(n596) );
  NOR2_X1 U688 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U689 ( .A1(n600), .A2(n599), .ZN(n603) );
  INV_X1 U690 ( .A(KEYINPUT83), .ZN(n601) );
  XNOR2_X1 U691 ( .A(n601), .B(KEYINPUT45), .ZN(n602) );
  XOR2_X1 U692 ( .A(KEYINPUT74), .B(KEYINPUT38), .Z(n604) );
  XNOR2_X1 U693 ( .A(n605), .B(n604), .ZN(n700) );
  NOR2_X1 U694 ( .A1(n606), .A2(n700), .ZN(n607) );
  NAND2_X1 U695 ( .A1(n701), .A2(n698), .ZN(n608) );
  XOR2_X1 U696 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n612) );
  NAND2_X1 U697 ( .A1(n687), .A2(n610), .ZN(n611) );
  XNOR2_X1 U698 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n609), .A2(n613), .ZN(n614) );
  XNOR2_X1 U700 ( .A(KEYINPUT109), .B(n614), .ZN(n622) );
  INV_X1 U701 ( .A(n622), .ZN(n615) );
  NAND2_X1 U702 ( .A1(n618), .A2(n357), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n669) );
  NOR2_X1 U704 ( .A1(n669), .A2(n623), .ZN(n624) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT48), .ZN(n632) );
  OR2_X1 U706 ( .A1(n629), .A2(n674), .ZN(n679) );
  AND2_X1 U707 ( .A1(n630), .A2(n679), .ZN(n631) );
  BUF_X2 U708 ( .A(n633), .Z(n680) );
  INV_X1 U709 ( .A(n639), .ZN(n635) );
  NAND2_X1 U710 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n640) );
  NOR2_X1 U713 ( .A1(KEYINPUT82), .A2(n640), .ZN(n637) );
  NOR2_X1 U714 ( .A1(KEYINPUT81), .A2(n637), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n351), .A2(G472), .ZN(n643) );
  XOR2_X1 U716 ( .A(KEYINPUT62), .B(n641), .Z(n642) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n644), .A2(n655), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U720 ( .A1(n727), .A2(G478), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(n649) );
  INV_X1 U722 ( .A(n655), .ZN(n738) );
  XNOR2_X1 U723 ( .A(n650), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U724 ( .A1(n351), .A2(G475), .ZN(n654) );
  XOR2_X1 U725 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n658) );
  XOR2_X1 U729 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n657) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(G60) );
  INV_X1 U731 ( .A(n659), .ZN(n660) );
  XOR2_X1 U732 ( .A(G101), .B(n660), .Z(G3) );
  XOR2_X1 U733 ( .A(G104), .B(n661), .Z(G6) );
  XNOR2_X1 U734 ( .A(n662), .B(KEYINPUT27), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(KEYINPUT26), .ZN(n664) );
  XNOR2_X1 U736 ( .A(G107), .B(n664), .ZN(G9) );
  NOR2_X1 U737 ( .A1(n669), .A2(n674), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n666) );
  XNOR2_X1 U739 ( .A(G128), .B(KEYINPUT111), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(G30) );
  NOR2_X1 U742 ( .A1(n669), .A2(n671), .ZN(n670) );
  XOR2_X1 U743 ( .A(G146), .B(n670), .Z(G48) );
  NOR2_X1 U744 ( .A1(n671), .A2(n673), .ZN(n672) );
  XOR2_X1 U745 ( .A(G113), .B(n672), .Z(G15) );
  NOR2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U747 ( .A(G116), .B(n675), .Z(G18) );
  XNOR2_X1 U748 ( .A(n676), .B(KEYINPUT112), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT37), .ZN(n678) );
  XNOR2_X1 U750 ( .A(G125), .B(n678), .ZN(G27) );
  XNOR2_X1 U751 ( .A(G134), .B(n679), .ZN(G36) );
  XOR2_X1 U752 ( .A(KEYINPUT2), .B(n680), .Z(n717) );
  XNOR2_X1 U753 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n681), .B(KEYINPUT51), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n685) );
  XNOR2_X1 U756 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n684) );
  XNOR2_X1 U757 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U758 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT114), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n572), .A2(n689), .ZN(n690) );
  XNOR2_X1 U761 ( .A(KEYINPUT50), .B(n690), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U764 ( .A(n696), .B(n695), .Z(n697) );
  NOR2_X1 U765 ( .A1(n712), .A2(n697), .ZN(n707) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U767 ( .A1(n700), .A2(n376), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U770 ( .A1(n713), .A2(n705), .ZN(n706) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U772 ( .A(n708), .B(KEYINPUT117), .Z(n709) );
  XNOR2_X1 U773 ( .A(KEYINPUT52), .B(n709), .ZN(n710) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U777 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U778 ( .A1(n718), .A2(G953), .ZN(n719) );
  XNOR2_X1 U779 ( .A(n719), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U780 ( .A1(n727), .A2(G210), .ZN(n724) );
  XOR2_X1 U781 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n721) );
  XOR2_X1 U782 ( .A(n721), .B(KEYINPUT55), .Z(n722) );
  XNOR2_X1 U783 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U784 ( .A(n726), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U785 ( .A1(n351), .A2(G469), .ZN(n733) );
  XOR2_X1 U786 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n730) );
  XNOR2_X1 U787 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n730), .B(n729), .ZN(n731) );
  XOR2_X1 U789 ( .A(n728), .B(n731), .Z(n732) );
  XNOR2_X1 U790 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U791 ( .A1(n738), .A2(n734), .ZN(G54) );
  NAND2_X1 U792 ( .A1(n351), .A2(G217), .ZN(n736) );
  XNOR2_X1 U793 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U794 ( .A1(n738), .A2(n737), .ZN(G66) );
  BUF_X1 U795 ( .A(n739), .Z(n741) );
  NAND2_X1 U796 ( .A1(n741), .A2(n740), .ZN(n746) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n742) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n742), .ZN(n743) );
  NAND2_X1 U799 ( .A1(n743), .A2(G898), .ZN(n744) );
  XOR2_X1 U800 ( .A(KEYINPUT125), .B(n744), .Z(n745) );
  NAND2_X1 U801 ( .A1(n746), .A2(n745), .ZN(n753) );
  XNOR2_X1 U802 ( .A(n747), .B(G101), .ZN(n748) );
  XOR2_X1 U803 ( .A(n749), .B(n748), .Z(n750) );
  NOR2_X1 U804 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U805 ( .A(n753), .B(n752), .ZN(G69) );
  XOR2_X1 U806 ( .A(n755), .B(n754), .Z(n756) );
  XOR2_X1 U807 ( .A(n757), .B(n756), .Z(n761) );
  XOR2_X1 U808 ( .A(n761), .B(n758), .Z(n760) );
  NAND2_X1 U809 ( .A1(n760), .A2(n759), .ZN(n765) );
  XNOR2_X1 U810 ( .A(G227), .B(n761), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n762), .A2(G900), .ZN(n763) );
  NAND2_X1 U812 ( .A1(G953), .A2(n763), .ZN(n764) );
  NAND2_X1 U813 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U814 ( .A(KEYINPUT126), .B(n766), .ZN(G72) );
  XOR2_X1 U815 ( .A(n767), .B(G122), .Z(G24) );
  XOR2_X1 U816 ( .A(G137), .B(n768), .Z(G39) );
  XOR2_X1 U817 ( .A(G131), .B(n769), .Z(G33) );
endmodule

