//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G137), .A4(new_n463), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n467), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n464), .A2(new_n463), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n469), .A2(new_n471), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n483), .A2(KEYINPUT66), .A3(new_n463), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT66), .B1(new_n483), .B2(new_n463), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n479), .B(new_n482), .C1(new_n487), .C2(G124), .ZN(G162));
  NAND4_X1  g063(.A1(new_n469), .A2(new_n471), .A3(G126), .A4(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n463), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n464), .A2(new_n496), .A3(G138), .A4(new_n463), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  AND2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G50), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n499), .A2(new_n500), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  OAI221_X1 g087(.A(new_n504), .B1(new_n509), .B2(new_n510), .C1(new_n511), .C2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n505), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n506), .A2(new_n507), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n505), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT68), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n526), .B1(new_n519), .B2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(G168));
  NOR2_X1   g103(.A1(new_n520), .A2(new_n501), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G90), .B1(G52), .B2(new_n503), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n511), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT69), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n517), .B1(new_n509), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n511), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n529), .A2(G91), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n506), .B2(new_n507), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n499), .C2(new_n500), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(KEYINPUT70), .B1(new_n559), .B2(KEYINPUT71), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND2_X1  g145(.A1(new_n529), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n503), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  INV_X1    g149(.A(G48), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n575), .A2(new_n517), .B1(new_n509), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT74), .Z(new_n579));
  NAND3_X1  g154(.A1(new_n508), .A2(KEYINPUT73), .A3(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT73), .B1(new_n508), .B2(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n577), .B1(new_n583), .B2(KEYINPUT75), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(G651), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G305));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n517), .B1(new_n509), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n511), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n594), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n592), .A2(new_n511), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT76), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n595), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n603), .A2(KEYINPUT77), .A3(new_n591), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G290));
  NAND3_X1  g180(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n509), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n520), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(G651), .B1(new_n503), .B2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g192(.A(new_n616), .B1(G171), .B2(G868), .ZN(G321));
  MUX2_X1   g193(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g194(.A(G280), .B(KEYINPUT78), .ZN(G297));
  AND2_X1   g195(.A1(new_n610), .A2(new_n614), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  OAI21_X1  g198(.A(KEYINPUT79), .B1(new_n543), .B2(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n622), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  MUX2_X1   g201(.A(KEYINPUT79), .B(new_n624), .S(new_n626), .Z(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n487), .A2(G123), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n463), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n478), .A2(G135), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n478), .A2(G2104), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n636), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n477), .B2(new_n468), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2100), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n642), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT15), .B(G2435), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT81), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n648), .A2(new_n649), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n649), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT82), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT16), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n657), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n660), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n647), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n658), .A2(new_n660), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(new_n646), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT83), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n674));
  NAND4_X1  g249(.A1(new_n666), .A2(new_n674), .A3(new_n671), .A4(new_n668), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n645), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AND3_X1   g251(.A1(new_n669), .A2(new_n670), .A3(new_n646), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n646), .B1(new_n669), .B2(new_n670), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n667), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g256(.A(KEYINPUT84), .B(new_n667), .C1(new_n677), .C2(new_n678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n676), .A2(new_n683), .ZN(G401));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  XNOR2_X1  g260(.A(G2067), .B(G2678), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(KEYINPUT17), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  AOI21_X1  g264(.A(KEYINPUT18), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2072), .B(G2078), .Z(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n687), .B2(KEYINPUT18), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2096), .B(G2100), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1956), .B(G2474), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT19), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n699), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n702), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n703), .A2(KEYINPUT20), .A3(new_n702), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n704), .B1(new_n702), .B2(new_n700), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT87), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n709), .B(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT86), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1991), .B(G1996), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT88), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n713), .A2(new_n718), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(G229));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G23), .ZN(new_n723));
  INV_X1    g298(.A(G288), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n722), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT33), .B(G1976), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT95), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n722), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n722), .ZN(new_n730));
  INV_X1    g305(.A(G1971), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n728), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n722), .A2(G6), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G305), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT32), .B(G1981), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT94), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n734), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n736), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(KEYINPUT34), .ZN(new_n743));
  INV_X1    g318(.A(G290), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(new_n722), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n722), .B2(G24), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT93), .B(G1986), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G25), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT89), .Z(new_n751));
  NAND3_X1  g326(.A1(new_n464), .A2(G131), .A3(new_n463), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n484), .A2(G119), .A3(new_n485), .ZN(new_n755));
  OR2_X1    g330(.A1(G95), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT35), .B(G1991), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT91), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT92), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n759), .B(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n746), .B2(new_n747), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n742), .A2(new_n743), .A3(new_n748), .A4(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n722), .A2(G19), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n543), .B2(new_n722), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1341), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT31), .B(G11), .Z(new_n771));
  NOR2_X1   g346(.A1(new_n634), .A2(new_n749), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n749), .B1(new_n773), .B2(G28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(KEYINPUT101), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(KEYINPUT101), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n773), .B2(G28), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n771), .B(new_n772), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  NOR2_X1   g354(.A1(G27), .A2(G29), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G164), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  INV_X1    g358(.A(G34), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT24), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(KEYINPUT24), .ZN(new_n786));
  AOI22_X1  g361(.A1(G160), .A2(G29), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n778), .B1(new_n779), .B2(new_n782), .C1(new_n783), .C2(new_n788), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n770), .B(new_n789), .C1(new_n779), .C2(new_n782), .ZN(new_n790));
  NOR2_X1   g365(.A1(G4), .A2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT97), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n615), .B2(new_n722), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT98), .B(G1348), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n793), .B(new_n794), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n749), .A2(G33), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT25), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n464), .A2(G127), .ZN(new_n799));
  NAND2_X1  g374(.A1(G115), .A2(G2104), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n463), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n798), .B(new_n801), .C1(G139), .C2(new_n478), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n749), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(G2072), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n803), .A2(G2072), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n804), .B(new_n805), .C1(new_n783), .C2(new_n788), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n790), .A2(new_n795), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n749), .A2(G35), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT102), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n749), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT29), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n811), .A2(G2090), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT103), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n749), .A2(G26), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT28), .ZN(new_n815));
  INV_X1    g390(.A(G128), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT99), .B1(new_n486), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n484), .A2(new_n818), .A3(new_n485), .A4(G128), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n463), .A2(G116), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n478), .A2(G140), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n815), .B1(new_n826), .B2(new_n749), .ZN(new_n827));
  INV_X1    g402(.A(G2067), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n749), .A2(G32), .ZN(new_n830));
  NAND3_X1  g405(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT26), .Z(new_n832));
  NAND3_X1  g407(.A1(new_n464), .A2(G141), .A3(new_n463), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n473), .A2(G105), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n484), .A2(G129), .A3(new_n485), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT100), .ZN(new_n837));
  AOI21_X1  g412(.A(KEYINPUT100), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n830), .B1(new_n839), .B2(new_n749), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT27), .B(G1996), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n722), .A2(G20), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT23), .Z(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G299), .B2(G16), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1956), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n813), .A2(new_n829), .A3(new_n842), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(G5), .A2(G16), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G171), .B2(G16), .ZN(new_n849));
  INV_X1    g424(.A(G1961), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(G16), .A2(G21), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G168), .B2(G16), .ZN(new_n853));
  INV_X1    g428(.A(G1966), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n851), .B(new_n855), .C1(new_n811), .C2(G2090), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n812), .A2(KEYINPUT103), .ZN(new_n857));
  NOR4_X1   g432(.A1(new_n807), .A2(new_n847), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n767), .A2(new_n858), .ZN(G311));
  NAND2_X1  g434(.A1(new_n767), .A2(new_n858), .ZN(G150));
  NAND2_X1  g435(.A1(new_n621), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  INV_X1    g437(.A(G55), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n863), .A2(new_n517), .B1(new_n509), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(new_n511), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n543), .A2(new_n868), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n542), .A2(new_n540), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n862), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n873));
  AOI21_X1  g448(.A(G860), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n873), .B2(new_n872), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT104), .ZN(new_n876));
  OAI21_X1  g451(.A(G860), .B1(new_n865), .B2(new_n867), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(G145));
  NAND2_X1  g454(.A1(new_n835), .A2(new_n836), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n802), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n802), .B1(new_n837), .B2(new_n838), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n495), .A2(new_n497), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n489), .A2(new_n492), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n820), .B2(new_n824), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n820), .A2(new_n886), .A3(new_n824), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n820), .A2(new_n886), .A3(new_n824), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n882), .B(new_n881), .C1(new_n891), .C2(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n478), .A2(G142), .ZN(new_n893));
  OR2_X1    g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n894), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  INV_X1    g472(.A(G130), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n486), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n484), .A2(KEYINPUT105), .A3(new_n485), .A4(G130), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n640), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n758), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n640), .A2(new_n754), .A3(new_n755), .A4(new_n757), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n899), .A2(new_n900), .ZN(new_n906));
  INV_X1    g481(.A(new_n896), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n903), .A2(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n890), .A2(new_n892), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n634), .B(G160), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(G162), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n890), .A2(new_n892), .ZN(new_n915));
  INV_X1    g490(.A(new_n909), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(KEYINPUT106), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n890), .A2(new_n892), .A3(new_n909), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n921), .A3(new_n917), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n922), .A2(KEYINPUT107), .A3(new_n913), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT107), .B1(new_n922), .B2(new_n913), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT77), .B1(new_n603), .B2(new_n591), .ZN(new_n928));
  AOI211_X1 g503(.A(new_n599), .B(new_n590), .C1(new_n602), .C2(new_n595), .ZN(new_n929));
  OAI21_X1  g504(.A(G288), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n600), .A2(new_n604), .A3(new_n724), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT108), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G305), .B(G303), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n933), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n937), .B2(new_n932), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n927), .B1(new_n939), .B2(KEYINPUT110), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n938), .B2(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n871), .B(new_n625), .Z(new_n944));
  NAND3_X1  g519(.A1(new_n563), .A2(new_n567), .A3(new_n621), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n557), .A2(new_n562), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n615), .B1(new_n946), .B2(new_n566), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n945), .A2(KEYINPUT41), .A3(new_n947), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT41), .B1(new_n945), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n944), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n927), .B(new_n941), .C1(new_n939), .C2(KEYINPUT110), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n943), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n943), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G868), .B2(new_n868), .ZN(G295));
  OAI21_X1  g533(.A(new_n957), .B1(G868), .B2(new_n868), .ZN(G331));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  NAND3_X1  g536(.A1(G171), .A2(new_n525), .A3(new_n527), .ZN(new_n962));
  NAND3_X1  g537(.A1(G168), .A2(new_n536), .A3(new_n535), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n871), .ZN(new_n965));
  INV_X1    g540(.A(new_n871), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n965), .B(new_n967), .C1(new_n951), .C2(new_n950), .ZN(new_n968));
  INV_X1    g543(.A(new_n967), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n962), .B2(new_n963), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n948), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n961), .B1(new_n972), .B2(new_n938), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n971), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n939), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n960), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n939), .B2(new_n974), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n938), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(KEYINPUT43), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n973), .A2(new_n975), .ZN(new_n982));
  NAND2_X1  g557(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n982), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(new_n984), .B2(new_n980), .ZN(G397));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n467), .A2(new_n989), .A3(new_n475), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n839), .A2(new_n986), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(KEYINPUT113), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n994), .A2(KEYINPUT113), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n825), .B(new_n828), .ZN(new_n997));
  INV_X1    g572(.A(new_n880), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n986), .B2(new_n998), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n995), .B(new_n996), .C1(new_n999), .C2(new_n992), .ZN(new_n1000));
  INV_X1    g575(.A(new_n992), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n758), .B(new_n761), .Z(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1986), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n744), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n744), .A2(new_n1004), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1001), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1003), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1012), .B(new_n1015), .C1(G166), .C2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(G303), .A2(new_n1013), .A3(new_n1014), .A4(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n886), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n988), .A2(new_n1022), .A3(new_n990), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n731), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n884), .B2(new_n885), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n990), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT116), .A3(new_n990), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1024), .B1(new_n1033), .B2(G2090), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1020), .B1(new_n1034), .B2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(G2090), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1030), .A2(new_n1031), .A3(new_n1036), .A4(new_n990), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1016), .B1(new_n1024), .B2(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1038), .A2(new_n1020), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1023), .B2(G2078), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1030), .A2(new_n1031), .A3(new_n990), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n850), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1022), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n990), .B1(new_n1025), .B2(KEYINPUT45), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(KEYINPUT118), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n988), .A2(new_n1049), .A3(new_n990), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G301), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n584), .A2(new_n1054), .A3(new_n586), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(new_n584), .B2(new_n586), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G305), .A2(G1981), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n584), .A2(new_n1054), .A3(new_n586), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n990), .A2(new_n1025), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1016), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n724), .A2(G1976), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT52), .B1(G288), .B2(new_n1067), .ZN(new_n1068));
  AND4_X1   g643(.A1(G8), .A2(new_n1066), .A3(new_n1068), .A4(new_n1061), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(KEYINPUT52), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1064), .A2(new_n1065), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1065), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1040), .B(new_n1052), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1043), .A2(G2084), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1047), .A2(KEYINPUT118), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1050), .A3(new_n1022), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1078), .B2(new_n854), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G286), .A2(G8), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1079), .B2(new_n1016), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1966), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT124), .B(G8), .C1(new_n1084), .C2(new_n1076), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n1084), .B2(new_n1076), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1080), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1087), .A2(new_n1088), .B1(KEYINPUT51), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1083), .A2(new_n1085), .A3(KEYINPUT125), .A4(new_n1086), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1081), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1075), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT62), .B(new_n1081), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1089), .A2(G286), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1040), .B(new_n1098), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1039), .A2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1038), .A2(new_n1020), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1102), .A2(new_n1104), .A3(new_n1098), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1039), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G288), .A2(G1976), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1055), .B1(new_n1064), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1063), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT115), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1107), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1101), .A2(new_n1106), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1023), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(KEYINPUT53), .A3(new_n779), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1044), .A3(new_n1042), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1116), .B1(new_n1052), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT126), .B(new_n1116), .C1(new_n1052), .C2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1045), .A2(G301), .A3(new_n1051), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1119), .A2(G171), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(KEYINPUT54), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1040), .B(new_n1128), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1956), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1033), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT57), .B1(new_n946), .B2(new_n566), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n567), .A2(new_n557), .A3(new_n1134), .A4(new_n562), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(G2072), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n988), .A2(new_n1022), .A3(new_n990), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1132), .A2(new_n1137), .A3(new_n1141), .ZN(new_n1142));
  NOR3_X1   g717(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1144));
  AOI21_X1  g719(.A(G1956), .B1(new_n1144), .B2(new_n1032), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1136), .B1(new_n1145), .B2(new_n1140), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(new_n1146), .A3(KEYINPUT61), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1043), .A2(new_n794), .B1(new_n1062), .B2(new_n828), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1148), .A2(new_n615), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n615), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT60), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n988), .A2(new_n1022), .A3(new_n986), .A4(new_n990), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1061), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n543), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1158), .A3(new_n543), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n615), .A2(KEYINPUT60), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1157), .A2(new_n1159), .B1(new_n1148), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1147), .A2(new_n1151), .A3(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1163));
  AOI21_X1  g738(.A(new_n1137), .B1(new_n1132), .B2(new_n1141), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1145), .A2(new_n1140), .A3(new_n1136), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT123), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1168), .B(new_n1163), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1162), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1150), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1146), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(KEYINPUT121), .B(new_n1146), .C1(new_n1165), .C2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1125), .B(new_n1130), .C1(new_n1170), .C2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1115), .B1(new_n1177), .B2(new_n1093), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1011), .B1(new_n1097), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1007), .A2(new_n1001), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT48), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1003), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n758), .A2(new_n761), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1000), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n826), .A2(new_n828), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1001), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1001), .B1(new_n997), .B2(new_n998), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n992), .A2(new_n986), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT46), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1188), .A2(KEYINPUT46), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT47), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1182), .A2(new_n1186), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1179), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g769(.A1(G227), .A2(new_n461), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n1196), .B1(new_n719), .B2(new_n720), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n676), .B2(new_n683), .ZN(new_n1198));
  NAND4_X1  g772(.A1(new_n925), .A2(new_n976), .A3(new_n1198), .A4(new_n979), .ZN(G225));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n1200));
  XNOR2_X1  g774(.A(G225), .B(new_n1200), .ZN(G308));
endmodule


