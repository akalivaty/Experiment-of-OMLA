

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738;

  BUF_X1 U366 ( .A(n711), .Z(n389) );
  AND2_X1 U367 ( .A1(n738), .A2(n408), .ZN(n407) );
  NOR2_X1 U368 ( .A1(n537), .A2(n538), .ZN(n533) );
  NOR2_X1 U369 ( .A1(n639), .A2(n662), .ZN(n381) );
  INV_X1 U370 ( .A(G953), .ZN(n725) );
  NOR2_X1 U371 ( .A1(n623), .A2(n706), .ZN(n627) );
  INV_X2 U372 ( .A(n379), .ZN(n481) );
  XNOR2_X2 U373 ( .A(G116), .B(KEYINPUT3), .ZN(n379) );
  XNOR2_X2 U374 ( .A(n531), .B(KEYINPUT35), .ZN(n733) );
  XNOR2_X2 U375 ( .A(n722), .B(n410), .ZN(n700) );
  INV_X1 U376 ( .A(n595), .ZN(n674) );
  NAND2_X1 U377 ( .A1(n525), .A2(n673), .ZN(n547) );
  BUF_X1 U378 ( .A(n555), .Z(n600) );
  NOR2_X1 U379 ( .A1(n611), .A2(n706), .ZN(n613) );
  NOR2_X1 U380 ( .A1(n617), .A2(n706), .ZN(n618) );
  AND2_X1 U381 ( .A1(n420), .A2(n419), .ZN(n356) );
  NAND2_X1 U382 ( .A1(n533), .A2(n523), .ZN(n388) );
  XNOR2_X1 U383 ( .A(n426), .B(n425), .ZN(n574) );
  XNOR2_X1 U384 ( .A(n406), .B(KEYINPUT1), .ZN(n525) );
  XNOR2_X1 U385 ( .A(n492), .B(n491), .ZN(n555) );
  XNOR2_X1 U386 ( .A(n362), .B(n501), .ZN(n670) );
  XNOR2_X1 U387 ( .A(n507), .B(n383), .ZN(n411) );
  XNOR2_X1 U388 ( .A(n384), .B(G140), .ZN(n383) );
  XNOR2_X1 U389 ( .A(n357), .B(G101), .ZN(n511) );
  XOR2_X1 U390 ( .A(G137), .B(G131), .Z(n512) );
  XNOR2_X2 U391 ( .A(n516), .B(n512), .ZN(n722) );
  INV_X1 U392 ( .A(G134), .ZN(n455) );
  XNOR2_X1 U393 ( .A(n511), .B(n510), .ZN(n514) );
  XNOR2_X1 U394 ( .A(n441), .B(G146), .ZN(n502) );
  INV_X1 U395 ( .A(KEYINPUT4), .ZN(n441) );
  XNOR2_X1 U396 ( .A(n385), .B(n354), .ZN(n711) );
  AND2_X1 U397 ( .A1(n540), .A2(n347), .ZN(n553) );
  XNOR2_X1 U398 ( .A(n570), .B(KEYINPUT69), .ZN(n585) );
  NAND2_X1 U399 ( .A1(n670), .A2(n569), .ZN(n570) );
  XNOR2_X1 U400 ( .A(n520), .B(G472), .ZN(n548) );
  XNOR2_X1 U401 ( .A(n365), .B(n364), .ZN(n449) );
  INV_X1 U402 ( .A(KEYINPUT8), .ZN(n364) );
  NAND2_X1 U403 ( .A1(n725), .A2(G234), .ZN(n365) );
  NOR2_X1 U404 ( .A1(n576), .A2(n659), .ZN(n396) );
  XOR2_X1 U405 ( .A(G478), .B(n457), .Z(n543) );
  XNOR2_X1 U406 ( .A(n470), .B(n469), .ZN(n541) );
  XNOR2_X1 U407 ( .A(n638), .B(KEYINPUT79), .ZN(n580) );
  INV_X1 U408 ( .A(KEYINPUT65), .ZN(n377) );
  INV_X1 U409 ( .A(n628), .ZN(n382) );
  INV_X1 U410 ( .A(KEYINPUT73), .ZN(n386) );
  XNOR2_X1 U411 ( .A(n515), .B(n519), .ZN(n397) );
  XNOR2_X1 U412 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U413 ( .A(n446), .B(n445), .ZN(n721) );
  XOR2_X1 U414 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n461) );
  XNOR2_X1 U415 ( .A(G131), .B(KEYINPUT97), .ZN(n458) );
  XOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n459) );
  XNOR2_X1 U417 ( .A(n465), .B(G122), .ZN(n405) );
  OR2_X1 U418 ( .A1(n497), .A2(G902), .ZN(n362) );
  XOR2_X1 U419 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n500) );
  XNOR2_X1 U420 ( .A(n721), .B(n403), .ZN(n464) );
  INV_X1 U421 ( .A(G146), .ZN(n403) );
  XNOR2_X1 U422 ( .A(n418), .B(n417), .ZN(n416) );
  XNOR2_X1 U423 ( .A(G137), .B(KEYINPUT24), .ZN(n418) );
  XNOR2_X1 U424 ( .A(KEYINPUT23), .B(G110), .ZN(n417) );
  XNOR2_X1 U425 ( .A(n415), .B(KEYINPUT92), .ZN(n414) );
  XNOR2_X1 U426 ( .A(G119), .B(G128), .ZN(n415) );
  OR2_X2 U427 ( .A1(n604), .A2(n389), .ZN(n419) );
  NAND2_X1 U428 ( .A1(n372), .A2(n370), .ZN(n420) );
  AND2_X1 U429 ( .A1(n359), .A2(n373), .ZN(n372) );
  NAND2_X1 U430 ( .A1(n371), .A2(n378), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n502), .B(n485), .ZN(n440) );
  XNOR2_X1 U432 ( .A(n439), .B(n438), .ZN(n437) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT76), .ZN(n439) );
  XNOR2_X1 U434 ( .A(G125), .B(KEYINPUT17), .ZN(n438) );
  XNOR2_X1 U435 ( .A(n482), .B(n483), .ZN(n707) );
  XNOR2_X1 U436 ( .A(n486), .B(G110), .ZN(n504) );
  INV_X1 U437 ( .A(n419), .ZN(n361) );
  XNOR2_X1 U438 ( .A(n567), .B(KEYINPUT41), .ZN(n692) );
  AND2_X1 U439 ( .A1(n584), .A2(n399), .ZN(n596) );
  AND2_X1 U440 ( .A1(n585), .A2(n400), .ZN(n399) );
  INV_X1 U441 ( .A(n658), .ZN(n400) );
  NOR2_X1 U442 ( .A1(n561), .A2(n568), .ZN(n563) );
  XNOR2_X1 U443 ( .A(n394), .B(KEYINPUT30), .ZN(n561) );
  OR2_X1 U444 ( .A1(n571), .A2(n658), .ZN(n394) );
  INV_X1 U445 ( .A(KEYINPUT108), .ZN(n425) );
  INV_X1 U446 ( .A(n548), .ZN(n680) );
  XNOR2_X1 U447 ( .A(n433), .B(KEYINPUT22), .ZN(n537) );
  AND2_X1 U448 ( .A1(n660), .A2(n435), .ZN(n434) );
  XNOR2_X1 U449 ( .A(n450), .B(n390), .ZN(n453) );
  NAND2_X1 U450 ( .A1(n356), .A2(G478), .ZN(n432) );
  NOR2_X1 U451 ( .A1(G953), .A2(G237), .ZN(n517) );
  OR2_X1 U452 ( .A1(G237), .A2(G902), .ZN(n490) );
  AND2_X1 U453 ( .A1(n737), .A2(n424), .ZN(n423) );
  INV_X1 U454 ( .A(n651), .ZN(n424) );
  NAND2_X1 U455 ( .A1(n421), .A2(n375), .ZN(n374) );
  NAND2_X1 U456 ( .A1(KEYINPUT2), .A2(n377), .ZN(n375) );
  NAND2_X1 U457 ( .A1(n602), .A2(n377), .ZN(n376) );
  AND2_X1 U458 ( .A1(n422), .A2(KEYINPUT65), .ZN(n378) );
  NAND2_X1 U459 ( .A1(n360), .A2(n345), .ZN(n359) );
  INV_X1 U460 ( .A(KEYINPUT67), .ZN(n357) );
  XNOR2_X1 U461 ( .A(n600), .B(n380), .ZN(n659) );
  INV_X1 U462 ( .A(KEYINPUT38), .ZN(n380) );
  NAND2_X1 U463 ( .A1(n528), .A2(n527), .ZN(n413) );
  XNOR2_X1 U464 ( .A(n547), .B(n526), .ZN(n528) );
  NAND2_X1 U465 ( .A1(n368), .A2(n585), .ZN(n367) );
  INV_X1 U466 ( .A(G469), .ZN(n508) );
  XOR2_X1 U467 ( .A(KEYINPUT6), .B(n680), .Z(n527) );
  INV_X1 U468 ( .A(n671), .ZN(n435) );
  NOR2_X1 U469 ( .A1(n543), .A2(n541), .ZN(n660) );
  XNOR2_X1 U470 ( .A(n451), .B(n391), .ZN(n390) );
  INV_X1 U471 ( .A(KEYINPUT7), .ZN(n391) );
  XOR2_X1 U472 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n451) );
  XNOR2_X1 U473 ( .A(n404), .B(n402), .ZN(n608) );
  INV_X1 U474 ( .A(n464), .ZN(n402) );
  XNOR2_X1 U475 ( .A(n466), .B(n405), .ZN(n404) );
  INV_X1 U476 ( .A(KEYINPUT91), .ZN(n384) );
  XOR2_X1 U477 ( .A(G104), .B(G107), .Z(n506) );
  INV_X1 U478 ( .A(KEYINPUT19), .ZN(n428) );
  XOR2_X1 U479 ( .A(n621), .B(n620), .Z(n443) );
  XNOR2_X1 U480 ( .A(n363), .B(n464), .ZN(n497) );
  XNOR2_X1 U481 ( .A(n447), .B(n448), .ZN(n363) );
  XNOR2_X1 U482 ( .A(n416), .B(n414), .ZN(n448) );
  XOR2_X1 U483 ( .A(n608), .B(KEYINPUT59), .Z(n610) );
  XNOR2_X1 U484 ( .A(n440), .B(n437), .ZN(n487) );
  NOR2_X1 U485 ( .A1(n654), .A2(n361), .ZN(n655) );
  XNOR2_X1 U486 ( .A(n572), .B(KEYINPUT42), .ZN(n736) );
  XNOR2_X1 U487 ( .A(n395), .B(n566), .ZN(n734) );
  AND2_X1 U488 ( .A1(n596), .A2(n398), .ZN(n586) );
  INV_X1 U489 ( .A(n600), .ZN(n398) );
  NAND2_X1 U490 ( .A1(n401), .A2(n541), .ZN(n640) );
  INV_X1 U491 ( .A(n543), .ZN(n401) );
  NOR2_X1 U492 ( .A1(n579), .A2(n600), .ZN(n638) );
  INV_X1 U493 ( .A(n541), .ZN(n542) );
  NOR2_X1 U494 ( .A1(n674), .A2(n368), .ZN(n532) );
  INV_X1 U495 ( .A(n640), .ZN(n642) );
  NOR2_X1 U496 ( .A1(n680), .A2(n546), .ZN(n631) );
  XNOR2_X1 U497 ( .A(n432), .B(n351), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n702), .B(n701), .ZN(n703) );
  AND2_X1 U499 ( .A1(n723), .A2(n355), .ZN(n345) );
  XOR2_X1 U500 ( .A(n406), .B(KEYINPUT107), .Z(n346) );
  XNOR2_X1 U501 ( .A(n548), .B(KEYINPUT102), .ZN(n571) );
  INV_X1 U502 ( .A(n571), .ZN(n368) );
  NOR2_X1 U503 ( .A1(n552), .A2(n382), .ZN(n347) );
  AND2_X1 U504 ( .A1(n423), .A2(n594), .ZN(n348) );
  AND2_X1 U505 ( .A1(n423), .A2(KEYINPUT48), .ZN(n349) );
  XOR2_X1 U506 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n350) );
  XOR2_X1 U507 ( .A(n705), .B(KEYINPUT120), .Z(n351) );
  XOR2_X1 U508 ( .A(n615), .B(n614), .Z(n352) );
  XOR2_X1 U509 ( .A(n497), .B(KEYINPUT122), .Z(n353) );
  INV_X1 U510 ( .A(n602), .ZN(n421) );
  XNOR2_X1 U511 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  XOR2_X1 U512 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n354) );
  NAND2_X1 U513 ( .A1(n376), .A2(n374), .ZN(n373) );
  AND2_X1 U514 ( .A1(n421), .A2(n377), .ZN(n355) );
  NOR2_X1 U515 ( .A1(G952), .A2(n725), .ZN(n706) );
  INV_X1 U516 ( .A(n706), .ZN(n430) );
  AND2_X2 U517 ( .A1(n420), .A2(n419), .ZN(n704) );
  XNOR2_X1 U518 ( .A(n413), .B(n529), .ZN(n668) );
  OR2_X1 U519 ( .A1(n711), .A2(n369), .ZN(n371) );
  NAND2_X2 U520 ( .A1(n393), .A2(n392), .ZN(n723) );
  INV_X1 U521 ( .A(n711), .ZN(n360) );
  XNOR2_X1 U522 ( .A(n605), .B(n353), .ZN(n606) );
  XNOR2_X1 U523 ( .A(n358), .B(KEYINPUT121), .ZN(G63) );
  NAND2_X1 U524 ( .A1(n431), .A2(n430), .ZN(n358) );
  XNOR2_X1 U525 ( .A(n367), .B(n366), .ZN(n427) );
  INV_X1 U526 ( .A(KEYINPUT28), .ZN(n366) );
  INV_X1 U527 ( .A(n723), .ZN(n369) );
  NAND2_X1 U528 ( .A1(n668), .A2(n549), .ZN(n412) );
  XNOR2_X1 U529 ( .A(n412), .B(n350), .ZN(n530) );
  XNOR2_X1 U530 ( .A(n616), .B(n352), .ZN(n617) );
  INV_X1 U531 ( .A(KEYINPUT2), .ZN(n422) );
  XNOR2_X1 U532 ( .A(n609), .B(n610), .ZN(n611) );
  XNOR2_X1 U533 ( .A(n516), .B(n397), .ZN(n619) );
  NOR2_X2 U534 ( .A1(n555), .A2(n658), .ZN(n429) );
  XNOR2_X1 U535 ( .A(n429), .B(n428), .ZN(n575) );
  NAND2_X1 U536 ( .A1(n736), .A2(n734), .ZN(n573) );
  NAND2_X1 U537 ( .A1(n593), .A2(n348), .ZN(n393) );
  XNOR2_X2 U538 ( .A(n534), .B(KEYINPUT103), .ZN(n732) );
  XNOR2_X1 U539 ( .A(n381), .B(KEYINPUT47), .ZN(n581) );
  XNOR2_X1 U540 ( .A(n387), .B(n386), .ZN(n554) );
  XNOR2_X2 U541 ( .A(G119), .B(KEYINPUT70), .ZN(n480) );
  NAND2_X1 U542 ( .A1(n553), .A2(n554), .ZN(n385) );
  NAND2_X1 U543 ( .A1(n535), .A2(n738), .ZN(n409) );
  NOR2_X2 U544 ( .A1(n732), .A2(n733), .ZN(n535) );
  NAND2_X1 U545 ( .A1(n407), .A2(n535), .ZN(n387) );
  XNOR2_X2 U546 ( .A(n388), .B(KEYINPUT32), .ZN(n738) );
  INV_X1 U547 ( .A(n524), .ZN(n436) );
  NAND2_X1 U548 ( .A1(n592), .A2(n349), .ZN(n392) );
  NAND2_X1 U549 ( .A1(n565), .A2(n642), .ZN(n395) );
  XNOR2_X1 U550 ( .A(n396), .B(n564), .ZN(n565) );
  XNOR2_X2 U551 ( .A(n503), .B(n502), .ZN(n516) );
  XNOR2_X2 U552 ( .A(n484), .B(n455), .ZN(n503) );
  NAND2_X1 U553 ( .A1(n406), .A2(n673), .ZN(n544) );
  XNOR2_X2 U554 ( .A(n509), .B(n508), .ZN(n406) );
  INV_X1 U555 ( .A(KEYINPUT44), .ZN(n408) );
  NAND2_X1 U556 ( .A1(n409), .A2(KEYINPUT44), .ZN(n540) );
  XNOR2_X1 U557 ( .A(n411), .B(n504), .ZN(n410) );
  NAND2_X1 U558 ( .A1(n436), .A2(n434), .ZN(n433) );
  NOR2_X2 U559 ( .A1(G902), .A2(n700), .ZN(n509) );
  INV_X1 U560 ( .A(n670), .ZN(n538) );
  NAND2_X1 U561 ( .A1(n427), .A2(n346), .ZN(n426) );
  NAND2_X1 U562 ( .A1(n575), .A2(n493), .ZN(n494) );
  XOR2_X1 U563 ( .A(n699), .B(n698), .Z(n442) );
  AND2_X1 U564 ( .A1(n517), .A2(G210), .ZN(n444) );
  XNOR2_X1 U565 ( .A(G113), .B(KEYINPUT5), .ZN(n510) );
  INV_X1 U566 ( .A(n512), .ZN(n513) );
  INV_X1 U567 ( .A(KEYINPUT104), .ZN(n526) );
  XNOR2_X1 U568 ( .A(n518), .B(n444), .ZN(n519) );
  XNOR2_X1 U569 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n529) );
  BUF_X1 U570 ( .A(n668), .Z(n691) );
  INV_X1 U571 ( .A(KEYINPUT39), .ZN(n564) );
  XNOR2_X1 U572 ( .A(n622), .B(n443), .ZN(n623) );
  NAND2_X1 U573 ( .A1(n606), .A2(n430), .ZN(n607) );
  XNOR2_X1 U574 ( .A(n607), .B(KEYINPUT123), .ZN(G66) );
  XOR2_X1 U575 ( .A(G140), .B(KEYINPUT10), .Z(n446) );
  XNOR2_X1 U576 ( .A(G125), .B(KEYINPUT68), .ZN(n445) );
  NAND2_X1 U577 ( .A1(G221), .A2(n449), .ZN(n447) );
  NAND2_X1 U578 ( .A1(G217), .A2(n449), .ZN(n450) );
  XOR2_X1 U579 ( .A(G122), .B(G107), .Z(n479) );
  XNOR2_X1 U580 ( .A(G116), .B(n479), .ZN(n452) );
  XNOR2_X1 U581 ( .A(n453), .B(n452), .ZN(n456) );
  XNOR2_X2 U582 ( .A(G128), .B(KEYINPUT78), .ZN(n454) );
  XNOR2_X2 U583 ( .A(n454), .B(G143), .ZN(n484) );
  XOR2_X1 U584 ( .A(n503), .B(n456), .Z(n705) );
  NOR2_X1 U585 ( .A1(G902), .A2(n705), .ZN(n457) );
  XNOR2_X1 U586 ( .A(n459), .B(n458), .ZN(n463) );
  NAND2_X1 U587 ( .A1(G214), .A2(n517), .ZN(n460) );
  XNOR2_X1 U588 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U589 ( .A(n463), .B(n462), .ZN(n466) );
  XOR2_X1 U590 ( .A(G113), .B(G104), .Z(n478) );
  XNOR2_X1 U591 ( .A(G143), .B(n478), .ZN(n465) );
  NOR2_X1 U592 ( .A1(n608), .A2(G902), .ZN(n470) );
  XOR2_X1 U593 ( .A(KEYINPUT13), .B(KEYINPUT100), .Z(n468) );
  XNOR2_X1 U594 ( .A(KEYINPUT99), .B(G475), .ZN(n467) );
  XNOR2_X1 U595 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U596 ( .A1(G898), .A2(n725), .ZN(n709) );
  NAND2_X1 U597 ( .A1(G234), .A2(G237), .ZN(n471) );
  XNOR2_X1 U598 ( .A(n471), .B(KEYINPUT14), .ZN(n474) );
  NAND2_X1 U599 ( .A1(G902), .A2(n474), .ZN(n472) );
  XNOR2_X1 U600 ( .A(n472), .B(KEYINPUT89), .ZN(n557) );
  NAND2_X1 U601 ( .A1(n709), .A2(n557), .ZN(n473) );
  XNOR2_X1 U602 ( .A(KEYINPUT90), .B(n473), .ZN(n476) );
  NAND2_X1 U603 ( .A1(G952), .A2(n474), .ZN(n689) );
  NOR2_X1 U604 ( .A1(G953), .A2(n689), .ZN(n475) );
  XOR2_X1 U605 ( .A(KEYINPUT88), .B(n475), .Z(n556) );
  NAND2_X1 U606 ( .A1(n476), .A2(n556), .ZN(n493) );
  NAND2_X1 U607 ( .A1(G214), .A2(n490), .ZN(n477) );
  XNOR2_X1 U608 ( .A(KEYINPUT87), .B(n477), .ZN(n658) );
  XOR2_X1 U609 ( .A(n479), .B(n478), .Z(n483) );
  XNOR2_X2 U610 ( .A(n481), .B(n480), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n518), .B(KEYINPUT16), .ZN(n482) );
  XNOR2_X1 U612 ( .A(n484), .B(n707), .ZN(n489) );
  NAND2_X1 U613 ( .A1(G224), .A2(n725), .ZN(n485) );
  XNOR2_X1 U614 ( .A(n511), .B(KEYINPUT71), .ZN(n486) );
  XOR2_X1 U615 ( .A(n487), .B(n504), .Z(n488) );
  XNOR2_X1 U616 ( .A(n489), .B(n488), .ZN(n615) );
  NAND2_X1 U617 ( .A1(n615), .A2(n602), .ZN(n492) );
  NAND2_X1 U618 ( .A1(G210), .A2(n490), .ZN(n491) );
  XNOR2_X1 U619 ( .A(n494), .B(KEYINPUT0), .ZN(n524) );
  NAND2_X1 U620 ( .A1(G234), .A2(n602), .ZN(n495) );
  XNOR2_X1 U621 ( .A(KEYINPUT20), .B(n495), .ZN(n498) );
  NAND2_X1 U622 ( .A1(G221), .A2(n498), .ZN(n496) );
  XNOR2_X1 U623 ( .A(n496), .B(KEYINPUT21), .ZN(n671) );
  NAND2_X1 U624 ( .A1(n498), .A2(G217), .ZN(n499) );
  XNOR2_X1 U625 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U626 ( .A1(G227), .A2(n725), .ZN(n505) );
  XNOR2_X1 U627 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U628 ( .A(n525), .ZN(n595) );
  XOR2_X1 U629 ( .A(KEYINPUT85), .B(n674), .Z(n587) );
  INV_X1 U630 ( .A(n587), .ZN(n522) );
  NOR2_X1 U631 ( .A1(n619), .A2(G902), .ZN(n520) );
  INV_X1 U632 ( .A(n527), .ZN(n583) );
  XNOR2_X1 U633 ( .A(KEYINPUT77), .B(n583), .ZN(n521) );
  NOR2_X1 U634 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U635 ( .A(n524), .ZN(n549) );
  NOR2_X1 U636 ( .A1(n671), .A2(n670), .ZN(n673) );
  AND2_X1 U637 ( .A1(n541), .A2(n543), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n530), .A2(n578), .ZN(n531) );
  NAND2_X1 U639 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U640 ( .A1(n595), .A2(n583), .ZN(n536) );
  NOR2_X1 U641 ( .A1(n537), .A2(n536), .ZN(n539) );
  NAND2_X1 U642 ( .A1(n539), .A2(n538), .ZN(n628) );
  NAND2_X1 U643 ( .A1(n543), .A2(n542), .ZN(n635) );
  INV_X1 U644 ( .A(n635), .ZN(n645) );
  NOR2_X1 U645 ( .A1(n642), .A2(n645), .ZN(n662) );
  XOR2_X1 U646 ( .A(n544), .B(KEYINPUT94), .Z(n562) );
  AND2_X1 U647 ( .A1(n549), .A2(n562), .ZN(n545) );
  XNOR2_X1 U648 ( .A(n545), .B(KEYINPUT95), .ZN(n546) );
  NOR2_X1 U649 ( .A1(n548), .A2(n547), .ZN(n682) );
  NAND2_X1 U650 ( .A1(n682), .A2(n549), .ZN(n550) );
  XNOR2_X1 U651 ( .A(KEYINPUT31), .B(n550), .ZN(n646) );
  NOR2_X1 U652 ( .A1(n631), .A2(n646), .ZN(n551) );
  NOR2_X1 U653 ( .A1(n662), .A2(n551), .ZN(n552) );
  INV_X1 U654 ( .A(n556), .ZN(n560) );
  NAND2_X1 U655 ( .A1(n557), .A2(G953), .ZN(n558) );
  NOR2_X1 U656 ( .A1(G900), .A2(n558), .ZN(n559) );
  NOR2_X1 U657 ( .A1(n560), .A2(n559), .ZN(n568) );
  NAND2_X1 U658 ( .A1(n563), .A2(n562), .ZN(n576) );
  AND2_X1 U659 ( .A1(n645), .A2(n565), .ZN(n651) );
  XOR2_X1 U660 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n566) );
  NOR2_X1 U661 ( .A1(n658), .A2(n659), .ZN(n664) );
  NAND2_X1 U662 ( .A1(n660), .A2(n664), .ZN(n567) );
  NOR2_X1 U663 ( .A1(n671), .A2(n568), .ZN(n569) );
  NAND2_X1 U664 ( .A1(n692), .A2(n574), .ZN(n572) );
  XNOR2_X1 U665 ( .A(n573), .B(KEYINPUT46), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n575), .A2(n574), .ZN(n639) );
  INV_X1 U667 ( .A(n576), .ZN(n577) );
  NAND2_X1 U668 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U669 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U670 ( .A(n582), .B(KEYINPUT75), .ZN(n589) );
  NOR2_X1 U671 ( .A1(n583), .A2(n640), .ZN(n584) );
  XNOR2_X1 U672 ( .A(n586), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n588), .A2(n587), .ZN(n649) );
  NAND2_X1 U674 ( .A1(n589), .A2(n649), .ZN(n590) );
  NOR2_X2 U675 ( .A1(n591), .A2(n590), .ZN(n592) );
  INV_X1 U676 ( .A(KEYINPUT48), .ZN(n594) );
  INV_X1 U677 ( .A(n592), .ZN(n593) );
  XOR2_X1 U678 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n598) );
  NAND2_X1 U679 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U680 ( .A(n598), .B(n597), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U682 ( .A(n601), .B(KEYINPUT106), .ZN(n737) );
  NAND2_X1 U683 ( .A1(n723), .A2(KEYINPUT2), .ZN(n603) );
  XNOR2_X1 U684 ( .A(KEYINPUT82), .B(n603), .ZN(n604) );
  NAND2_X1 U685 ( .A1(G217), .A2(n356), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n704), .A2(G475), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(G60) );
  NAND2_X1 U689 ( .A1(n704), .A2(G210), .ZN(n616) );
  XOR2_X1 U690 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n614) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U692 ( .A1(n704), .A2(G472), .ZN(n622) );
  XOR2_X1 U693 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n621) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT84), .ZN(n620) );
  XOR2_X1 U695 ( .A(KEYINPUT83), .B(KEYINPUT111), .Z(n625) );
  XNOR2_X1 U696 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(G57) );
  XNOR2_X1 U699 ( .A(G101), .B(KEYINPUT112), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(G3) );
  NAND2_X1 U701 ( .A1(n631), .A2(n642), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n630), .B(G104), .ZN(G6) );
  XOR2_X1 U703 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n633) );
  NAND2_X1 U704 ( .A1(n631), .A2(n645), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U706 ( .A(G107), .B(n634), .ZN(G9) );
  NOR2_X1 U707 ( .A1(n635), .A2(n639), .ZN(n637) );
  XNOR2_X1 U708 ( .A(G128), .B(KEYINPUT29), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(G30) );
  XOR2_X1 U710 ( .A(G143), .B(n638), .Z(G45) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U712 ( .A(G146), .B(n641), .Z(G48) );
  XOR2_X1 U713 ( .A(G113), .B(KEYINPUT113), .Z(n644) );
  NAND2_X1 U714 ( .A1(n646), .A2(n642), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(G15) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n647), .B(G116), .ZN(G18) );
  XOR2_X1 U718 ( .A(KEYINPUT37), .B(KEYINPUT114), .Z(n648) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U720 ( .A(G125), .B(n650), .ZN(G27) );
  XOR2_X1 U721 ( .A(G134), .B(n651), .Z(G36) );
  NAND2_X1 U722 ( .A1(n389), .A2(n422), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n652), .B(KEYINPUT80), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n723), .A2(KEYINPUT2), .ZN(n653) );
  XOR2_X1 U725 ( .A(KEYINPUT81), .B(n653), .Z(n654) );
  NAND2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n657), .A2(n725), .ZN(n696) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n666) );
  INV_X1 U730 ( .A(n662), .ZN(n663) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(KEYINPUT116), .ZN(n669) );
  NAND2_X1 U734 ( .A1(n669), .A2(n691), .ZN(n686) );
  AND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U736 ( .A(KEYINPUT49), .B(n672), .ZN(n678) );
  XOR2_X1 U737 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n676) );
  OR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U739 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U743 ( .A(KEYINPUT51), .B(n683), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n684), .A2(n692), .ZN(n685) );
  NAND2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U746 ( .A(KEYINPUT52), .B(n687), .Z(n688) );
  NOR2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U748 ( .A(n690), .B(KEYINPUT117), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U751 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U752 ( .A(n697), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U753 ( .A1(n356), .A2(G469), .ZN(n702) );
  XOR2_X1 U754 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n699) );
  XNOR2_X1 U755 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n700), .B(n442), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n706), .A2(n703), .ZN(G54) );
  XNOR2_X1 U758 ( .A(G101), .B(n707), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n708), .B(G110), .ZN(n710) );
  NOR2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n720) );
  NOR2_X1 U761 ( .A1(G953), .A2(n389), .ZN(n712) );
  XNOR2_X1 U762 ( .A(KEYINPUT125), .B(n712), .ZN(n717) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U765 ( .A1(n714), .A2(G898), .ZN(n715) );
  XNOR2_X1 U766 ( .A(KEYINPUT124), .B(n715), .ZN(n716) );
  NAND2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(KEYINPUT126), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(G69) );
  XOR2_X1 U770 ( .A(n722), .B(n721), .Z(n727) );
  INV_X1 U771 ( .A(n727), .ZN(n724) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(n725), .ZN(n731) );
  XNOR2_X1 U774 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U778 ( .A(n732), .B(G110), .Z(G12) );
  XOR2_X1 U779 ( .A(n733), .B(G122), .Z(G24) );
  XOR2_X1 U780 ( .A(G131), .B(n734), .Z(n735) );
  XNOR2_X1 U781 ( .A(KEYINPUT127), .B(n735), .ZN(G33) );
  XNOR2_X1 U782 ( .A(G137), .B(n736), .ZN(G39) );
  XNOR2_X1 U783 ( .A(G140), .B(n737), .ZN(G42) );
  XNOR2_X1 U784 ( .A(n738), .B(G119), .ZN(G21) );
endmodule

