//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n205), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n223), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  AND2_X1   g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT66), .B1(new_n247), .B2(new_n211), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n252), .A2(new_n253), .A3(G1), .A4(G13), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n248), .A2(new_n251), .A3(G274), .A4(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n248), .A2(new_n254), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n257), .B2(new_n217), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n260), .B2(new_n262), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G97), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT68), .B(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n267), .B(new_n268), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n247), .A2(new_n211), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n258), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI211_X1 g0076(.A(KEYINPUT13), .B(new_n258), .C1(new_n272), .C2(new_n273), .ZN(new_n277));
  OAI21_X1  g0077(.A(G169), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT14), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n274), .B2(new_n275), .ZN(new_n282));
  INV_X1    g0082(.A(new_n277), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n280), .A2(G179), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(G169), .C1(new_n276), .C2(new_n277), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n279), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n216), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT12), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n211), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n288), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n249), .A2(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G68), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G50), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n303), .A2(new_n304), .B1(new_n212), .B2(G68), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n212), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(G77), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n293), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n300), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n280), .A2(G190), .A3(new_n282), .A4(new_n283), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n276), .A2(new_n277), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n313), .B2(G200), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n287), .A2(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n255), .B1(new_n257), .B2(new_n271), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n261), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT67), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(G1698), .A3(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G223), .ZN(new_n325));
  INV_X1    g0125(.A(new_n270), .ZN(new_n326));
  INV_X1    g0126(.A(new_n266), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n326), .A2(G222), .B1(G77), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n316), .B1(new_n329), .B2(new_n273), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G190), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G58), .A2(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n212), .B1(new_n332), .B2(new_n304), .ZN(new_n333));
  INV_X1    g0133(.A(G150), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n303), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT8), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G58), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n306), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n333), .B(new_n335), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n294), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n296), .A2(G50), .A3(new_n297), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G50), .B2(new_n288), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT9), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G200), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n331), .B(new_n347), .C1(new_n348), .C2(new_n330), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT10), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n329), .A2(new_n273), .ZN(new_n351));
  INV_X1    g0151(.A(new_n316), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n346), .B1(new_n353), .B2(G200), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n331), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n353), .A2(G179), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n330), .A2(G169), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n358), .A2(new_n345), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n296), .A2(G77), .A3(new_n297), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n339), .B(KEYINPUT70), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n302), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n340), .B1(G20), .B2(G77), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n294), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n362), .B(new_n368), .C1(new_n307), .C2(new_n289), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n217), .B1(new_n322), .B2(new_n323), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n266), .A2(G232), .A3(new_n269), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n266), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n273), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n256), .A2(G244), .A3(new_n250), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n375), .A2(new_n255), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G169), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(new_n380), .A3(new_n376), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(G200), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n369), .C1(new_n384), .C2(new_n377), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AND4_X1   g0186(.A1(new_n315), .A2(new_n357), .A3(new_n361), .A4(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n222), .A2(new_n216), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n332), .ZN(new_n389));
  INV_X1    g0189(.A(G159), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n303), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT3), .B(G33), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(G20), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n260), .A2(new_n262), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n391), .B1(new_n397), .B2(G68), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n294), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n319), .B2(new_n320), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n396), .B1(new_n400), .B2(KEYINPUT7), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n391), .B1(new_n401), .B2(G68), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n339), .A2(new_n297), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n295), .A2(new_n404), .B1(new_n288), .B2(new_n339), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n269), .A2(G223), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G226), .A2(G1698), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n395), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n259), .A2(new_n218), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n273), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n248), .A2(G232), .A3(new_n250), .A4(new_n254), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n255), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT74), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n255), .A2(new_n416), .A3(KEYINPUT74), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G169), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n380), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n410), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT18), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n407), .A2(new_n427), .A3(new_n408), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n403), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n421), .A2(G200), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n269), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n431), .A2(new_n395), .B1(new_n259), .B2(new_n218), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(new_n273), .B1(new_n417), .B2(new_n418), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(G190), .A3(new_n420), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n426), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n403), .A2(new_n409), .A3(new_n430), .A4(new_n434), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT17), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n348), .B1(new_n433), .B2(new_n420), .ZN(new_n439));
  AND4_X1   g0239(.A1(G190), .A2(new_n415), .A3(new_n419), .A4(new_n420), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n441), .A2(KEYINPUT75), .A3(new_n403), .A4(new_n428), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT76), .A4(new_n442), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n425), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n387), .A2(KEYINPUT77), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT77), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n315), .A2(new_n357), .A3(new_n361), .A4(new_n386), .ZN(new_n450));
  INV_X1    g0250(.A(new_n425), .ZN(new_n451));
  AND4_X1   g0251(.A1(new_n403), .A2(new_n430), .A3(new_n428), .A4(new_n434), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(KEYINPUT75), .B1(new_n437), .B2(KEYINPUT17), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT76), .B1(new_n453), .B2(new_n436), .ZN(new_n454));
  INV_X1    g0254(.A(new_n446), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n449), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G41), .ZN(new_n462));
  INV_X1    g0262(.A(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n256), .A2(KEYINPUT88), .A3(G264), .A4(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(new_n248), .A3(G264), .A4(new_n254), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT88), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n269), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n395), .ZN(new_n472));
  INV_X1    g0272(.A(G294), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n259), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n273), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT89), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n460), .A2(new_n462), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n464), .B(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n256), .A2(G274), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT89), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n470), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n477), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n470), .A2(new_n475), .A3(new_n481), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n484), .A2(new_n380), .B1(new_n378), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n393), .A2(new_n212), .A3(G87), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT87), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT22), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n487), .B2(KEYINPUT22), .ZN(new_n490));
  OR3_X1    g0290(.A1(new_n218), .A2(KEYINPUT22), .A3(G20), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n489), .A2(new_n490), .B1(new_n327), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT23), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n212), .B2(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n372), .A2(KEYINPUT23), .A3(G20), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G116), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n495), .A2(new_n496), .B1(new_n498), .B2(new_n212), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n492), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n493), .B1(new_n492), .B2(new_n499), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n293), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n296), .B1(G1), .B2(new_n259), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT25), .B1(new_n289), .B2(new_n372), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n289), .A2(KEYINPUT25), .A3(new_n372), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n504), .A2(G107), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n486), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n484), .A2(new_n348), .B1(new_n384), .B2(new_n485), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n509), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT90), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n486), .A2(new_n509), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT90), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(new_n515), .C1(new_n509), .C2(new_n511), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  INV_X1    g0318(.A(new_n273), .ZN(new_n519));
  AND2_X1   g0319(.A1(KEYINPUT4), .A2(G244), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n319), .A2(new_n320), .A3(new_n269), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n319), .A2(G250), .A3(G1698), .A4(new_n320), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n393), .A2(new_n269), .A3(G244), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT78), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n393), .A2(new_n269), .A3(KEYINPUT78), .A4(G244), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n519), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n256), .A2(new_n465), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n481), .B1(new_n225), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n518), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n530), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n273), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n533), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT80), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n378), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n288), .A2(G97), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n503), .B2(new_n224), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n372), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  XOR2_X1   g0345(.A(G97), .B(G107), .Z(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(KEYINPUT6), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G20), .B1(G77), .B2(new_n302), .ZN(new_n548));
  INV_X1    g0348(.A(new_n396), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n212), .B1(new_n264), .B2(new_n265), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n392), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n372), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n544), .B1(new_n552), .B2(new_n293), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n537), .A2(new_n538), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(new_n380), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n293), .ZN(new_n557));
  INV_X1    g0357(.A(new_n544), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(G200), .B2(new_n554), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n534), .A2(new_n539), .A3(G190), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n541), .A2(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT21), .ZN(new_n563));
  INV_X1    g0363(.A(G116), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n289), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n503), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(G20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n293), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(KEYINPUT85), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n259), .A2(G97), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n212), .A3(new_n523), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT86), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n570), .A2(new_n573), .A3(new_n212), .A4(new_n523), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(KEYINPUT85), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n566), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n465), .A2(new_n248), .A3(G270), .A4(new_n254), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n269), .A2(G257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n395), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n319), .B2(new_n320), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n273), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n585), .A2(new_n481), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G169), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n563), .B1(new_n582), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(G200), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n582), .B(new_n595), .C1(new_n384), .C2(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n504), .A2(G116), .ZN(new_n597));
  INV_X1    g0397(.A(new_n581), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n565), .B(new_n597), .C1(new_n598), .C2(new_n579), .ZN(new_n599));
  AND4_X1   g0399(.A1(G179), .A2(new_n585), .A3(new_n481), .A4(new_n591), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n599), .A2(KEYINPUT21), .A3(G169), .A4(new_n592), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n594), .A2(new_n596), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n393), .A2(new_n212), .A3(G68), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n212), .B1(new_n268), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G87), .B2(new_n203), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n306), .B2(new_n224), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n293), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n365), .A2(new_n289), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(KEYINPUT82), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT82), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(new_n365), .B2(new_n503), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n219), .B1(new_n459), .B2(G1), .ZN(new_n616));
  OR3_X1    g0416(.A1(new_n459), .A2(G1), .A3(G274), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n256), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(G244), .A2(G1698), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n497), .B1(new_n395), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n393), .A2(new_n269), .A3(G238), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT81), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n393), .A2(new_n269), .A3(KEYINPUT81), .A4(G238), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n618), .B1(new_n625), .B2(new_n519), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n380), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n378), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n615), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n610), .A2(new_n611), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT82), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n612), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(G200), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n503), .A2(new_n218), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(KEYINPUT83), .B1(G190), .B2(new_n627), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT83), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n634), .A2(new_n635), .A3(new_n640), .A4(new_n637), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n630), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n562), .A2(new_n603), .A3(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n458), .A2(new_n517), .A3(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n287), .A2(new_n311), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n314), .A2(new_n312), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n382), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n454), .B2(new_n455), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n451), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n360), .B1(new_n649), .B2(new_n357), .ZN(new_n650));
  INV_X1    g0450(.A(new_n458), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT92), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n559), .B1(new_n554), .B2(G179), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n378), .B2(new_n540), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n642), .A2(new_n652), .A3(KEYINPUT26), .A4(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n654), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT91), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n626), .A2(new_n657), .A3(new_n378), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n626), .B2(new_n378), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n628), .B(new_n615), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n627), .A2(G190), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(new_n634), .A3(new_n635), .A4(new_n637), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n541), .A2(new_n556), .A3(new_n660), .A4(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT92), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n655), .B1(new_n656), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n660), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n541), .A2(new_n556), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n560), .A2(new_n561), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n662), .B1(new_n511), .B2(new_n509), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n602), .A2(new_n594), .A3(new_n601), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n514), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n667), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n666), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n650), .B1(new_n651), .B2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(new_n509), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n249), .A2(new_n212), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G343), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT93), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n517), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n514), .B2(new_n685), .ZN(new_n687));
  INV_X1    g0487(.A(new_n685), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n599), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n603), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n673), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n673), .A2(new_n688), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n517), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n510), .A2(new_n685), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n206), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n209), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n642), .A2(new_n654), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n664), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n664), .B2(new_n663), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n688), .B1(new_n709), .B2(new_n675), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n688), .B1(new_n666), .B2(new_n675), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(KEYINPUT29), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT95), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n600), .A2(new_n477), .A3(new_n483), .A4(new_n627), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT94), .B1(new_n540), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT94), .B(new_n718), .C1(new_n540), .C2(new_n715), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n627), .A2(G179), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n484), .A2(new_n554), .A3(new_n720), .A4(new_n592), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT31), .B1(new_n722), .B2(new_n688), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n714), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n688), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT95), .A3(new_n723), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n643), .A2(new_n513), .A3(new_n516), .A4(new_n685), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n713), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n706), .B1(new_n735), .B2(G1), .ZN(G364));
  INV_X1    g0536(.A(G13), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n249), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n701), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n693), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n691), .ZN(new_n743));
  INV_X1    g0543(.A(new_n741), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n211), .B1(G20), .B2(new_n378), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n212), .A2(new_n380), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n748), .A2(new_n384), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G322), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n748), .A2(new_n348), .A3(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n212), .A2(G179), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n752), .B(new_n758), .C1(G329), .C2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n759), .A2(new_n384), .A3(G200), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n589), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n380), .A2(new_n348), .A3(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n767), .B1(G294), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n748), .A2(new_n384), .A3(new_n348), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n747), .A2(new_n760), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n771), .A2(G326), .B1(G311), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n763), .A2(new_n327), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n771), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n754), .A2(new_n216), .B1(new_n776), .B2(new_n304), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n750), .A2(new_n222), .B1(new_n772), .B2(new_n307), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n766), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n327), .B1(G87), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n765), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n782), .A2(G107), .B1(new_n769), .B2(G97), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n761), .A2(new_n390), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n746), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n745), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n327), .A2(new_n700), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(G355), .B1(new_n564), .B2(new_n700), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n245), .A2(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n700), .A2(new_n393), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G45), .B2(new_n209), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n744), .B(new_n787), .C1(new_n791), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n790), .B(KEYINPUT96), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n691), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n743), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  OR2_X1    g0602(.A1(new_n369), .A2(new_n685), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n385), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n382), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n379), .A2(new_n381), .A3(new_n685), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(KEYINPUT99), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT99), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n385), .A2(new_n803), .B1(new_n381), .B2(new_n379), .ZN(new_n809));
  INV_X1    g0609(.A(new_n806), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n712), .B(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(new_n733), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT100), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n741), .B1(new_n813), .B2(new_n733), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n745), .A2(new_n788), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n753), .A2(G150), .B1(G159), .B2(new_n773), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n776), .C1(new_n822), .C2(new_n750), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n765), .A2(new_n216), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  INV_X1    g0626(.A(new_n769), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n393), .B1(new_n761), .B2(new_n826), .C1(new_n827), .C2(new_n222), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n825), .B(new_n828), .C1(G50), .C2(new_n780), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n765), .A2(new_n218), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n327), .B1(new_n224), .B2(new_n827), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(G107), .C2(new_n780), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n753), .A2(G283), .B1(G116), .B2(new_n773), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n833), .A2(KEYINPUT97), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n749), .A2(G294), .B1(G311), .B2(new_n762), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n589), .B2(new_n776), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(KEYINPUT97), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n824), .A2(new_n829), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n741), .B1(G77), .B2(new_n819), .C1(new_n839), .C2(new_n746), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT98), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n812), .B2(new_n789), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n817), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n738), .A2(new_n249), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n731), .A2(new_n729), .A3(new_n723), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n311), .B(new_n688), .C1(new_n646), .C2(new_n287), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n311), .A2(new_n688), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n315), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n845), .A2(new_n812), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n399), .B1(KEYINPUT16), .B2(new_n398), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n409), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT102), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT102), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n851), .A2(new_n854), .A3(new_n409), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n683), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n456), .A2(KEYINPUT103), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT103), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n447), .B2(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n853), .B(new_n855), .C1(new_n423), .C2(new_n683), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n437), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n424), .A2(new_n437), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  INV_X1    g0666(.A(new_n410), .ZN(new_n867));
  INV_X1    g0667(.A(new_n683), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n410), .A2(KEYINPUT104), .A3(new_n683), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n864), .B1(new_n871), .B2(new_n862), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n861), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n875), .B(new_n872), .C1(new_n858), .C2(new_n860), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n850), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n451), .A2(new_n443), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n869), .A3(new_n870), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n871), .B(new_n862), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n872), .B1(new_n858), .B2(new_n860), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(KEYINPUT38), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n845), .A2(KEYINPUT40), .A3(new_n849), .A4(new_n812), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n879), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n458), .A2(new_n845), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT107), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(G330), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n887), .B2(new_n889), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n645), .A2(new_n688), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT39), .B1(new_n874), .B2(new_n876), .ZN(new_n896));
  XNOR2_X1  g0696(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n885), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n849), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n676), .A2(new_n685), .A3(new_n812), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n806), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n874), .B2(new_n876), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n451), .A2(new_n683), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT106), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT103), .B1(new_n456), .B2(new_n857), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n447), .A2(new_n859), .A3(new_n856), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n873), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n875), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT38), .B(new_n873), .C1(new_n909), .C2(new_n910), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n883), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n913), .A2(new_n915), .A3(new_n897), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n894), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n913), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n904), .B1(new_n919), .B2(new_n902), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n907), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n458), .B(new_n711), .C1(KEYINPUT29), .C2(new_n712), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n650), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  AOI21_X1  g0725(.A(new_n844), .B1(new_n893), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n893), .B2(new_n925), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n547), .B(KEYINPUT101), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT35), .ZN(new_n929));
  OAI211_X1 g0729(.A(G116), .B(new_n213), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n929), .B2(new_n928), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT36), .Z(new_n932));
  NOR3_X1   g0732(.A1(new_n388), .A2(new_n209), .A3(new_n307), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n216), .A2(G50), .ZN(new_n934));
  OAI211_X1 g0734(.A(G1), .B(new_n737), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n927), .A2(new_n932), .A3(new_n935), .ZN(G367));
  AND2_X1   g0736(.A1(new_n237), .A2(new_n795), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n791), .B1(new_n206), .B2(new_n365), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n741), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n772), .A2(new_n764), .B1(new_n761), .B2(new_n755), .ZN(new_n940));
  XNOR2_X1  g0740(.A(KEYINPUT110), .B(G311), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n750), .A2(new_n589), .B1(new_n776), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n766), .A2(new_n564), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n940), .B(new_n942), .C1(KEYINPUT46), .C2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT111), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n765), .A2(new_n224), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n395), .B1(new_n754), .B2(new_n473), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n947), .B(new_n948), .C1(G107), .C2(new_n769), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n944), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT112), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT112), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n266), .B1(new_n821), .B2(new_n761), .C1(new_n754), .C2(new_n390), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n749), .A2(G150), .B1(G50), .B2(new_n773), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n822), .B2(new_n776), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n827), .A2(new_n216), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n222), .A2(new_n766), .B1(new_n765), .B2(new_n307), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT113), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n951), .A2(new_n952), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT47), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n939), .B1(new_n961), .B2(new_n745), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT114), .Z(new_n963));
  AOI21_X1  g0763(.A(new_n685), .B1(new_n634), .B2(new_n637), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n667), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n964), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n660), .A3(new_n662), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n963), .B1(new_n799), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n562), .B1(new_n553), .B2(new_n685), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n654), .A2(new_n688), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n698), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n698), .A2(new_n974), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n694), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n696), .B1(new_n687), .B2(new_n695), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n693), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n976), .A2(new_n982), .A3(new_n979), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n984), .A2(new_n735), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(new_n735), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n701), .B(KEYINPUT41), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n739), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT43), .B1(new_n968), .B2(KEYINPUT108), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(KEYINPUT108), .B2(new_n968), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n696), .A2(new_n973), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT42), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n510), .A2(new_n669), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n688), .B1(new_n998), .B2(new_n668), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  MUX2_X1   g0800(.A(new_n995), .B(new_n993), .S(new_n1000), .Z(new_n1001));
  NAND2_X1  g0801(.A1(new_n981), .A2(new_n974), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n970), .B1(new_n991), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(G387));
  NAND2_X1  g0805(.A1(new_n986), .A2(new_n735), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n701), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n986), .A2(new_n735), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n687), .A2(new_n799), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n363), .A2(new_n304), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n703), .B(new_n459), .C1(new_n216), .C2(new_n307), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n795), .B1(new_n233), .B2(new_n459), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n703), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n792), .A2(new_n1015), .B1(new_n372), .B2(new_n700), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(KEYINPUT115), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n791), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT115), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n741), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n754), .A2(new_n941), .B1(new_n776), .B2(new_n751), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(KEYINPUT116), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(KEYINPUT116), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n749), .A2(G317), .B1(G303), .B2(new_n773), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT48), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(KEYINPUT48), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n780), .A2(G294), .B1(new_n769), .B2(G283), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n765), .A2(new_n564), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n393), .B(new_n1033), .C1(G326), .C2(new_n762), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n395), .B(new_n947), .C1(G150), .C2(new_n762), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n749), .A2(G50), .B1(G68), .B2(new_n773), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n339), .A2(new_n753), .B1(new_n771), .B2(G159), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n780), .A2(G77), .B1(new_n366), .B2(new_n769), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1020), .B1(new_n1041), .B2(new_n745), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n986), .A2(new_n740), .B1(new_n1010), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1009), .A2(new_n1043), .ZN(G393));
  NAND2_X1  g0844(.A1(new_n980), .A2(new_n981), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n976), .A2(new_n694), .A3(new_n979), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n1006), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n701), .A3(new_n988), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1045), .A2(new_n740), .A3(new_n1046), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n973), .A2(new_n790), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n754), .A2(new_n589), .B1(new_n761), .B2(new_n751), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G294), .B2(new_n773), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n266), .B1(G107), .B2(new_n782), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n780), .A2(G283), .B1(new_n769), .B2(G116), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n749), .A2(G311), .B1(new_n771), .B2(G317), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n749), .A2(G159), .B1(new_n771), .B2(G150), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n827), .A2(new_n307), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n830), .B(new_n1061), .C1(G68), .C2(new_n780), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n363), .A2(new_n773), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n393), .B1(new_n761), .B2(new_n822), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n753), .B2(G50), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1056), .A2(new_n1058), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n745), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n795), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n791), .B1(new_n224), .B2(new_n206), .C1(new_n241), .C2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1051), .A2(new_n741), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n1071), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1049), .B1(new_n1073), .B2(new_n1074), .ZN(G390));
  AND4_X1   g0875(.A1(G330), .A2(new_n845), .A3(new_n812), .A4(new_n849), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n810), .B1(new_n712), .B2(new_n812), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n895), .B1(new_n1078), .B2(new_n900), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n896), .A2(new_n898), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n913), .A2(new_n915), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n810), .B1(new_n710), .B2(new_n812), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n895), .C1(new_n900), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1077), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n732), .A2(G330), .A3(new_n812), .A4(new_n849), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1080), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n845), .A2(G330), .A3(new_n812), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n900), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1086), .A2(new_n1082), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n732), .A2(G330), .A3(new_n812), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1076), .B1(new_n1092), .B2(new_n900), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1093), .B2(new_n1078), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n845), .A2(G330), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n458), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1096), .B(new_n650), .C1(new_n651), .C2(new_n713), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1088), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n1087), .A3(new_n1085), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n701), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n896), .A2(new_n898), .A3(new_n788), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n741), .B1(new_n339), .B2(new_n819), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n750), .A2(new_n564), .B1(new_n761), .B2(new_n473), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G283), .B2(new_n771), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n825), .B(new_n1061), .C1(G87), .C2(new_n780), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n753), .A2(G107), .B1(G97), .B2(new_n773), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1107), .A2(new_n327), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n750), .A2(new_n826), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n327), .B(new_n1111), .C1(G125), .C2(new_n762), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n773), .A2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n753), .A2(G137), .B1(new_n771), .B2(G128), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n782), .A2(G50), .B1(new_n769), .B2(G159), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n780), .A2(G150), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT53), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1110), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1105), .B1(new_n1121), .B2(new_n745), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1104), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT118), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1085), .A2(new_n740), .A3(new_n1087), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1124), .A2(new_n1125), .A3(KEYINPUT119), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT119), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1103), .B1(new_n1126), .B2(new_n1127), .ZN(G378));
  NAND2_X1  g0928(.A1(new_n395), .A2(new_n463), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1129), .B(new_n956), .C1(new_n366), .C2(new_n773), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n222), .B2(new_n765), .C1(new_n307), .C2(new_n766), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n750), .A2(new_n372), .B1(new_n761), .B2(new_n764), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n754), .A2(new_n224), .B1(new_n776), .B2(new_n564), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT58), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n753), .A2(G132), .B1(new_n771), .B2(G125), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n749), .A2(G128), .B1(G137), .B2(new_n773), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n780), .A2(new_n1114), .B1(new_n769), .B2(G150), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n782), .A2(G159), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G33), .B(G41), .C1(new_n762), .C2(G124), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1134), .A2(KEYINPUT58), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1129), .B(new_n304), .C1(G33), .C2(G41), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1135), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n745), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n744), .B1(new_n304), .B2(new_n818), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n357), .A2(new_n361), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n345), .A2(new_n868), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT120), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1152), .B(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1148), .B(new_n1149), .C1(new_n1155), .C2(new_n789), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT122), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n907), .A2(new_n921), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1155), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT40), .B1(new_n919), .B2(new_n850), .ZN(new_n1161));
  OAI21_X1  g0961(.A(G330), .B1(new_n885), .B2(new_n886), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT121), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT121), .ZN(new_n1164));
  INV_X1    g0964(.A(G330), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n886), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1081), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n879), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1160), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1159), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1161), .A2(new_n1162), .A3(KEYINPUT121), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1164), .B1(new_n879), .B2(new_n1167), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1155), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n1170), .C1(new_n922), .C2(KEYINPUT122), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1157), .B1(new_n1177), .B2(new_n740), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1102), .A2(new_n1098), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n922), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1175), .A2(new_n921), .A3(new_n907), .A4(new_n1170), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1080), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1099), .A2(new_n1184), .A3(new_n1084), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1097), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n701), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1178), .B1(new_n1180), .B2(new_n1187), .ZN(G375));
  NAND2_X1  g0988(.A1(new_n900), .A2(new_n788), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n741), .B1(G68), .B2(new_n819), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT123), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n564), .A2(new_n754), .B1(new_n750), .B2(new_n764), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G107), .B2(new_n773), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n771), .A2(G294), .B1(G303), .B2(new_n762), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n327), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n782), .A2(G77), .B1(new_n366), .B2(new_n769), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n224), .B2(new_n766), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n749), .A2(G137), .B1(G128), .B2(new_n762), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n826), .B2(new_n776), .C1(new_n754), .C2(new_n1113), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n780), .A2(G159), .B1(new_n769), .B2(G50), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n395), .B1(new_n773), .B2(G150), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n222), .C2(new_n765), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1195), .A2(new_n1197), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1191), .B1(new_n1203), .B2(new_n745), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1094), .A2(new_n740), .B1(new_n1189), .B2(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1101), .A2(new_n990), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1097), .B(new_n1091), .C1(new_n1093), .C2(new_n1078), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1205), .B1(new_n1206), .B2(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(new_n1074), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1072), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1009), .A2(new_n801), .A3(new_n1043), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(G384), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .A4(new_n1049), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(G387), .A2(G381), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(G375), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1103), .A2(new_n1125), .A3(new_n1124), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(G407));
  INV_X1    g1019(.A(G343), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(G213), .A3(new_n1220), .A4(new_n1218), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(new_n1221), .A3(G213), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT124), .Z(G409));
  OAI211_X1 g1023(.A(G378), .B(new_n1178), .C1(new_n1180), .C2(new_n1187), .ZN(new_n1224));
  AOI221_X4 g1024(.A(new_n990), .B1(new_n1098), .B2(new_n1102), .C1(new_n1172), .C2(new_n1176), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1156), .B1(new_n1183), .B2(new_n739), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1218), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1220), .A2(G213), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  OAI211_X1 g1031(.A(KEYINPUT125), .B(new_n1207), .C1(new_n1101), .C2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1231), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n1208), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n702), .B1(new_n1208), .B2(KEYINPUT60), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1232), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1237), .A2(G384), .A3(new_n1205), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G384), .B1(new_n1237), .B2(new_n1205), .ZN(new_n1239));
  INV_X1    g1039(.A(G2897), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1238), .A2(new_n1239), .B1(new_n1240), .B2(new_n1229), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1205), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1214), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1237), .A2(G384), .A3(new_n1205), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1229), .A2(new_n1240), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT126), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1241), .A2(new_n1246), .A3(KEYINPUT126), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1230), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT62), .B1(new_n1230), .B2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1224), .A2(new_n1227), .B1(G213), .B2(new_n1220), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n801), .B1(new_n1009), .B2(new_n1043), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1211), .B(new_n1049), .C1(new_n1213), .C2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1261), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G390), .A2(new_n1212), .A3(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1262), .A2(new_n1004), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1004), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1253), .A2(new_n1260), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1228), .A2(KEYINPUT63), .A3(new_n1229), .A4(new_n1254), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT63), .B1(new_n1257), .B2(new_n1254), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(new_n1253), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1229), .A2(new_n1228), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT61), .B1(new_n1275), .B2(new_n1250), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT127), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1267), .B1(new_n1273), .B2(new_n1277), .ZN(G405));
  NAND2_X1  g1078(.A1(G375), .A2(new_n1218), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1224), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(new_n1254), .Z(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1269), .ZN(G402));
endmodule


