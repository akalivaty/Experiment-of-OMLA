//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT65), .B(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(KEYINPUT65), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(new_n473), .A3(new_n467), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n465), .A2(new_n480), .ZN(G160));
  NAND3_X1  g056(.A1(new_n478), .A2(G2105), .A3(new_n467), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  INV_X1    g059(.A(new_n479), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT67), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n473), .A2(KEYINPUT68), .A3(G114), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n478), .A2(G126), .A3(G2105), .A4(new_n467), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR4_X1   g074(.A1(new_n470), .A2(KEYINPUT4), .A3(new_n499), .A4(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n478), .A2(G138), .A3(new_n473), .A4(new_n467), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n502), .B2(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n498), .B1(new_n503), .B2(new_n505), .ZN(G164));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(new_n514), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(G166));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n521), .A2(G51), .B1(new_n509), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(KEYINPUT71), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(KEYINPUT71), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(new_n521), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n518), .A2(G90), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n525), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  OAI211_X1 g119(.A(G43), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n545));
  OAI211_X1 g120(.A(G81), .B(new_n509), .C1(new_n515), .C2(new_n516), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT72), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n507), .A2(new_n508), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n549), .A2(new_n550), .B1(new_n524), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT74), .Z(G188));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n507), .A2(new_n566), .A3(new_n508), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(G78), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n518), .A2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n573));
  NAND2_X1  g148(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n527), .B(new_n578), .ZN(G303));
  NAND2_X1  g154(.A1(new_n518), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n521), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT78), .ZN(G288));
  OAI211_X1 g159(.A(G86), .B(new_n509), .C1(new_n515), .C2(new_n516), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n586), .B2(new_n525), .C1(new_n520), .C2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n552), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n518), .A2(G85), .B1(new_n524), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n521), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G301), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n517), .A2(KEYINPUT79), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT79), .B1(new_n517), .B2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n521), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n565), .A2(new_n567), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n605), .B2(new_n511), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT80), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n596), .B1(new_n610), .B2(new_n595), .ZN(G284));
  AOI21_X1  g186(.A(new_n596), .B1(new_n610), .B2(new_n595), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n576), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n576), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n610), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n483), .A2(G123), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n473), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G135), .B2(new_n485), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT82), .Z(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NOR3_X1   g203(.A1(new_n470), .A2(new_n462), .A3(G2105), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n631), .B1(KEYINPUT81), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(KEYINPUT81), .ZN(new_n634));
  MUX2_X1   g209(.A(new_n633), .B(new_n631), .S(new_n634), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT83), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT17), .Z(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  INV_X1    g234(.A(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(new_n654), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n658), .B(new_n659), .C1(new_n657), .C2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n654), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  INV_X1    g259(.A(G34), .ZN(new_n685));
  AOI21_X1  g260(.A(G29), .B1(new_n685), .B2(KEYINPUT24), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(KEYINPUT24), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G160), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G2084), .ZN(new_n691));
  INV_X1    g266(.A(G104), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n692), .A2(new_n473), .A3(KEYINPUT90), .ZN(new_n693));
  AOI21_X1  g268(.A(KEYINPUT90), .B1(new_n692), .B2(new_n473), .ZN(new_n694));
  OAI221_X1 g269(.A(G2104), .B1(G116), .B2(new_n473), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G140), .ZN(new_n696));
  INV_X1    g271(.A(G128), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n695), .B1(new_n479), .B2(new_n696), .C1(new_n697), .C2(new_n482), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n689), .A2(G26), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT91), .B(G2067), .ZN(new_n703));
  OAI22_X1  g278(.A1(new_n690), .A2(new_n691), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT25), .Z(new_n706));
  INV_X1    g281(.A(G139), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n706), .B1(new_n479), .B2(new_n707), .C1(new_n708), .C2(new_n473), .ZN(new_n709));
  MUX2_X1   g284(.A(G33), .B(new_n709), .S(G29), .Z(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G2072), .Z(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NOR2_X1   g288(.A1(G171), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G5), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n689), .A2(G32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n485), .A2(G141), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n483), .A2(G129), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT26), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n463), .A2(G105), .ZN(new_n722));
  NOR4_X1   g297(.A1(new_n718), .A2(new_n719), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n689), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n711), .B1(new_n712), .B2(new_n715), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n704), .B(new_n727), .C1(new_n702), .C2(new_n703), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n726), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n715), .A2(new_n712), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n690), .A2(new_n691), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(KEYINPUT97), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n713), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n555), .B2(new_n713), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G11), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT94), .B(G28), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(new_n689), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n737), .B1(new_n739), .B2(new_n741), .C1(new_n627), .C2(new_n689), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n728), .A2(new_n733), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n713), .A2(G20), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT23), .Z(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G299), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n689), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n689), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT29), .Z(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n749), .B1(new_n753), .B2(G2090), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n713), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n713), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G1966), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT96), .ZN(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n752), .A2(new_n759), .B1(G1966), .B2(new_n756), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n754), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G27), .A2(G29), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G164), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT98), .B(G2078), .Z(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n732), .A2(KEYINPUT97), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n744), .A2(new_n761), .A3(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G24), .B(G290), .S(G16), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT86), .ZN(new_n771));
  INV_X1    g346(.A(G1986), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n689), .A2(G25), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n485), .A2(G131), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n483), .A2(G119), .ZN(new_n777));
  OR2_X1    g352(.A1(G95), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(new_n689), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT35), .B(G1991), .Z(new_n783));
  XOR2_X1   g358(.A(new_n782), .B(new_n783), .Z(new_n784));
  AND2_X1   g359(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n773), .A2(new_n774), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n713), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n713), .ZN(new_n788));
  INV_X1    g363(.A(G1971), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n713), .A2(G23), .ZN(new_n791));
  INV_X1    g366(.A(new_n583), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n713), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G6), .B(G305), .S(G16), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n790), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n786), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n769), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n713), .A2(G4), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n610), .B2(new_n713), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT89), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n808), .A2(new_n813), .ZN(G311));
  INV_X1    g389(.A(G311), .ZN(G150));
  NAND2_X1  g390(.A1(new_n610), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(new_n525), .ZN(new_n819));
  OAI211_X1 g394(.A(G55), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n820));
  OAI211_X1 g395(.A(G93), .B(new_n509), .C1(new_n515), .C2(new_n516), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(KEYINPUT100), .B1(new_n555), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n554), .A2(new_n524), .ZN(new_n824));
  INV_X1    g399(.A(new_n550), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT72), .B1(new_n545), .B2(new_n546), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n828));
  INV_X1    g403(.A(new_n822), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(KEYINPUT99), .B1(new_n827), .B2(new_n829), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n555), .A2(new_n833), .A3(new_n822), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n817), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n822), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT101), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  OR2_X1    g418(.A1(new_n840), .A2(new_n843), .ZN(G145));
  NAND2_X1  g419(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n845));
  INV_X1    g420(.A(new_n500), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n505), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n498), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n723), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n780), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n483), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n473), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G142), .B2(new_n485), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(new_n630), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n698), .B(KEYINPUT102), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n709), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n851), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n627), .B(new_n490), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G160), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n861), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g441(.A1(new_n822), .A2(new_n595), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n609), .A2(G299), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n576), .A2(new_n602), .A3(new_n608), .A4(new_n607), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n868), .A2(KEYINPUT41), .A3(new_n869), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(new_n868), .B2(new_n869), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n618), .B(new_n836), .ZN(new_n875));
  MUX2_X1   g450(.A(new_n871), .B(new_n874), .S(new_n875), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n527), .B(new_n583), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(G290), .B(G305), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G290), .B(G305), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT42), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n880), .A2(KEYINPUT103), .A3(new_n882), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n880), .B2(new_n882), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n887), .B2(KEYINPUT42), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n876), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n867), .B1(new_n889), .B2(new_n595), .ZN(G295));
  OAI21_X1  g465(.A(new_n867), .B1(new_n889), .B2(new_n595), .ZN(G331));
  OAI211_X1 g466(.A(G171), .B(new_n530), .C1(new_n535), .C2(new_n536), .ZN(new_n892));
  NAND2_X1  g467(.A1(G286), .A2(G301), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n836), .A2(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n823), .A2(new_n830), .B1(new_n832), .B2(new_n834), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(KEYINPUT104), .A3(new_n897), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n900), .A2(new_n874), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n898), .A3(KEYINPUT105), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n896), .A2(KEYINPUT105), .A3(new_n897), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n870), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n906), .B2(new_n886), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n887), .B1(new_n902), .B2(new_n905), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n836), .A2(new_n894), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n901), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n871), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n903), .A2(new_n904), .A3(new_n874), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n911), .B1(new_n918), .B2(new_n887), .ZN(new_n919));
  AOI211_X1 g494(.A(KEYINPUT106), .B(new_n886), .C1(new_n916), .C2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n907), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n910), .B1(KEYINPUT43), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n921), .B2(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n907), .A2(KEYINPUT107), .A3(new_n927), .A4(new_n908), .ZN(new_n928));
  INV_X1    g503(.A(new_n905), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n900), .A2(new_n874), .A3(new_n901), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n886), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n908), .A3(new_n927), .A4(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n925), .A2(new_n926), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n926), .B1(new_n925), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n924), .B1(new_n937), .B2(new_n938), .ZN(G397));
  XOR2_X1   g514(.A(KEYINPUT109), .B(G1384), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n849), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G40), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n465), .A2(new_n943), .A3(new_n480), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n723), .B(G1996), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n698), .B(G2067), .Z(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n780), .B(new_n783), .Z(new_n951));
  OAI21_X1  g526(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n592), .A2(new_n772), .A3(new_n593), .ZN(new_n953));
  NAND2_X1  g528(.A1(G290), .A2(G1986), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT110), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT111), .Z(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(G164), .B2(G1384), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT4), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n504), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n962), .A2(new_n963), .A3(new_n500), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT112), .B(new_n961), .C1(new_n964), .C2(new_n498), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n849), .A2(new_n961), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n944), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G2078), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(KEYINPUT53), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G160), .A2(G40), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(KEYINPUT50), .B2(new_n967), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n960), .A2(new_n965), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n712), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n849), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n968), .B1(G164), .B2(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n944), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n982), .B2(G2078), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n972), .A2(new_n978), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(G171), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n942), .A2(new_n979), .A3(G2078), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n944), .A3(new_n980), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n978), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(G171), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n990));
  INV_X1    g565(.A(G1966), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n966), .B2(new_n969), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n974), .A2(new_n976), .A3(new_n691), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(G168), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G8), .ZN(new_n995));
  AOI21_X1  g570(.A(G168), .B1(new_n992), .B2(new_n993), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n998), .A3(G8), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n989), .A2(new_n990), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT112), .B1(new_n849), .B2(new_n961), .ZN(new_n1005));
  NOR3_X1   g580(.A1(G164), .A2(new_n959), .A3(G1384), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT50), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n975), .B(new_n961), .C1(new_n964), .C2(new_n498), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n849), .A2(KEYINPUT116), .A3(new_n975), .A4(new_n961), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1012), .A3(new_n944), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(KEYINPUT117), .ZN(new_n1014));
  AOI21_X1  g589(.A(G2090), .B1(new_n1013), .B2(KEYINPUT117), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1014), .A2(new_n1015), .B1(new_n789), .B2(new_n982), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1004), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n960), .A2(new_n965), .A3(new_n944), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  XNOR2_X1  g596(.A(G305), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1024), .A3(KEYINPUT115), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  OR2_X1    g601(.A1(G305), .A2(G1981), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(G305), .A2(G1981), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1023), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1022), .A2(KEYINPUT49), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1019), .A2(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1026), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1025), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT114), .B1(new_n792), .B2(G1976), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1020), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G288), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1020), .A2(new_n1038), .A3(new_n1036), .A4(new_n1040), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1035), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n982), .A2(new_n789), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n977), .B2(G2090), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1003), .A2(new_n1046), .A3(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT113), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1003), .A2(new_n1046), .A3(new_n1049), .A4(G8), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1044), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n988), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT125), .B1(new_n988), .B2(G171), .ZN(new_n1053));
  OAI221_X1 g628(.A(KEYINPUT54), .B1(G171), .B2(new_n984), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1000), .A2(new_n1018), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT119), .B1(new_n572), .B2(new_n575), .ZN(new_n1056));
  INV_X1    g631(.A(new_n574), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n573), .B(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT57), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1058), .A2(new_n1061), .A3(new_n571), .A4(new_n570), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1056), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n960), .A2(new_n965), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n973), .B1(new_n1066), .B2(KEYINPUT50), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1956), .B1(new_n1067), .B2(new_n1012), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT56), .B(G2072), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT120), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n980), .A2(new_n981), .A3(new_n944), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1065), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1013), .A2(new_n748), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1065), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1073), .A2(new_n1076), .A3(KEYINPUT61), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT61), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  NAND2_X1  g656(.A1(new_n1019), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1996), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n980), .A2(new_n981), .A3(new_n1083), .A4(new_n944), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1082), .A2(KEYINPUT121), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT121), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n555), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1082), .A2(KEYINPUT121), .A3(new_n1084), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT122), .A3(new_n555), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1089), .A2(new_n1095), .A3(KEYINPUT59), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1087), .A2(new_n1088), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1079), .A2(new_n1080), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1075), .B1(new_n1074), .B2(new_n1071), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1072), .B(new_n1065), .C1(new_n1013), .C2(new_n748), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1073), .A2(new_n1076), .A3(KEYINPUT61), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1098), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT122), .B1(new_n1094), .B2(new_n555), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT123), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1019), .A2(G2067), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n977), .B2(new_n812), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  OR3_X1    g688(.A1(new_n1112), .A2(KEYINPUT124), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n609), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT124), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT124), .B(new_n609), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1099), .A2(new_n1109), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1111), .A2(new_n609), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1076), .B1(new_n1101), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1055), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1017), .B(G286), .C1(new_n992), .C2(new_n993), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1046), .A2(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1004), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1051), .A2(KEYINPUT63), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1051), .A2(new_n1018), .A3(new_n1125), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(KEYINPUT63), .ZN(new_n1130));
  AOI211_X1 g705(.A(G1976), .B(G288), .C1(new_n1025), .C2(new_n1034), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1020), .B1(new_n1131), .B2(new_n1028), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1044), .ZN(new_n1134));
  INV_X1    g709(.A(new_n985), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1051), .A2(new_n1018), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n997), .A2(new_n1137), .A3(new_n999), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n997), .B2(new_n999), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1134), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1130), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n958), .B1(new_n1124), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n946), .A2(KEYINPUT46), .A3(new_n1083), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n945), .B2(G1996), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n723), .A2(new_n948), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1144), .B(new_n1146), .C1(new_n945), .C2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT47), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n781), .A2(new_n783), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT126), .Z(new_n1151));
  OAI22_X1  g726(.A1(new_n950), .A2(new_n1151), .B1(G2067), .B2(new_n698), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1152), .A2(new_n946), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n952), .B(KEYINPUT127), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n945), .A2(new_n953), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n1155), .B(KEYINPUT48), .Z(new_n1156));
  AOI211_X1 g731(.A(new_n1149), .B(new_n1153), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1143), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g733(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n1160), .A2(new_n922), .A3(new_n865), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


