

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  AND2_X2 U322 ( .A1(n450), .A2(n530), .ZN(n451) );
  XNOR2_X1 U323 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U324 ( .A(n327), .B(n326), .ZN(n575) );
  XNOR2_X1 U325 ( .A(n451), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U326 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U327 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U328 ( .A(G141GAT), .B(G22GAT), .Z(n332) );
  XOR2_X1 U329 ( .A(G78GAT), .B(G148GAT), .Z(n291) );
  XNOR2_X1 U330 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n290) );
  XNOR2_X1 U331 ( .A(n291), .B(n290), .ZN(n317) );
  XOR2_X1 U332 ( .A(n332), .B(n317), .Z(n293) );
  NAND2_X1 U333 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U335 ( .A(n294), .B(KEYINPUT92), .Z(n298) );
  XOR2_X1 U336 ( .A(G204GAT), .B(G211GAT), .Z(n296) );
  XNOR2_X1 U337 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n396) );
  XNOR2_X1 U339 ( .A(n396), .B(KEYINPUT88), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U341 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n300) );
  XNOR2_X1 U342 ( .A(G50GAT), .B(KEYINPUT94), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U344 ( .A(n302), .B(n301), .Z(n312) );
  XOR2_X1 U345 ( .A(G155GAT), .B(KEYINPUT3), .Z(n304) );
  XNOR2_X1 U346 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U348 ( .A(n305), .B(KEYINPUT89), .Z(n307) );
  XNOR2_X1 U349 ( .A(KEYINPUT2), .B(G162GAT), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n307), .B(n306), .ZN(n425) );
  XOR2_X1 U351 ( .A(KEYINPUT93), .B(KEYINPUT22), .Z(n309) );
  XNOR2_X1 U352 ( .A(G197GAT), .B(KEYINPUT24), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n425), .B(n310), .ZN(n311) );
  XNOR2_X1 U355 ( .A(n312), .B(n311), .ZN(n464) );
  XOR2_X1 U356 ( .A(KEYINPUT13), .B(G57GAT), .Z(n374) );
  XOR2_X1 U357 ( .A(KEYINPUT73), .B(G85GAT), .Z(n314) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(KEYINPUT72), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n316) );
  INV_X1 U360 ( .A(G92GAT), .ZN(n315) );
  XNOR2_X1 U361 ( .A(n316), .B(n315), .ZN(n361) );
  XOR2_X1 U362 ( .A(G176GAT), .B(G64GAT), .Z(n402) );
  XNOR2_X1 U363 ( .A(n361), .B(n402), .ZN(n319) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XOR2_X1 U365 ( .A(n435), .B(n317), .Z(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n374), .B(n320), .ZN(n327) );
  XOR2_X1 U368 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n322) );
  NAND2_X1 U369 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U371 ( .A(KEYINPUT74), .B(n323), .Z(n325) );
  XOR2_X1 U372 ( .A(G204GAT), .B(KEYINPUT31), .Z(n324) );
  INV_X1 U373 ( .A(KEYINPUT64), .ZN(n328) );
  XNOR2_X1 U374 ( .A(n575), .B(n328), .ZN(n329) );
  XNOR2_X1 U375 ( .A(n329), .B(KEYINPUT41), .ZN(n498) );
  XOR2_X1 U376 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n331) );
  XNOR2_X1 U377 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U379 ( .A(KEYINPUT65), .B(G113GAT), .Z(n334) );
  XOR2_X1 U380 ( .A(G15GAT), .B(G1GAT), .Z(n375) );
  XNOR2_X1 U381 ( .A(n332), .B(n375), .ZN(n333) );
  XNOR2_X1 U382 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U383 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U384 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U385 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U386 ( .A(n339), .B(KEYINPUT69), .Z(n342) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(G197GAT), .ZN(n340) );
  XOR2_X1 U388 ( .A(n340), .B(G8GAT), .Z(n407) );
  XOR2_X1 U389 ( .A(n407), .B(KEYINPUT68), .Z(n341) );
  XNOR2_X1 U390 ( .A(n342), .B(n341), .ZN(n347) );
  XOR2_X1 U391 ( .A(G29GAT), .B(KEYINPUT8), .Z(n344) );
  XNOR2_X1 U392 ( .A(G43GAT), .B(G36GAT), .ZN(n343) );
  XNOR2_X1 U393 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U394 ( .A(G50GAT), .B(KEYINPUT7), .Z(n345) );
  XOR2_X1 U395 ( .A(n346), .B(n345), .Z(n351) );
  XOR2_X1 U396 ( .A(n347), .B(n351), .Z(n570) );
  NAND2_X1 U397 ( .A1(n498), .A2(n570), .ZN(n349) );
  XOR2_X1 U398 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U400 ( .A(KEYINPUT114), .B(n350), .ZN(n385) );
  INV_X1 U401 ( .A(n351), .ZN(n365) );
  XOR2_X1 U402 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n353) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(G106GAT), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U405 ( .A(n354), .B(KEYINPUT77), .Z(n356) );
  XOR2_X1 U406 ( .A(G190GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U407 ( .A(n436), .B(G162GAT), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n358) );
  NAND2_X1 U410 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U412 ( .A(n360), .B(n359), .Z(n363) );
  XNOR2_X1 U413 ( .A(n361), .B(KEYINPUT78), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U415 ( .A(n365), .B(n364), .Z(n556) );
  XOR2_X1 U416 ( .A(G78GAT), .B(G155GAT), .Z(n367) );
  XNOR2_X1 U417 ( .A(G183GAT), .B(G71GAT), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U419 ( .A(KEYINPUT79), .B(G64GAT), .Z(n369) );
  XNOR2_X1 U420 ( .A(G8GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U422 ( .A(n371), .B(n370), .ZN(n383) );
  XOR2_X1 U423 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n373) );
  XNOR2_X1 U424 ( .A(KEYINPUT80), .B(KEYINPUT15), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n379) );
  XOR2_X1 U426 ( .A(n374), .B(G211GAT), .Z(n377) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(n375), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U429 ( .A(n379), .B(n378), .Z(n381) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U431 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U432 ( .A(n383), .B(n382), .Z(n578) );
  NOR2_X1 U433 ( .A1(n556), .A2(n578), .ZN(n384) );
  AND2_X1 U434 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U435 ( .A(n386), .B(KEYINPUT47), .ZN(n392) );
  INV_X1 U436 ( .A(n578), .ZN(n457) );
  XNOR2_X1 U437 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n387) );
  XNOR2_X1 U438 ( .A(n387), .B(n556), .ZN(n583) );
  NOR2_X1 U439 ( .A1(n457), .A2(n583), .ZN(n388) );
  XOR2_X1 U440 ( .A(KEYINPUT45), .B(n388), .Z(n389) );
  NOR2_X1 U441 ( .A1(n575), .A2(n389), .ZN(n390) );
  INV_X1 U442 ( .A(n570), .ZN(n499) );
  XOR2_X1 U443 ( .A(n499), .B(KEYINPUT70), .Z(n559) );
  INV_X1 U444 ( .A(n559), .ZN(n455) );
  NAND2_X1 U445 ( .A1(n390), .A2(n455), .ZN(n391) );
  NAND2_X1 U446 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(KEYINPUT48), .B(n393), .ZN(n547) );
  XOR2_X1 U448 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n395) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U451 ( .A(n397), .B(n396), .Z(n401) );
  XOR2_X1 U452 ( .A(G183GAT), .B(KEYINPUT17), .Z(n399) );
  XNOR2_X1 U453 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n440) );
  XNOR2_X1 U455 ( .A(G36GAT), .B(n440), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n405) );
  XNOR2_X1 U458 ( .A(G190GAT), .B(G92GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U460 ( .A(n407), .B(n406), .Z(n520) );
  INV_X1 U461 ( .A(n520), .ZN(n490) );
  NAND2_X1 U462 ( .A1(n547), .A2(n490), .ZN(n409) );
  XOR2_X1 U463 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n431) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XOR2_X1 U466 ( .A(G148GAT), .B(G120GAT), .Z(n411) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(G141GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U469 ( .A(G134GAT), .B(G85GAT), .Z(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n430) );
  XOR2_X1 U472 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n417) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G57GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U475 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n428) );
  XOR2_X1 U479 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n423) );
  XNOR2_X1 U480 ( .A(KEYINPUT83), .B(G127GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U482 ( .A(G113GAT), .B(n424), .Z(n448) );
  INV_X1 U483 ( .A(n448), .ZN(n426) );
  XOR2_X1 U484 ( .A(n426), .B(n425), .Z(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n517) );
  INV_X1 U487 ( .A(n517), .ZN(n546) );
  NOR2_X2 U488 ( .A1(n431), .A2(n546), .ZN(n569) );
  NAND2_X1 U489 ( .A1(n464), .A2(n569), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n432), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U491 ( .A(G176GAT), .B(KEYINPUT84), .Z(n434) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(KEYINPUT85), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n447) );
  XOR2_X1 U494 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n438) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U497 ( .A(n439), .B(G99GAT), .Z(n445) );
  XOR2_X1 U498 ( .A(n440), .B(G15GAT), .Z(n442) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U504 ( .A(n449), .B(n448), .Z(n522) );
  INV_X1 U505 ( .A(n522), .ZN(n530) );
  NAND2_X1 U506 ( .A1(n566), .A2(n556), .ZN(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n452) );
  OR2_X1 U508 ( .A1(n455), .A2(n575), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n456), .B(KEYINPUT75), .ZN(n486) );
  NOR2_X1 U510 ( .A1(n457), .A2(n556), .ZN(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT81), .B(n458), .Z(n459) );
  XNOR2_X1 U512 ( .A(KEYINPUT16), .B(n459), .ZN(n472) );
  XNOR2_X1 U513 ( .A(n520), .B(KEYINPUT99), .ZN(n460) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(n460), .ZN(n467) );
  XOR2_X1 U515 ( .A(n464), .B(KEYINPUT28), .Z(n496) );
  INV_X1 U516 ( .A(n496), .ZN(n527) );
  NAND2_X1 U517 ( .A1(n467), .A2(n527), .ZN(n531) );
  NOR2_X1 U518 ( .A1(n530), .A2(n531), .ZN(n461) );
  NOR2_X1 U519 ( .A1(n517), .A2(n461), .ZN(n471) );
  NAND2_X1 U520 ( .A1(n530), .A2(n490), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n464), .A2(n462), .ZN(n463) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n463), .Z(n468) );
  XNOR2_X1 U523 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n530), .A2(n464), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n466), .B(n465), .ZN(n568) );
  NAND2_X1 U526 ( .A1(n568), .A2(n467), .ZN(n548) );
  NAND2_X1 U527 ( .A1(n468), .A2(n548), .ZN(n469) );
  NOR2_X1 U528 ( .A1(n546), .A2(n469), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n484) );
  NAND2_X1 U530 ( .A1(n472), .A2(n484), .ZN(n500) );
  INV_X1 U531 ( .A(n500), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n486), .A2(n473), .ZN(n480) );
  NOR2_X1 U533 ( .A1(n517), .A2(n480), .ZN(n475) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n520), .A2(n480), .ZN(n477) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U539 ( .A1(n522), .A2(n480), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n527), .A2(n480), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT102), .B(n481), .Z(n482) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n583), .A2(n578), .ZN(n483) );
  NAND2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n485), .ZN(n516) );
  NAND2_X1 U548 ( .A1(n516), .A2(n486), .ZN(n487) );
  XOR2_X1 U549 ( .A(KEYINPUT38), .B(n487), .Z(n495) );
  NAND2_X1 U550 ( .A1(n546), .A2(n495), .ZN(n489) );
  XOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .Z(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n495), .A2(n490), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  NAND2_X1 U556 ( .A1(n495), .A2(n530), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U559 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  NAND2_X1 U561 ( .A1(n498), .A2(n499), .ZN(n514) );
  NOR2_X1 U562 ( .A1(n514), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(n501), .Z(n510) );
  NOR2_X1 U564 ( .A1(n510), .A2(n517), .ZN(n505) );
  XOR2_X1 U565 ( .A(KEYINPUT105), .B(KEYINPUT107), .Z(n503) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n510), .A2(n520), .ZN(n506) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n506), .Z(n507) );
  XNOR2_X1 U571 ( .A(KEYINPUT108), .B(n507), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n510), .A2(n522), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n510), .A2(n527), .ZN(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  INV_X1 U579 ( .A(n514), .ZN(n515) );
  NAND2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n526) );
  NOR2_X1 U581 ( .A1(n517), .A2(n526), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n526), .ZN(n521) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n525) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(n529), .B(n528), .Z(G1339GAT) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT117), .Z(n536) );
  NAND2_X1 U594 ( .A1(n530), .A2(n546), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n533), .A2(n547), .ZN(n534) );
  XOR2_X1 U597 ( .A(KEYINPUT116), .B(n534), .Z(n543) );
  NAND2_X1 U598 ( .A1(n543), .A2(n559), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n538) );
  NAND2_X1 U601 ( .A1(n498), .A2(n543), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(n539), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n541) );
  NAND2_X1 U605 ( .A1(n543), .A2(n578), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U609 ( .A1(n543), .A2(n556), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n549) );
  NOR2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U613 ( .A(n550), .B(KEYINPUT120), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n557), .A2(n570), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U617 ( .A1(n498), .A2(n557), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n578), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n562) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT123), .B(n563), .Z(n565) );
  NAND2_X1 U630 ( .A1(n498), .A2(n566), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n578), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n582) );
  INV_X1 U635 ( .A(n582), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n579), .A2(n570), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U642 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

