//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT30), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT64), .A2(G134), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(G134), .A2(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n192), .A2(new_n193), .ZN(new_n201));
  OAI211_X1 g015(.A(G131), .B(new_n200), .C1(new_n201), .C2(G137), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n199), .B2(new_n202), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(KEYINPUT1), .A3(G146), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n212), .B(new_n213), .C1(G128), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n204), .A2(new_n205), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(KEYINPUT0), .A3(G128), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G128), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n194), .A2(new_n196), .A3(new_n198), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n222), .B2(new_n199), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n189), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n211), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n206), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n213), .A4(new_n212), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n199), .A3(new_n202), .ZN(new_n231));
  INV_X1    g045(.A(new_n223), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(KEYINPUT30), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n236), .A3(new_n232), .ZN(new_n239));
  INV_X1    g053(.A(G210), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n240), .A2(G237), .A3(G953), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT27), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT26), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n238), .A2(new_n239), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n238), .A2(KEYINPUT67), .A3(new_n239), .A4(new_n245), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n188), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n199), .A2(new_n202), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n225), .B2(new_n229), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n252), .A2(new_n223), .A3(new_n237), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n215), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT30), .B1(new_n256), .B2(new_n232), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n252), .A2(new_n223), .A3(new_n189), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n253), .B1(new_n259), .B2(new_n237), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n188), .A3(new_n245), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n236), .B1(new_n256), .B2(new_n232), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT28), .B1(new_n262), .B2(new_n253), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n239), .A2(KEYINPUT68), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n253), .B2(KEYINPUT28), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n245), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n187), .B1(new_n250), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT69), .B(new_n187), .C1(new_n250), .C2(new_n271), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT32), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G472), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n267), .A2(new_n265), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n237), .B1(new_n252), .B2(new_n223), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n239), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(KEYINPUT28), .ZN(new_n284));
  AOI211_X1 g098(.A(KEYINPUT71), .B(new_n264), .C1(new_n239), .C2(new_n282), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n278), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT72), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n238), .A2(new_n239), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n290), .B2(new_n269), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n263), .A2(new_n265), .A3(new_n267), .A4(new_n245), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n257), .A2(new_n258), .A3(new_n236), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n269), .B1(new_n294), .B2(new_n253), .ZN(new_n295));
  AND4_X1   g109(.A1(new_n289), .A2(new_n295), .A3(new_n279), .A4(new_n292), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n288), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n286), .A2(KEYINPUT72), .A3(new_n287), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n277), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT32), .B(new_n187), .C1(new_n250), .C2(new_n271), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n276), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G125), .B(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n210), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(KEYINPUT75), .ZN(new_n305));
  INV_X1    g119(.A(G125), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n306), .A2(KEYINPUT16), .A3(G140), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(new_n303), .B2(KEYINPUT16), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G146), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n206), .A2(G119), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT23), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n206), .A2(G119), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G110), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT74), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n314), .A2(new_n312), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT24), .B(G110), .Z(new_n320));
  OR2_X1    g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n311), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n308), .B(new_n210), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(new_n319), .B2(new_n320), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n316), .B2(new_n315), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G953), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(G221), .A3(G234), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT22), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(G137), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n331), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n322), .B2(new_n326), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT25), .B1(new_n335), .B2(G902), .ZN(new_n336));
  NAND2_X1  g150(.A1(G217), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(G217), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT73), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n332), .A2(new_n341), .A3(new_n287), .A4(new_n334), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n340), .A2(G902), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT76), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n332), .A2(new_n345), .A3(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT77), .B1(new_n302), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n220), .A2(G125), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(G125), .B2(new_n215), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n328), .A2(G224), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n353));
  XOR2_X1   g167(.A(G110), .B(G122), .Z(new_n354));
  INV_X1    g168(.A(G104), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G107), .ZN(new_n356));
  INV_X1    g170(.A(G107), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n357), .A2(KEYINPUT3), .A3(G104), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT3), .B1(new_n357), .B2(G104), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G101), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n244), .B(new_n356), .C1(new_n358), .C2(new_n359), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n355), .B2(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(KEYINPUT3), .A3(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n244), .B1(new_n367), .B2(new_n356), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT79), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n365), .A2(new_n366), .B1(new_n355), .B2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n372));
  NOR4_X1   g186(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT4), .A4(new_n244), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n237), .B(new_n363), .C1(new_n370), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n357), .B2(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n357), .A2(G104), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n355), .A2(KEYINPUT80), .A3(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT81), .B1(new_n379), .B2(G101), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(G101), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n362), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n382), .B2(KEYINPUT81), .ZN(new_n383));
  INV_X1    g197(.A(new_n234), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n235), .ZN(new_n385));
  INV_X1    g199(.A(G116), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n386), .A2(KEYINPUT5), .A3(G119), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n234), .B2(KEYINPUT5), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n385), .B1(G113), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n374), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n391), .B1(new_n374), .B2(new_n390), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n354), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n374), .A2(new_n390), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n395), .A2(new_n354), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n353), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(KEYINPUT86), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n374), .A2(new_n390), .A3(new_n391), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n400), .B2(new_n354), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n352), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n351), .A2(KEYINPUT7), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n350), .B(new_n403), .Z(new_n404));
  XOR2_X1   g218(.A(new_n383), .B(new_n389), .Z(new_n405));
  XNOR2_X1  g219(.A(new_n354), .B(KEYINPUT8), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n404), .B(new_n396), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n287), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n402), .A2(new_n287), .A3(new_n409), .A4(new_n407), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G214), .B1(G237), .B2(G902), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT9), .B(G234), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G221), .B1(new_n417), .B2(G902), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n328), .A2(G227), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT78), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n316), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n421), .B(G140), .Z(new_n422));
  INV_X1    g236(.A(KEYINPUT10), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n225), .B2(new_n229), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n424), .A2(new_n425), .A3(new_n383), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n424), .B2(new_n383), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n222), .A2(new_n199), .ZN(new_n429));
  INV_X1    g243(.A(new_n220), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n363), .B(new_n430), .C1(new_n370), .C2(new_n373), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n381), .B2(new_n362), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n433), .A2(new_n216), .A3(new_n380), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n434), .B2(KEYINPUT10), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n429), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n383), .A2(new_n230), .A3(KEYINPUT10), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n424), .A2(new_n425), .A3(new_n383), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n435), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n422), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n422), .B1(new_n447), .B2(new_n437), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT12), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n383), .A2(new_n215), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n216), .B1(new_n433), .B2(new_n380), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n449), .B(new_n437), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n451), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT12), .B1(new_n453), .B2(new_n429), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n448), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT84), .B(new_n422), .C1(new_n436), .C2(new_n443), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n446), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n457), .A2(new_n458), .A3(new_n287), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n450), .A2(new_n423), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n431), .C1(new_n426), .C2(new_n427), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n429), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n462), .A2(new_n429), .B1(new_n454), .B2(new_n452), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n448), .A2(new_n463), .B1(new_n464), .B2(new_n422), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n460), .B(G469), .C1(new_n465), .C2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n422), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n447), .A2(new_n437), .ZN(new_n468));
  INV_X1    g282(.A(new_n422), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n470), .A3(G469), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n458), .A2(new_n287), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(KEYINPUT83), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n418), .B1(new_n459), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(KEYINPUT85), .B(new_n418), .C1(new_n459), .C2(new_n475), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n415), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n274), .A2(new_n275), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT32), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n297), .A2(new_n298), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G472), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n485), .A3(new_n300), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n487));
  INV_X1    g301(.A(new_n347), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n490));
  INV_X1    g304(.A(G237), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n328), .A3(G214), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n208), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G131), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(G143), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n195), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n490), .B1(new_n497), .B2(KEYINPUT17), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n493), .A2(KEYINPUT17), .A3(G131), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT87), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n498), .A2(new_n499), .A3(new_n501), .A4(new_n323), .ZN(new_n502));
  XNOR2_X1  g316(.A(G113), .B(G122), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n355), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT18), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n495), .B1(new_n505), .B2(new_n195), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n303), .A2(new_n210), .ZN(new_n507));
  OAI221_X1 g321(.A(new_n506), .B1(new_n494), .B2(new_n505), .C1(new_n305), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n502), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n303), .B(KEYINPUT19), .Z(new_n510));
  OAI21_X1  g324(.A(new_n497), .B1(G146), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n508), .B1(new_n310), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n504), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n287), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT20), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n509), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n504), .B1(new_n502), .B2(new_n508), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n287), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G475), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n515), .A2(KEYINPUT20), .A3(new_n516), .A4(new_n287), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G122), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT88), .B1(new_n526), .B2(G116), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT88), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n386), .A3(G122), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n527), .A2(new_n529), .B1(G116), .B2(new_n526), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n357), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n192), .A2(new_n193), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n208), .A2(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n206), .A2(G143), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n533), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n206), .A2(G143), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n534), .B1(new_n539), .B2(KEYINPUT13), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(KEYINPUT13), .ZN(new_n543));
  OAI211_X1 g357(.A(KEYINPUT89), .B(new_n534), .C1(new_n539), .C2(KEYINPUT13), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G134), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n531), .B(new_n538), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n526), .A2(G116), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n357), .B1(new_n548), .B2(KEYINPUT14), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n530), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n538), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n536), .A2(new_n537), .A3(new_n532), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n416), .A2(G217), .A3(new_n328), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n547), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n287), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  NOR2_X1   g375(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n565), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n287), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(G234), .A2(G237), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(G952), .A3(new_n328), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT92), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT21), .B(G898), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT93), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(G902), .A3(G953), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n525), .A2(new_n569), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n348), .A2(new_n480), .A3(new_n489), .A4(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G101), .ZN(G3));
  OAI21_X1  g394(.A(new_n287), .B1(new_n250), .B2(new_n271), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n481), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n478), .B2(new_n479), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n415), .A2(new_n577), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n584), .A2(new_n488), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n555), .B2(KEYINPUT94), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n558), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n557), .B1(new_n547), .B2(new_n553), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n556), .A2(new_n558), .A3(new_n589), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n561), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n561), .A2(new_n287), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n561), .B(new_n287), .C1(new_n591), .C2(new_n592), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n587), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n598), .ZN(new_n600));
  NOR4_X1   g414(.A1(new_n595), .A2(new_n600), .A3(KEYINPUT95), .A4(new_n596), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT96), .A3(new_n525), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT96), .B1(new_n602), .B2(new_n525), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n586), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  AOI21_X1  g423(.A(new_n525), .B1(new_n566), .B2(new_n568), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n586), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT97), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT35), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n357), .ZN(G9));
  INV_X1    g428(.A(new_n583), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n333), .A2(KEYINPUT36), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n327), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n327), .A2(new_n616), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n345), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n617), .A2(KEYINPUT98), .A3(new_n345), .A4(new_n618), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n343), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n480), .A2(new_n578), .A3(new_n615), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT37), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n316), .ZN(G12));
  INV_X1    g440(.A(new_n623), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n478), .B2(new_n479), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n276), .A2(new_n301), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n415), .B1(new_n629), .B2(new_n485), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n572), .B1(G900), .B2(new_n575), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n610), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  OR2_X1    g449(.A1(new_n413), .A2(KEYINPUT99), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n413), .A2(KEYINPUT99), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n636), .A2(KEYINPUT38), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n525), .A2(new_n569), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n627), .A2(new_n414), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT67), .B1(new_n260), .B2(new_n245), .ZN(new_n647));
  INV_X1    g461(.A(new_n249), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n269), .B2(new_n283), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n650), .B2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n629), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(KEYINPUT100), .B2(new_n644), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT101), .B1(new_n646), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n478), .A2(new_n479), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n632), .B(KEYINPUT39), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n653), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n661), .A3(new_n642), .A4(new_n645), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n654), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  OAI211_X1 g478(.A(new_n525), .B(new_n632), .C1(new_n599), .C2(new_n601), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n631), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G146), .ZN(G48));
  AOI21_X1  g482(.A(new_n347), .B1(new_n629), .B2(new_n485), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n457), .A2(new_n287), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n457), .A2(new_n458), .A3(new_n287), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n418), .A3(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n673), .A2(new_n415), .A3(new_n577), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n669), .A2(new_n606), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND4_X1  g491(.A1(new_n674), .A2(new_n486), .A3(new_n488), .A4(new_n610), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT103), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n669), .A2(new_n680), .A3(new_n610), .A4(new_n674), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  OAI21_X1  g497(.A(KEYINPUT104), .B1(new_n673), .B2(new_n415), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n458), .B1(new_n457), .B2(new_n287), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n459), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n687));
  INV_X1    g501(.A(new_n414), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n411), .B2(new_n412), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n687), .A3(new_n418), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n578), .A3(new_n486), .A4(new_n623), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NOR2_X1   g507(.A1(new_n284), .A2(new_n285), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n267), .A2(new_n265), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n269), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n261), .B(new_n696), .C1(new_n649), .C2(new_n188), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n187), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n582), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n347), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n643), .B(KEYINPUT105), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n674), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  NAND4_X1  g517(.A1(new_n666), .A2(new_n623), .A3(new_n582), .A4(new_n698), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n691), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT106), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n691), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  AND2_X1   g525(.A1(new_n411), .A2(new_n412), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n465), .A2(KEYINPUT107), .A3(G469), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n471), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n672), .A2(new_n716), .A3(new_n473), .ZN(new_n717));
  INV_X1    g531(.A(new_n418), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n688), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n712), .A2(new_n666), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n272), .A2(new_n482), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n300), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n721), .A2(KEYINPUT109), .A3(new_n300), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n485), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n720), .A2(new_n726), .A3(KEYINPUT42), .A4(new_n488), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT110), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n669), .A2(new_n720), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n669), .A2(new_n732), .A3(new_n720), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  AND3_X1   g550(.A1(new_n717), .A2(new_n712), .A3(new_n719), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n486), .A2(new_n737), .A3(new_n488), .A4(new_n633), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n546), .ZN(G36));
  INV_X1    g555(.A(new_n525), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n602), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT43), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n615), .A3(new_n627), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n413), .A2(new_n688), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n745), .B2(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n465), .A2(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n467), .A2(new_n470), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n753), .A3(G469), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n750), .A2(new_n753), .A3(KEYINPUT112), .A4(G469), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n473), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(KEYINPUT46), .A3(new_n473), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n672), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n418), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n746), .A2(new_n749), .A3(new_n656), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  NAND2_X1  g581(.A1(new_n764), .A2(KEYINPUT47), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n486), .A2(new_n488), .A3(new_n748), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n770), .A3(new_n418), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n768), .A2(new_n666), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  NOR2_X1   g587(.A1(new_n642), .A2(new_n347), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n629), .A2(new_n651), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n743), .A2(new_n718), .A3(new_n688), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n686), .B(KEYINPUT49), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n675), .A2(new_n702), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n682), .A3(new_n692), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n569), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n566), .A2(KEYINPUT113), .A3(new_n568), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n525), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n689), .A2(new_n576), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT114), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n488), .A3(new_n584), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n602), .A2(new_n525), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n584), .A2(new_n488), .A3(new_n585), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n579), .A2(new_n624), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n627), .A2(new_n699), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n720), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n525), .B1(new_n783), .B2(new_n782), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n747), .A2(new_n632), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n628), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n486), .B1(new_n795), .B2(KEYINPUT115), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n780), .A2(new_n791), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n628), .B(new_n630), .C1(new_n633), .C2(new_n666), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n701), .A2(new_n689), .A3(new_n632), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n627), .A2(new_n717), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n418), .A3(new_n652), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n710), .A2(KEYINPUT52), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n708), .B1(new_n691), .B2(new_n705), .ZN(new_n806));
  AOI211_X1 g620(.A(KEYINPUT106), .B(new_n704), .C1(new_n684), .C2(new_n690), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n801), .B(new_n804), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n740), .B1(new_n728), .B2(new_n734), .ZN(new_n812));
  XNOR2_X1  g626(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n800), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT117), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n791), .A2(new_n799), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n779), .A2(new_n682), .A3(new_n692), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n812), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n819), .A3(new_n811), .A4(new_n813), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n812), .A2(new_n816), .A3(new_n817), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n808), .B(KEYINPUT52), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n815), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n800), .A2(new_n811), .A3(new_n821), .A4(new_n812), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT54), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n748), .A2(new_n673), .A3(new_n572), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n775), .A2(new_n488), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT120), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n525), .A3(new_n602), .ZN(new_n835));
  INV_X1    g649(.A(new_n744), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(new_n832), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n792), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n686), .A2(new_n418), .A3(new_n688), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n642), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n744), .A2(new_n572), .A3(new_n347), .A4(new_n699), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n768), .A2(new_n771), .ZN(new_n850));
  INV_X1    g664(.A(new_n686), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(new_n418), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n843), .A2(new_n747), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n848), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n846), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n838), .A2(new_n849), .A3(new_n854), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n852), .A2(KEYINPUT121), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n852), .A2(KEYINPUT121), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n853), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n855), .A2(new_n846), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(KEYINPUT51), .A3(new_n864), .A4(new_n838), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n328), .A2(G952), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT122), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n834), .A2(new_n605), .A3(new_n604), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n726), .A2(new_n488), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n837), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT48), .Z(new_n872));
  AOI211_X1 g686(.A(new_n868), .B(new_n872), .C1(new_n691), .C2(new_n843), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n860), .A2(new_n865), .A3(new_n867), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n831), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(G952), .A2(G953), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n778), .B1(new_n875), .B2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n397), .A2(new_n401), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT123), .Z(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT55), .Z(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n352), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n827), .A2(G902), .A3(new_n828), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n240), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n883), .B2(KEYINPUT56), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n328), .A2(G952), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n827), .A2(KEYINPUT124), .A3(G902), .A4(new_n828), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n892), .B2(new_n410), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n887), .A2(new_n893), .ZN(G51));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n756), .A3(new_n757), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n472), .B(KEYINPUT57), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n829), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n457), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n885), .B1(new_n895), .B2(new_n899), .ZN(G54));
  NAND2_X1  g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n515), .B1(new_n892), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n515), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n901), .C1(new_n890), .C2(new_n891), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n905), .A3(new_n885), .ZN(G60));
  XOR2_X1   g720(.A(new_n596), .B(KEYINPUT59), .Z(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n897), .B2(new_n829), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n593), .A2(new_n594), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n886), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n831), .A2(new_n907), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n909), .ZN(G63));
  XOR2_X1   g726(.A(new_n337), .B(KEYINPUT60), .Z(new_n913));
  NAND3_X1  g727(.A1(new_n827), .A2(new_n828), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n617), .A2(new_n618), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n335), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n886), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n916), .A2(KEYINPUT61), .A3(new_n886), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(G66));
  AOI21_X1  g736(.A(new_n328), .B1(new_n574), .B2(G224), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n780), .A2(new_n791), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT125), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n926), .B2(new_n328), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n879), .B1(G898), .B2(new_n328), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT126), .Z(new_n929));
  XNOR2_X1  g743(.A(new_n927), .B(new_n929), .ZN(G69));
  NAND2_X1  g744(.A1(new_n701), .A2(new_n689), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n765), .A2(new_n656), .A3(new_n870), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n812), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n766), .A2(new_n772), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n710), .A2(new_n801), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n937), .A3(new_n328), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n259), .B(new_n510), .Z(new_n939));
  NAND2_X1  g753(.A1(G900), .A2(G953), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n942));
  INV_X1    g756(.A(new_n663), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n936), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n663), .A2(KEYINPUT62), .A3(new_n710), .A4(new_n801), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n657), .A2(new_n748), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n789), .A2(new_n785), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n947), .A2(new_n348), .A3(new_n489), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(G953), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n941), .B(KEYINPUT127), .C1(new_n950), .C2(new_n939), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n328), .B1(G227), .B2(G900), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G72));
  NAND3_X1  g767(.A1(new_n925), .A2(new_n937), .A3(new_n934), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  AOI21_X1  g770(.A(new_n290), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n885), .B1(new_n957), .B2(new_n269), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n946), .A2(new_n925), .A3(new_n949), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n956), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n290), .A3(new_n245), .ZN(new_n961));
  INV_X1    g775(.A(new_n295), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n825), .B(new_n956), .C1(new_n649), .C2(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n958), .A2(new_n961), .A3(new_n963), .ZN(G57));
endmodule


