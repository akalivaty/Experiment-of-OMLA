

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(n659), .ZN(n627) );
  NOR2_X2 U551 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U552 ( .A1(n525), .A2(n524), .ZN(n790) );
  XNOR2_X1 U553 ( .A(n596), .B(KEYINPUT13), .ZN(n515) );
  AND2_X1 U554 ( .A1(n603), .A2(n602), .ZN(n613) );
  INV_X1 U555 ( .A(KEYINPUT94), .ZN(n611) );
  INV_X1 U556 ( .A(KEYINPUT99), .ZN(n736) );
  XNOR2_X1 U557 ( .A(n737), .B(n736), .ZN(n750) );
  NOR2_X1 U558 ( .A1(G651), .A2(n525), .ZN(n794) );
  NOR2_X1 U559 ( .A1(n600), .A2(n599), .ZN(n961) );
  NOR2_X1 U560 ( .A1(n549), .A2(n548), .ZN(G160) );
  INV_X1 U561 ( .A(G651), .ZN(n524) );
  NOR2_X1 U562 ( .A1(G543), .A2(n524), .ZN(n516) );
  XOR2_X1 U563 ( .A(KEYINPUT1), .B(n516), .Z(n797) );
  XNOR2_X1 U564 ( .A(G543), .B(KEYINPUT0), .ZN(n517) );
  XNOR2_X1 U565 ( .A(n517), .B(KEYINPUT65), .ZN(n525) );
  NAND2_X1 U566 ( .A1(G49), .A2(n794), .ZN(n519) );
  NAND2_X1 U567 ( .A1(G87), .A2(n525), .ZN(n518) );
  NAND2_X1 U568 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U569 ( .A1(n797), .A2(n520), .ZN(n522) );
  NAND2_X1 U570 ( .A1(G651), .A2(G74), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(G288) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n789) );
  NAND2_X1 U573 ( .A1(n789), .A2(G88), .ZN(n523) );
  XNOR2_X1 U574 ( .A(n523), .B(KEYINPUT78), .ZN(n527) );
  NAND2_X1 U575 ( .A1(G75), .A2(n790), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U577 ( .A(KEYINPUT79), .B(n528), .ZN(n532) );
  NAND2_X1 U578 ( .A1(G50), .A2(n794), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G62), .A2(n797), .ZN(n529) );
  AND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(G303) );
  INV_X1 U582 ( .A(G2104), .ZN(n536) );
  AND2_X1 U583 ( .A1(n536), .A2(G2105), .ZN(n988) );
  NAND2_X1 U584 ( .A1(G126), .A2(n988), .ZN(n534) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n989) );
  NAND2_X1 U586 ( .A1(G114), .A2(n989), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U588 ( .A(KEYINPUT84), .B(n535), .ZN(n542) );
  NOR2_X4 U589 ( .A1(G2105), .A2(n536), .ZN(n992) );
  NAND2_X1 U590 ( .A1(G102), .A2(n992), .ZN(n540) );
  NOR2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XOR2_X1 U592 ( .A(n537), .B(KEYINPUT17), .Z(n538) );
  XNOR2_X1 U593 ( .A(KEYINPUT64), .B(n538), .ZN(n878) );
  NAND2_X1 U594 ( .A1(G138), .A2(n878), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U596 ( .A1(n542), .A2(n541), .ZN(G164) );
  NAND2_X1 U597 ( .A1(G137), .A2(n878), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G125), .A2(n988), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n549) );
  NAND2_X1 U600 ( .A1(n989), .A2(G113), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G101), .A2(n992), .ZN(n545) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(n545), .Z(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G52), .A2(n794), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G64), .A2(n797), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G90), .A2(n789), .ZN(n553) );
  NAND2_X1 U608 ( .A1(G77), .A2(n790), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U612 ( .A(KEYINPUT66), .B(n557), .ZN(G171) );
  NAND2_X1 U613 ( .A1(n789), .A2(G89), .ZN(n558) );
  XNOR2_X1 U614 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G76), .A2(n790), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n561), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U618 ( .A1(n797), .A2(G63), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT70), .ZN(n564) );
  NAND2_X1 U620 ( .A1(G51), .A2(n794), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U622 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U624 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U625 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U626 ( .A1(G86), .A2(n789), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G61), .A2(n797), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n790), .A2(G73), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT2), .B(n571), .Z(n572) );
  NOR2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U632 ( .A(KEYINPUT77), .B(n574), .Z(n576) );
  NAND2_X1 U633 ( .A1(n794), .A2(G48), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(G305) );
  AND2_X1 U635 ( .A1(n794), .A2(G47), .ZN(n580) );
  NAND2_X1 U636 ( .A1(G85), .A2(n789), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G72), .A2(n790), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U639 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n797), .A2(G60), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n582), .A2(n581), .ZN(G290) );
  NOR2_X1 U642 ( .A1(G1976), .A2(G288), .ZN(n681) );
  NOR2_X1 U643 ( .A1(G1971), .A2(G303), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n681), .A2(n583), .ZN(n906) );
  NOR2_X1 U645 ( .A1(G164), .A2(G1384), .ZN(n704) );
  NAND2_X1 U646 ( .A1(G160), .A2(G40), .ZN(n703) );
  INV_X1 U647 ( .A(n703), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n704), .A2(n584), .ZN(n659) );
  NOR2_X1 U649 ( .A1(G2084), .A2(n659), .ZN(n646) );
  NAND2_X1 U650 ( .A1(G8), .A2(n646), .ZN(n657) );
  NAND2_X1 U651 ( .A1(G8), .A2(n659), .ZN(n729) );
  NOR2_X1 U652 ( .A1(G1966), .A2(n729), .ZN(n655) );
  NAND2_X1 U653 ( .A1(G1996), .A2(n627), .ZN(n585) );
  XNOR2_X1 U654 ( .A(KEYINPUT26), .B(n585), .ZN(n589) );
  INV_X1 U655 ( .A(KEYINPUT26), .ZN(n587) );
  INV_X1 U656 ( .A(G1341), .ZN(n586) );
  NOR2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n659), .A2(n588), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n589), .A2(n591), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n590), .A2(KEYINPUT92), .ZN(n603) );
  INV_X1 U661 ( .A(n591), .ZN(n592) );
  OR2_X1 U662 ( .A1(KEYINPUT92), .A2(n592), .ZN(n601) );
  NAND2_X1 U663 ( .A1(n789), .A2(G81), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n593), .B(KEYINPUT12), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G68), .A2(n790), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G43), .A2(n794), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n515), .A2(n597), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n797), .A2(G56), .ZN(n598) );
  XOR2_X1 U670 ( .A(KEYINPUT14), .B(n598), .Z(n599) );
  AND2_X1 U671 ( .A1(n601), .A2(n961), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G92), .A2(n789), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G79), .A2(n790), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G54), .A2(n794), .ZN(n607) );
  NAND2_X1 U676 ( .A1(G66), .A2(n797), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U679 ( .A(KEYINPUT15), .B(n610), .Z(n962) );
  NOR2_X1 U680 ( .A1(n613), .A2(n962), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(n611), .ZN(n620) );
  NAND2_X1 U682 ( .A1(n613), .A2(n962), .ZN(n618) );
  AND2_X1 U683 ( .A1(n659), .A2(G1348), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n614), .B(KEYINPUT93), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n627), .A2(G2067), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n620), .A2(n619), .ZN(n634) );
  NAND2_X1 U689 ( .A1(G53), .A2(n794), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G65), .A2(n797), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U692 ( .A1(G91), .A2(n789), .ZN(n624) );
  NAND2_X1 U693 ( .A1(G78), .A2(n790), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U695 ( .A1(n626), .A2(n625), .ZN(n1025) );
  INV_X1 U696 ( .A(KEYINPUT91), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G2072), .A2(n627), .ZN(n628) );
  XNOR2_X1 U698 ( .A(KEYINPUT27), .B(n628), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n632) );
  AND2_X1 U700 ( .A1(n659), .A2(G1956), .ZN(n631) );
  NOR2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n1025), .A2(n635), .ZN(n633) );
  NAND2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n638) );
  NOR2_X1 U704 ( .A1(n1025), .A2(n635), .ZN(n636) );
  XOR2_X1 U705 ( .A(n636), .B(KEYINPUT28), .Z(n637) );
  NAND2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n639), .B(KEYINPUT29), .ZN(n643) );
  XNOR2_X1 U708 ( .A(G2078), .B(KEYINPUT25), .ZN(n854) );
  NOR2_X1 U709 ( .A1(n659), .A2(n854), .ZN(n641) );
  INV_X1 U710 ( .A(G1961), .ZN(n934) );
  NOR2_X1 U711 ( .A1(n627), .A2(n934), .ZN(n640) );
  NOR2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n645) );
  AND2_X1 U713 ( .A1(n645), .A2(G171), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n644), .B(KEYINPUT95), .ZN(n667) );
  NOR2_X1 U715 ( .A1(n645), .A2(G171), .ZN(n652) );
  NOR2_X1 U716 ( .A1(n655), .A2(n646), .ZN(n647) );
  XNOR2_X1 U717 ( .A(KEYINPUT96), .B(n647), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n648), .A2(G8), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT30), .B(n649), .ZN(n650) );
  NOR2_X1 U720 ( .A1(G168), .A2(n650), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U722 ( .A(KEYINPUT31), .B(n653), .Z(n665) );
  AND2_X1 U723 ( .A1(n667), .A2(n665), .ZN(n654) );
  NOR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n674) );
  INV_X1 U726 ( .A(G8), .ZN(n664) );
  NOR2_X1 U727 ( .A1(G1971), .A2(n729), .ZN(n658) );
  XOR2_X1 U728 ( .A(KEYINPUT97), .B(n658), .Z(n661) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n659), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n662), .A2(G303), .ZN(n663) );
  OR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U733 ( .A1(n665), .A2(n668), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n671) );
  INV_X1 U735 ( .A(n668), .ZN(n669) );
  OR2_X1 U736 ( .A1(n669), .A2(G286), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(KEYINPUT32), .B(n672), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n725) );
  NAND2_X1 U740 ( .A1(n906), .A2(n725), .ZN(n676) );
  INV_X1 U741 ( .A(KEYINPUT98), .ZN(n675) );
  XNOR2_X1 U742 ( .A(n676), .B(n675), .ZN(n679) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n905) );
  INV_X1 U744 ( .A(n729), .ZN(n677) );
  NAND2_X1 U745 ( .A1(n905), .A2(n677), .ZN(n678) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n680), .A2(KEYINPUT33), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n681), .A2(KEYINPUT33), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n682), .A2(n729), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n722) );
  XOR2_X1 U751 ( .A(G1981), .B(G305), .Z(n919) );
  NAND2_X1 U752 ( .A1(G119), .A2(n988), .ZN(n686) );
  NAND2_X1 U753 ( .A1(G107), .A2(n989), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n992), .A2(G95), .ZN(n687) );
  XOR2_X1 U756 ( .A(KEYINPUT88), .B(n687), .Z(n688) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n691) );
  BUF_X1 U758 ( .A(n878), .Z(n993) );
  NAND2_X1 U759 ( .A1(G131), .A2(n993), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n1000) );
  AND2_X1 U761 ( .A1(n1000), .A2(G1991), .ZN(n702) );
  XOR2_X1 U762 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n693) );
  NAND2_X1 U763 ( .A1(G105), .A2(n992), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n693), .B(n692), .ZN(n698) );
  NAND2_X1 U765 ( .A1(G129), .A2(n988), .ZN(n695) );
  NAND2_X1 U766 ( .A1(G117), .A2(n989), .ZN(n694) );
  NAND2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U768 ( .A(KEYINPUT89), .B(n696), .Z(n697) );
  NOR2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U770 ( .A1(G141), .A2(n993), .ZN(n699) );
  NAND2_X1 U771 ( .A1(n700), .A2(n699), .ZN(n1010) );
  AND2_X1 U772 ( .A1(n1010), .A2(G1996), .ZN(n701) );
  NOR2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n866) );
  NOR2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n747) );
  INV_X1 U775 ( .A(n747), .ZN(n705) );
  NOR2_X1 U776 ( .A1(n866), .A2(n705), .ZN(n740) );
  NAND2_X1 U777 ( .A1(G104), .A2(n992), .ZN(n707) );
  NAND2_X1 U778 ( .A1(G140), .A2(n993), .ZN(n706) );
  NAND2_X1 U779 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U780 ( .A(KEYINPUT34), .B(n708), .ZN(n714) );
  NAND2_X1 U781 ( .A1(n989), .A2(G116), .ZN(n709) );
  XNOR2_X1 U782 ( .A(n709), .B(KEYINPUT86), .ZN(n711) );
  NAND2_X1 U783 ( .A1(G128), .A2(n988), .ZN(n710) );
  NAND2_X1 U784 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U785 ( .A(KEYINPUT35), .B(n712), .Z(n713) );
  NOR2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U787 ( .A(KEYINPUT36), .B(n715), .ZN(n1013) );
  XOR2_X1 U788 ( .A(G2067), .B(KEYINPUT37), .Z(n716) );
  XNOR2_X1 U789 ( .A(KEYINPUT85), .B(n716), .ZN(n745) );
  NOR2_X1 U790 ( .A1(n1013), .A2(n745), .ZN(n869) );
  NAND2_X1 U791 ( .A1(n869), .A2(n747), .ZN(n717) );
  XOR2_X1 U792 ( .A(KEYINPUT87), .B(n717), .Z(n743) );
  XNOR2_X1 U793 ( .A(G1986), .B(G290), .ZN(n913) );
  NAND2_X1 U794 ( .A1(n747), .A2(n913), .ZN(n718) );
  NAND2_X1 U795 ( .A1(n743), .A2(n718), .ZN(n719) );
  OR2_X1 U796 ( .A1(n740), .A2(n719), .ZN(n733) );
  INV_X1 U797 ( .A(n733), .ZN(n720) );
  AND2_X1 U798 ( .A1(n919), .A2(n720), .ZN(n721) );
  NAND2_X1 U799 ( .A1(n722), .A2(n721), .ZN(n735) );
  NOR2_X1 U800 ( .A1(G2090), .A2(G303), .ZN(n723) );
  NAND2_X1 U801 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n726) );
  AND2_X1 U803 ( .A1(n726), .A2(n729), .ZN(n731) );
  NOR2_X1 U804 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XOR2_X1 U805 ( .A(n727), .B(KEYINPUT24), .Z(n728) );
  NOR2_X1 U806 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n732) );
  OR2_X1 U808 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n737) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n1010), .ZN(n893) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n738) );
  NOR2_X1 U812 ( .A1(G1991), .A2(n1000), .ZN(n870) );
  NOR2_X1 U813 ( .A1(n738), .A2(n870), .ZN(n739) );
  NOR2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U815 ( .A1(n893), .A2(n741), .ZN(n742) );
  XNOR2_X1 U816 ( .A(KEYINPUT39), .B(n742), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n1013), .A2(n745), .ZN(n890) );
  NAND2_X1 U819 ( .A1(n746), .A2(n890), .ZN(n748) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U822 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U823 ( .A(G2427), .B(G2446), .Z(n753) );
  XNOR2_X1 U824 ( .A(G1341), .B(G2430), .ZN(n752) );
  XNOR2_X1 U825 ( .A(n753), .B(n752), .ZN(n754) );
  XOR2_X1 U826 ( .A(n754), .B(G2435), .Z(n756) );
  XNOR2_X1 U827 ( .A(G1348), .B(G2438), .ZN(n755) );
  XNOR2_X1 U828 ( .A(n756), .B(n755), .ZN(n760) );
  XOR2_X1 U829 ( .A(G2454), .B(G2451), .Z(n758) );
  XNOR2_X1 U830 ( .A(KEYINPUT100), .B(G2443), .ZN(n757) );
  XNOR2_X1 U831 ( .A(n758), .B(n757), .ZN(n759) );
  XOR2_X1 U832 ( .A(n760), .B(n759), .Z(n761) );
  AND2_X1 U833 ( .A1(G14), .A2(n761), .ZN(G401) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U835 ( .A(G57), .ZN(G237) );
  INV_X1 U836 ( .A(G132), .ZN(G219) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n762) );
  XNOR2_X1 U839 ( .A(n762), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n830) );
  NAND2_X1 U841 ( .A1(n830), .A2(G567), .ZN(n763) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n763), .Z(G234) );
  NAND2_X1 U843 ( .A1(G860), .A2(n961), .ZN(n764) );
  XOR2_X1 U844 ( .A(KEYINPUT67), .B(n764), .Z(G153) );
  XOR2_X1 U845 ( .A(G171), .B(KEYINPUT68), .Z(G301) );
  NOR2_X1 U846 ( .A1(n962), .A2(G868), .ZN(n765) );
  XNOR2_X1 U847 ( .A(n765), .B(KEYINPUT69), .ZN(n767) );
  NAND2_X1 U848 ( .A1(G868), .A2(G301), .ZN(n766) );
  NAND2_X1 U849 ( .A1(n767), .A2(n766), .ZN(G284) );
  INV_X1 U850 ( .A(G868), .ZN(n812) );
  NAND2_X1 U851 ( .A1(n1025), .A2(n812), .ZN(n768) );
  XNOR2_X1 U852 ( .A(n768), .B(KEYINPUT71), .ZN(n770) );
  NOR2_X1 U853 ( .A1(n812), .A2(G286), .ZN(n769) );
  NOR2_X1 U854 ( .A1(n770), .A2(n769), .ZN(G297) );
  INV_X1 U855 ( .A(G860), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n771), .A2(G559), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n772), .A2(n962), .ZN(n773) );
  XNOR2_X1 U858 ( .A(n773), .B(KEYINPUT16), .ZN(n774) );
  XNOR2_X1 U859 ( .A(KEYINPUT72), .B(n774), .ZN(G148) );
  NAND2_X1 U860 ( .A1(n962), .A2(G868), .ZN(n775) );
  NOR2_X1 U861 ( .A1(G559), .A2(n775), .ZN(n777) );
  AND2_X1 U862 ( .A1(n812), .A2(n961), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(G282) );
  NAND2_X1 U864 ( .A1(G123), .A2(n988), .ZN(n778) );
  XNOR2_X1 U865 ( .A(n778), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G99), .A2(n992), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT73), .B(n779), .Z(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G111), .A2(n989), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G135), .A2(n993), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n1005) );
  XNOR2_X1 U873 ( .A(n1005), .B(G2096), .ZN(n787) );
  INV_X1 U874 ( .A(G2100), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(G156) );
  NAND2_X1 U876 ( .A1(G559), .A2(n962), .ZN(n788) );
  XOR2_X1 U877 ( .A(n961), .B(n788), .Z(n808) );
  NOR2_X1 U878 ( .A1(G860), .A2(n808), .ZN(n802) );
  NAND2_X1 U879 ( .A1(G93), .A2(n789), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G80), .A2(n790), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(KEYINPUT75), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G55), .A2(n794), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n797), .A2(G67), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT76), .B(n798), .Z(n799) );
  OR2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n813) );
  XOR2_X1 U888 ( .A(n813), .B(KEYINPUT74), .Z(n801) );
  XNOR2_X1 U889 ( .A(n802), .B(n801), .ZN(G145) );
  INV_X1 U890 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U891 ( .A(n1025), .B(G290), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(G288), .ZN(n804) );
  XNOR2_X1 U893 ( .A(KEYINPUT19), .B(n804), .ZN(n806) );
  XOR2_X1 U894 ( .A(G305), .B(n813), .Z(n805) );
  XNOR2_X1 U895 ( .A(n806), .B(n805), .ZN(n807) );
  XNOR2_X1 U896 ( .A(G166), .B(n807), .ZN(n965) );
  XNOR2_X1 U897 ( .A(n965), .B(KEYINPUT80), .ZN(n809) );
  XNOR2_X1 U898 ( .A(n809), .B(n808), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n810), .A2(G868), .ZN(n811) );
  XOR2_X1 U900 ( .A(KEYINPUT81), .B(n811), .Z(n815) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U903 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n817), .ZN(n819) );
  XNOR2_X1 U906 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n818) );
  XNOR2_X1 U907 ( .A(n819), .B(n818), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G2072), .A2(n820), .ZN(G158) );
  XNOR2_X1 U909 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U910 ( .A1(G220), .A2(G219), .ZN(n821) );
  XOR2_X1 U911 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U912 ( .A1(G218), .A2(n822), .ZN(n823) );
  XOR2_X1 U913 ( .A(KEYINPUT83), .B(n823), .Z(n824) );
  NAND2_X1 U914 ( .A1(G96), .A2(n824), .ZN(n959) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n959), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G108), .A2(G120), .ZN(n825) );
  NOR2_X1 U917 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G69), .A2(n826), .ZN(n960) );
  NAND2_X1 U919 ( .A1(G567), .A2(n960), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n987) );
  NAND2_X1 U921 ( .A1(G661), .A2(G483), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n987), .A2(n829), .ZN(n833) );
  NAND2_X1 U923 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U929 ( .A(G120), .B(KEYINPUT101), .ZN(G236) );
  NAND2_X1 U931 ( .A1(n993), .A2(G136), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n834), .B(KEYINPUT106), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n836) );
  NAND2_X1 U934 ( .A1(G124), .A2(n988), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G112), .A2(n989), .ZN(n840) );
  NAND2_X1 U938 ( .A1(G100), .A2(n992), .ZN(n839) );
  NAND2_X1 U939 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U940 ( .A(KEYINPUT107), .B(n841), .Z(n842) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(G162) );
  XOR2_X1 U942 ( .A(G29), .B(KEYINPUT120), .Z(n865) );
  XOR2_X1 U943 ( .A(G2084), .B(G34), .Z(n844) );
  XNOR2_X1 U944 ( .A(KEYINPUT54), .B(n844), .ZN(n861) );
  XNOR2_X1 U945 ( .A(G2090), .B(G35), .ZN(n859) );
  XNOR2_X1 U946 ( .A(KEYINPUT117), .B(G2067), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n845), .B(G26), .ZN(n853) );
  XNOR2_X1 U948 ( .A(G1996), .B(G32), .ZN(n847) );
  XNOR2_X1 U949 ( .A(G1991), .B(G25), .ZN(n846) );
  NOR2_X1 U950 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U951 ( .A1(G28), .A2(n848), .ZN(n851) );
  XNOR2_X1 U952 ( .A(KEYINPUT118), .B(G2072), .ZN(n849) );
  XNOR2_X1 U953 ( .A(G33), .B(n849), .ZN(n850) );
  NOR2_X1 U954 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U955 ( .A1(n853), .A2(n852), .ZN(n856) );
  XOR2_X1 U956 ( .A(G27), .B(n854), .Z(n855) );
  NOR2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U958 ( .A(KEYINPUT53), .B(n857), .ZN(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n862), .B(KEYINPUT55), .ZN(n863) );
  XNOR2_X1 U962 ( .A(KEYINPUT119), .B(n863), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n902) );
  XNOR2_X1 U964 ( .A(G160), .B(G2084), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n872) );
  NOR2_X1 U967 ( .A1(n870), .A2(n1005), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U969 ( .A(KEYINPUT114), .B(n873), .ZN(n889) );
  NAND2_X1 U970 ( .A1(G127), .A2(n988), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G115), .A2(n989), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n877) );
  XOR2_X1 U973 ( .A(KEYINPUT110), .B(KEYINPUT47), .Z(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n883) );
  NAND2_X1 U975 ( .A1(G103), .A2(n992), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U978 ( .A(KEYINPUT109), .B(n881), .Z(n882) );
  NOR2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n1008) );
  XNOR2_X1 U980 ( .A(G2072), .B(n1008), .ZN(n885) );
  XNOR2_X1 U981 ( .A(G164), .B(G2078), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U983 ( .A(n886), .B(KEYINPUT115), .Z(n887) );
  XNOR2_X1 U984 ( .A(KEYINPUT50), .B(n887), .ZN(n888) );
  NOR2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n891) );
  NAND2_X1 U986 ( .A1(n891), .A2(n890), .ZN(n896) );
  XOR2_X1 U987 ( .A(G2090), .B(G162), .Z(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(KEYINPUT51), .B(n894), .ZN(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U991 ( .A(KEYINPUT52), .B(n897), .Z(n898) );
  NOR2_X1 U992 ( .A1(KEYINPUT55), .A2(n898), .ZN(n899) );
  XOR2_X1 U993 ( .A(KEYINPUT116), .B(n899), .Z(n900) );
  NAND2_X1 U994 ( .A1(G29), .A2(n900), .ZN(n901) );
  NAND2_X1 U995 ( .A1(n902), .A2(n901), .ZN(n956) );
  XNOR2_X1 U996 ( .A(G16), .B(KEYINPUT56), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n903), .B(KEYINPUT121), .ZN(n927) );
  XNOR2_X1 U998 ( .A(G171), .B(G1961), .ZN(n916) );
  INV_X1 U999 ( .A(G1971), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G166), .A2(n904), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1002 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(KEYINPUT122), .B(n909), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n1025), .B(G1956), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1007 ( .A(KEYINPUT123), .B(n914), .Z(n915) );
  NAND2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n925) );
  XOR2_X1 U1009 ( .A(n961), .B(G1341), .Z(n918) );
  XOR2_X1 U1010 ( .A(G1348), .B(n962), .Z(n917) );
  NOR2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n923) );
  XNOR2_X1 U1012 ( .A(G1966), .B(G168), .ZN(n920) );
  NAND2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(n921), .B(KEYINPUT57), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1016 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1017 ( .A1(n927), .A2(n926), .ZN(n953) );
  XNOR2_X1 U1018 ( .A(G1986), .B(G24), .ZN(n932) );
  XNOR2_X1 U1019 ( .A(G1971), .B(G22), .ZN(n929) );
  XNOR2_X1 U1020 ( .A(G23), .B(G1976), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(KEYINPUT125), .B(n930), .ZN(n931) );
  NOR2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(KEYINPUT58), .B(n933), .ZN(n936) );
  XNOR2_X1 U1025 ( .A(n934), .B(G5), .ZN(n935) );
  NAND2_X1 U1026 ( .A1(n936), .A2(n935), .ZN(n948) );
  XOR2_X1 U1027 ( .A(G1966), .B(G21), .Z(n946) );
  XOR2_X1 U1028 ( .A(G19), .B(G1341), .Z(n940) );
  XNOR2_X1 U1029 ( .A(G1956), .B(G20), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(G6), .B(G1981), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1033 ( .A(KEYINPUT59), .B(G1348), .Z(n941) );
  XNOR2_X1 U1034 ( .A(G4), .B(n941), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(n944), .B(KEYINPUT60), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1039 ( .A(KEYINPUT61), .B(n949), .Z(n951) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT124), .ZN(n950) );
  NOR2_X1 U1041 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1042 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1043 ( .A(KEYINPUT126), .B(n954), .Z(n955) );
  NOR2_X1 U1044 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1045 ( .A1(n957), .A2(G11), .ZN(n958) );
  XOR2_X1 U1046 ( .A(KEYINPUT62), .B(n958), .Z(G311) );
  XNOR2_X1 U1047 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1048 ( .A(G108), .ZN(G238) );
  INV_X1 U1049 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(G325) );
  INV_X1 U1051 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1052 ( .A(G286), .B(n961), .Z(n964) );
  XOR2_X1 U1053 ( .A(G171), .B(n962), .Z(n963) );
  XNOR2_X1 U1054 ( .A(n964), .B(n963), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(n966), .B(n965), .ZN(n967) );
  NOR2_X1 U1056 ( .A1(G37), .A2(n967), .ZN(G397) );
  XOR2_X1 U1057 ( .A(G2100), .B(G2096), .Z(n969) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G2090), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(n969), .B(n968), .ZN(n973) );
  XOR2_X1 U1060 ( .A(G2678), .B(KEYINPUT42), .Z(n971) );
  XNOR2_X1 U1061 ( .A(G2072), .B(KEYINPUT43), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n971), .B(n970), .ZN(n972) );
  XOR2_X1 U1063 ( .A(n973), .B(n972), .Z(n975) );
  XNOR2_X1 U1064 ( .A(G2078), .B(G2084), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n975), .B(n974), .ZN(G227) );
  XOR2_X1 U1066 ( .A(G2474), .B(KEYINPUT103), .Z(n977) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G1976), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n977), .B(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(n978), .B(G1956), .Z(n980) );
  XNOR2_X1 U1070 ( .A(G1996), .B(G1961), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n980), .B(n979), .ZN(n984) );
  XOR2_X1 U1072 ( .A(KEYINPUT104), .B(KEYINPUT41), .Z(n982) );
  XNOR2_X1 U1073 ( .A(G1986), .B(G1971), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n982), .B(n981), .ZN(n983) );
  XOR2_X1 U1075 ( .A(n984), .B(n983), .Z(n986) );
  XNOR2_X1 U1076 ( .A(G1991), .B(G1981), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n986), .B(n985), .ZN(G229) );
  XOR2_X1 U1078 ( .A(KEYINPUT102), .B(n987), .Z(G319) );
  NAND2_X1 U1079 ( .A1(G130), .A2(n988), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(G118), .A2(n989), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n999) );
  NAND2_X1 U1082 ( .A1(G106), .A2(n992), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(G142), .A2(n993), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1085 ( .A(KEYINPUT45), .B(n996), .Z(n997) );
  XNOR2_X1 U1086 ( .A(KEYINPUT108), .B(n997), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XOR2_X1 U1088 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1002) );
  XOR2_X1 U1089 ( .A(n1000), .B(G162), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(n1002), .B(n1001), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(n1004), .B(n1003), .Z(n1007) );
  XNOR2_X1 U1092 ( .A(G160), .B(n1005), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1007), .B(n1006), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(n1009), .B(n1008), .Z(n1012) );
  XOR2_X1 U1095 ( .A(G164), .B(n1010), .Z(n1011) );
  XNOR2_X1 U1096 ( .A(n1012), .B(n1011), .ZN(n1014) );
  XOR2_X1 U1097 ( .A(n1014), .B(n1013), .Z(n1015) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1015), .ZN(G395) );
  XNOR2_X1 U1099 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n1017) );
  NOR2_X1 U1100 ( .A1(G227), .A2(G229), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NOR2_X1 U1102 ( .A1(G397), .A2(n1018), .ZN(n1022) );
  INV_X1 U1103 ( .A(G319), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(G401), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT111), .B(n1020), .Z(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(G395), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(n1024), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U1109 ( .A(G225), .ZN(G308) );
  INV_X1 U1110 ( .A(G69), .ZN(G235) );
  INV_X1 U1111 ( .A(n1025), .ZN(G299) );
endmodule

