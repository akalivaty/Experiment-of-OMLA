//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n202), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G97), .C2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G77), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G1), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G257), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n218), .B(new_n230), .C1(new_n231), .C2(new_n214), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n224), .ZN(new_n234));
  INV_X1    g0034(.A(new_n201), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  AOI22_X1  g0037(.A1(new_n232), .A2(KEYINPUT0), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n228), .B(new_n238), .C1(KEYINPUT0), .C2(new_n232), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n207), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G250), .B(G257), .Z(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n260), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n261), .A2(new_n264), .B1(new_n265), .B2(new_n217), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n223), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n233), .ZN(new_n276));
  NAND3_X1  g0076(.A1(KEYINPUT66), .A2(G33), .A3(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(new_n269), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G232), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n268), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G169), .ZN(new_n282));
  INV_X1    g0082(.A(G179), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(new_n281), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT79), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT7), .B1(new_n264), .B2(new_n224), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT7), .ZN(new_n287));
  NOR4_X1   g0087(.A1(new_n262), .A2(new_n263), .A3(new_n287), .A4(G20), .ZN(new_n288));
  OAI21_X1  g0088(.A(G68), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G159), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G58), .A2(G68), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n224), .B1(new_n235), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n285), .B1(new_n295), .B2(KEYINPUT80), .ZN(new_n296));
  OR2_X1    g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n224), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n287), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n293), .B1(new_n302), .B2(G68), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT79), .B1(new_n303), .B2(new_n291), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT16), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n233), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT16), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT80), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n303), .B2(new_n291), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n310), .B2(new_n285), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT81), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT68), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n306), .B2(new_n233), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n306), .A2(new_n314), .A3(new_n233), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n223), .A2(G13), .A3(G20), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n224), .A2(G1), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT70), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT8), .B(G58), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n322), .A2(new_n326), .B1(new_n321), .B2(new_n325), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n312), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n313), .B1(new_n312), .B2(new_n327), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n284), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT18), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n281), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G190), .B2(new_n281), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n312), .A2(new_n327), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n312), .A2(KEYINPUT17), .A3(new_n327), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT18), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n284), .C1(new_n328), .C2(new_n329), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n331), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n324), .A2(new_n202), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n322), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n265), .A2(G20), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT69), .ZN(new_n347));
  INV_X1    g0147(.A(G150), .ZN(new_n348));
  INV_X1    g0148(.A(new_n290), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n347), .A2(new_n325), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(G20), .B2(new_n203), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n345), .B1(G50), .B2(new_n320), .C1(new_n351), .C2(new_n318), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n279), .A2(G226), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n297), .A2(new_n298), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G223), .A2(G1698), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT67), .B(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(G222), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n267), .C1(new_n220), .C2(new_n354), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n353), .A2(new_n359), .A3(new_n272), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n360), .A2(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n283), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n352), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(G190), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n360), .A2(new_n332), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n352), .B(KEYINPUT9), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT10), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n363), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n343), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n260), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n377));
  INV_X1    g0177(.A(G97), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n377), .A2(new_n264), .B1(new_n265), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n271), .B1(new_n379), .B2(new_n267), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n279), .A2(G238), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(KEYINPUT74), .A3(KEYINPUT13), .A4(new_n381), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n356), .A2(new_n212), .B1(new_n207), .B2(new_n256), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n354), .B1(G33), .B2(G97), .ZN(new_n384));
  INV_X1    g0184(.A(new_n267), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n381), .B(new_n272), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT13), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G179), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT78), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n380), .A2(KEYINPUT13), .A3(new_n381), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n388), .A2(new_n395), .A3(G169), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(KEYINPUT14), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(KEYINPUT78), .A3(G179), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(KEYINPUT14), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n394), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n290), .A2(G50), .ZN(new_n401));
  INV_X1    g0201(.A(G77), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n401), .B1(new_n224), .B2(G68), .C1(new_n347), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n319), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT11), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT77), .B1(new_n321), .B2(new_n208), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT12), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n403), .A2(new_n319), .A3(new_n406), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n324), .A2(new_n321), .A3(new_n307), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(G68), .B1(new_n410), .B2(new_n409), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n408), .A2(new_n411), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n400), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n391), .A2(G190), .ZN(new_n417));
  INV_X1    g0217(.A(new_n415), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n388), .A2(new_n395), .A3(G200), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT15), .B(G87), .Z(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n346), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n422), .B1(new_n221), .B2(new_n224), .C1(new_n349), .C2(new_n325), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n307), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n221), .A2(new_n321), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n413), .A2(G77), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n271), .B1(new_n279), .B2(G244), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n354), .B1(new_n209), .B2(new_n256), .C1(new_n356), .C2(new_n207), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n267), .C1(G107), .C2(new_n354), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OR3_X1    g0231(.A1(new_n431), .A2(KEYINPUT71), .A3(G179), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT71), .B1(new_n431), .B2(G179), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G169), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n431), .A2(G200), .ZN(new_n438));
  INV_X1    g0238(.A(G190), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n427), .B(new_n438), .C1(new_n439), .C2(new_n431), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n416), .A2(new_n420), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n376), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G283), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n224), .C1(G33), .C2(new_n378), .ZN(new_n445));
  INV_X1    g0245(.A(G116), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G20), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n307), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT20), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT89), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n448), .A2(new_n449), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT89), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n453), .A3(new_n449), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n321), .A2(new_n446), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT82), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n265), .B2(G1), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n223), .A2(KEYINPUT82), .A3(G33), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n307), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(G116), .A4(new_n320), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n354), .B1(new_n214), .B2(new_n256), .C1(new_n356), .C2(new_n231), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT88), .B(G303), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n264), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n267), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(G274), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n471), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n278), .A2(new_n474), .A3(G270), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n468), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n463), .A2(G169), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n476), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n463), .A2(new_n480), .A3(G179), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n463), .A2(KEYINPUT21), .A3(G169), .A4(new_n476), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n213), .A2(G20), .ZN(new_n484));
  XOR2_X1   g0284(.A(new_n484), .B(KEYINPUT23), .Z(new_n485));
  AOI21_X1  g0285(.A(G20), .B1(new_n297), .B2(new_n298), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT90), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT22), .A4(G87), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n346), .A2(G116), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n354), .A2(new_n487), .A3(new_n224), .A4(G87), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT22), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n489), .A2(KEYINPUT24), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(new_n490), .A3(new_n488), .A4(new_n485), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n497), .A3(new_n307), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n223), .A2(G13), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT25), .B1(new_n499), .B2(new_n484), .ZN(new_n500));
  OR3_X1    g0300(.A1(new_n499), .A2(new_n484), .A3(KEYINPUT25), .ZN(new_n501));
  INV_X1    g0301(.A(new_n317), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n320), .B(new_n460), .C1(new_n502), .C2(new_n315), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n500), .B(new_n501), .C1(new_n503), .C2(new_n213), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT91), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n318), .A2(G107), .A3(new_n320), .A4(new_n460), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT91), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n506), .A2(new_n507), .A3(new_n500), .A4(new_n501), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n218), .B1(new_n257), .B2(new_n259), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n231), .A2(new_n256), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n354), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n385), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n278), .A2(new_n474), .A3(G264), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G190), .A3(new_n473), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n356), .A2(new_n218), .B1(new_n231), .B2(new_n256), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n354), .B1(G33), .B2(G294), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n473), .B(new_n515), .C1(new_n520), .C2(new_n385), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n498), .A2(new_n509), .A3(new_n518), .A4(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n455), .A2(new_n462), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n476), .A2(G200), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n468), .A2(G190), .A3(new_n473), .A4(new_n475), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n456), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n470), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n278), .A2(G250), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT86), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n278), .A2(KEYINPUT86), .A3(G250), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n470), .A2(G274), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n265), .A2(new_n446), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n356), .A2(new_n209), .B1(new_n219), .B2(new_n256), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n354), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n538), .B2(new_n385), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n435), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n538), .A2(new_n385), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(new_n283), .A3(new_n535), .A4(new_n533), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n486), .A2(G68), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT87), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g0345(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(G20), .B1(G33), .B2(G97), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT19), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OR3_X1    g0348(.A1(new_n265), .A2(new_n378), .A3(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(G20), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n486), .A2(KEYINPUT87), .A3(G68), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n307), .ZN(new_n553));
  INV_X1    g0353(.A(new_n421), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n321), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n503), .A2(new_n554), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n540), .A2(new_n542), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n523), .A2(new_n527), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n473), .ZN(new_n560));
  NOR4_X1   g0360(.A1(new_n514), .A2(new_n516), .A3(G179), .A4(new_n560), .ZN(new_n561));
  AOI221_X4 g0361(.A(new_n561), .B1(new_n435), .B2(new_n521), .C1(new_n498), .C2(new_n509), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n483), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n503), .A2(new_n378), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n302), .A2(G107), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n290), .A2(G77), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n378), .A2(new_n213), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n565), .B(new_n566), .C1(new_n224), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n564), .B1(new_n573), .B2(new_n307), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n354), .A2(new_n260), .A3(G244), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n354), .A2(G250), .A3(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n354), .A2(new_n260), .A3(KEYINPUT4), .A4(G244), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n444), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n267), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n278), .A2(new_n474), .A3(G257), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n278), .A2(new_n474), .A3(KEYINPUT83), .A4(G257), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n560), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  OAI221_X1 g0387(.A(new_n574), .B1(G97), .B2(new_n320), .C1(new_n587), .C2(new_n332), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n581), .A2(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT84), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n581), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT85), .B1(new_n594), .B2(G190), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n581), .A2(new_n592), .A3(new_n586), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n592), .B1(new_n581), .B2(new_n586), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT85), .B(G190), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n589), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n591), .A2(new_n435), .A3(new_n593), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n574), .B1(G97), .B2(new_n320), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n587), .A2(new_n283), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n534), .A2(new_n539), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n332), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n534), .A2(new_n539), .A3(new_n439), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n553), .B(new_n555), .C1(new_n217), .C2(new_n503), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n563), .A2(new_n600), .A3(new_n604), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n443), .A2(new_n611), .ZN(G372));
  INV_X1    g0412(.A(new_n363), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n312), .A2(new_n327), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n284), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n341), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(KEYINPUT18), .A3(new_n284), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n437), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n400), .A2(new_n415), .B1(new_n619), .B2(new_n420), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(new_n339), .ZN(new_n621));
  INV_X1    g0421(.A(new_n374), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n372), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n613), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(G190), .B1(new_n596), .B2(new_n597), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n588), .B1(new_n627), .B2(new_n598), .ZN(new_n628));
  INV_X1    g0428(.A(new_n604), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n628), .A2(new_n629), .A3(new_n609), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n479), .A2(new_n482), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n498), .A2(new_n509), .B1(new_n435), .B2(new_n521), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G179), .B2(new_n521), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n633), .A3(new_n481), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n634), .A3(new_n523), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n604), .A2(new_n609), .A3(KEYINPUT26), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT26), .B1(new_n604), .B2(new_n609), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n636), .A2(new_n558), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n624), .B1(new_n443), .B2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(G13), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(G20), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n223), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n463), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g0450(.A(new_n483), .B(new_n650), .Z(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(new_n527), .ZN(new_n652));
  XOR2_X1   g0452(.A(KEYINPUT92), .B(G330), .Z(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n649), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n562), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n523), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n498), .B2(new_n509), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n659), .B2(new_n562), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n483), .A2(new_n655), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n656), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n661), .A2(new_n665), .ZN(G399));
  NOR2_X1   g0466(.A1(new_n230), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n546), .A2(new_n446), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT93), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n236), .B2(new_n668), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n639), .A2(new_n655), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT29), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(KEYINPUT95), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT96), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n634), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n631), .A2(new_n633), .A3(KEYINPUT96), .A4(new_n481), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n630), .A2(new_n523), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n638), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .A3(new_n655), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT95), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n649), .B1(new_n635), .B2(new_n638), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(KEYINPUT29), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n677), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  NOR4_X1   g0487(.A1(new_n476), .A2(new_n283), .A3(new_n514), .A4(new_n516), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n594), .A2(new_n605), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(KEYINPUT94), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n605), .A2(G179), .A3(new_n480), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n590), .A3(new_n521), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(KEYINPUT94), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n594), .A2(new_n605), .A3(new_n694), .A4(new_n688), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n649), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT31), .B(new_n697), .C1(new_n611), .C2(new_n649), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n699), .A3(new_n649), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n653), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n687), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n674), .B1(new_n703), .B2(G1), .ZN(G364));
  AOI21_X1  g0504(.A(new_n223), .B1(new_n643), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n667), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G13), .A2(G33), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n652), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n233), .B1(G20), .B2(new_n435), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n224), .A2(new_n439), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n283), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n354), .B1(new_n718), .B2(G322), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n283), .A2(new_n332), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n224), .A2(G190), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G317), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT33), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(KEYINPUT33), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G294), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n224), .B1(new_n729), .B2(G190), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n719), .B(new_n727), .C1(new_n728), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n332), .A2(G179), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n721), .A2(new_n729), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(G283), .A2(new_n734), .B1(new_n736), .B2(G329), .ZN(new_n737));
  INV_X1    g0537(.A(G303), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n715), .A2(new_n732), .ZN(new_n739));
  INV_X1    g0539(.A(G311), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n721), .A2(new_n716), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n737), .B1(new_n738), .B2(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n715), .A2(new_n720), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n731), .B(new_n742), .C1(G326), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n734), .A2(G107), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n746), .B1(new_n202), .B2(new_n743), .C1(new_n217), .C2(new_n739), .ZN(new_n747));
  INV_X1    g0547(.A(G159), .ZN(new_n748));
  OR3_X1    g0548(.A1(new_n735), .A2(KEYINPUT32), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT32), .B1(new_n735), .B2(new_n748), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n749), .B(new_n750), .C1(new_n378), .C2(new_n730), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n354), .B1(new_n717), .B2(new_n206), .C1(new_n208), .C2(new_n722), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n221), .A2(new_n741), .ZN(new_n753));
  NOR4_X1   g0553(.A1(new_n747), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n708), .B(new_n713), .C1(new_n714), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n230), .A2(new_n354), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n237), .B2(new_n469), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(new_n251), .B2(new_n469), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n229), .A2(G355), .A3(new_n354), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n760), .B(new_n761), .C1(G116), .C2(new_n229), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n711), .A2(new_n714), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n652), .A2(new_n653), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n707), .B1(new_n652), .B2(new_n653), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n756), .A2(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(G396));
  OAI211_X1 g0569(.A(new_n437), .B(new_n440), .C1(new_n427), .C2(new_n655), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT99), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n437), .B2(new_n655), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n434), .A2(KEYINPUT99), .A3(new_n436), .A4(new_n649), .ZN(new_n773));
  AND3_X1   g0573(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n685), .B(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(new_n702), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n708), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n354), .B1(new_n739), .B2(new_n202), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n733), .A2(new_n208), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n206), .B2(new_n730), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G143), .A2(new_n718), .B1(new_n723), .B2(G150), .ZN(new_n782));
  INV_X1    g0582(.A(G137), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n782), .B1(new_n783), .B2(new_n743), .C1(new_n748), .C2(new_n741), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT98), .Z(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n785), .B2(KEYINPUT34), .ZN(new_n786));
  INV_X1    g0586(.A(G132), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n786), .B1(KEYINPUT34), .B2(new_n785), .C1(new_n787), .C2(new_n735), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n354), .B1(new_n718), .B2(G294), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n789), .B1(new_n378), .B2(new_n730), .C1(new_n790), .C2(new_n722), .ZN(new_n791));
  INV_X1    g0591(.A(new_n741), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G116), .A2(new_n792), .B1(new_n734), .B2(G87), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n213), .B2(new_n739), .C1(new_n740), .C2(new_n735), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n791), .B(new_n794), .C1(G303), .C2(new_n744), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT97), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n788), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n708), .B1(new_n797), .B2(new_n714), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n714), .A2(new_n709), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n798), .B1(G77), .B2(new_n800), .C1(new_n801), .C2(new_n710), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n777), .A2(new_n802), .ZN(G384));
  NAND2_X1  g0603(.A1(new_n415), .A2(new_n649), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n416), .A2(new_n420), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n420), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n415), .B(new_n649), .C1(new_n400), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n698), .A2(new_n808), .A3(new_n700), .A4(new_n801), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT38), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n305), .A2(new_n319), .A3(new_n311), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n327), .ZN(new_n813));
  INV_X1    g0613(.A(new_n647), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n284), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n816), .A3(new_n335), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT37), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n328), .A2(new_n329), .B1(new_n284), .B2(new_n814), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT37), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n335), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n815), .ZN(new_n823));
  AOI221_X4 g0623(.A(new_n811), .B1(new_n818), .B2(new_n822), .C1(new_n343), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n343), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n818), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT38), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n810), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT40), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n814), .B1(new_n328), .B2(new_n329), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT100), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n339), .A2(new_n831), .B1(new_n616), .B2(new_n617), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n337), .A2(KEYINPUT100), .A3(new_n338), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n830), .A2(new_n335), .A3(new_n615), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(KEYINPUT37), .B1(new_n821), .B2(new_n819), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n811), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n825), .A2(KEYINPUT38), .A3(new_n826), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n829), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n828), .A2(new_n829), .B1(new_n839), .B2(new_n810), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n442), .A2(new_n701), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n653), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n442), .A2(new_n677), .A3(new_n683), .A4(new_n686), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n624), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT101), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n843), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n825), .A2(new_n826), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n811), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(KEYINPUT39), .A3(new_n838), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n339), .A2(new_n831), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n618), .A3(new_n833), .ZN(new_n853));
  INV_X1    g0653(.A(new_n329), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n312), .A2(new_n313), .A3(new_n327), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n647), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n615), .A2(new_n335), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n822), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n851), .B1(new_n824), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n416), .A2(new_n649), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n850), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n616), .A2(new_n617), .A3(new_n647), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n523), .B1(new_n483), .B2(new_n562), .ZN(new_n866));
  NOR4_X1   g0666(.A1(new_n866), .A2(new_n628), .A3(new_n629), .A4(new_n609), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n636), .A2(new_n558), .A3(new_n637), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n655), .B(new_n801), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n437), .B2(new_n649), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(new_n808), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n824), .B2(new_n827), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(new_n865), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n847), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n223), .B2(new_n643), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT35), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n224), .B(new_n233), .C1(new_n572), .C2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n877), .B(G116), .C1(new_n876), .C2(new_n572), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT36), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n220), .A2(new_n292), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n880), .A2(new_n236), .B1(G50), .B2(new_n208), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n642), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n879), .A3(new_n882), .ZN(G367));
  NOR2_X1   g0683(.A1(new_n739), .A2(new_n446), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT46), .ZN(new_n885));
  INV_X1    g0685(.A(new_n730), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(G107), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n718), .A2(new_n465), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n741), .A2(new_n790), .B1(new_n735), .B2(new_n724), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(G97), .B2(new_n734), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n264), .B1(new_n722), .B2(new_n728), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(G311), .B2(new_n744), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n887), .A2(new_n888), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n735), .A2(new_n783), .ZN(new_n894));
  INV_X1    g0694(.A(G143), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n743), .A2(new_n895), .B1(new_n739), .B2(new_n206), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n894), .B(new_n896), .C1(new_n220), .C2(new_n734), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n897), .B1(new_n208), .B2(new_n730), .C1(new_n348), .C2(new_n717), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n722), .A2(new_n748), .B1(new_n741), .B2(new_n202), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT105), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n354), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n893), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT47), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n708), .B1(new_n903), .B2(new_n714), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n763), .B1(new_n229), .B2(new_n554), .C1(new_n758), .C2(new_n247), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n610), .A2(new_n558), .B1(new_n608), .B2(new_n649), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n558), .A2(new_n608), .A3(new_n649), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n904), .B(new_n905), .C1(new_n908), .C2(new_n712), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n628), .A2(new_n629), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n602), .A2(new_n649), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n910), .A2(new_n911), .B1(new_n629), .B2(new_n649), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n665), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT45), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n665), .A2(new_n912), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT44), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n661), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n916), .ZN(new_n918));
  INV_X1    g0718(.A(new_n661), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n913), .B(KEYINPUT45), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(KEYINPUT104), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n654), .A2(KEYINPUT104), .A3(new_n660), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n660), .B(new_n662), .Z(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n654), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT103), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n703), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n667), .B(KEYINPUT41), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n706), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n919), .A2(new_n912), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n912), .A2(new_n664), .A3(KEYINPUT42), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT42), .B1(new_n912), .B2(new_n664), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n629), .B1(new_n600), .B2(new_n562), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n936), .B(new_n937), .C1(new_n649), .C2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n941), .B1(new_n939), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n909), .B1(new_n933), .B2(new_n948), .ZN(G387));
  AND2_X1   g0749(.A1(new_n925), .A2(new_n929), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(new_n703), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n703), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n667), .A3(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n736), .A2(G326), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n886), .A2(G283), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G311), .A2(new_n723), .B1(new_n718), .B2(G317), .ZN(new_n956));
  INV_X1    g0756(.A(G322), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n956), .B1(new_n957), .B2(new_n743), .C1(new_n466), .C2(new_n741), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT48), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n955), .B1(new_n728), .B2(new_n739), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT108), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n959), .B2(new_n958), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n264), .B1(new_n446), .B2(new_n733), .C1(new_n962), .C2(KEYINPUT49), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n954), .B(new_n963), .C1(KEYINPUT49), .C2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n886), .A2(new_n421), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n202), .B2(new_n717), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT107), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n741), .A2(new_n208), .ZN(new_n968));
  INV_X1    g0768(.A(new_n739), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G159), .A2(new_n744), .B1(new_n969), .B2(new_n220), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n348), .B2(new_n735), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n354), .B1(new_n733), .B2(new_n378), .C1(new_n325), .C2(new_n722), .ZN(new_n972));
  NOR4_X1   g0772(.A1(new_n967), .A2(new_n968), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n714), .B1(new_n964), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n325), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n202), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n977));
  AOI21_X1  g0777(.A(G45), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n670), .B(new_n979), .C1(G68), .C2(G77), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n758), .B(new_n980), .C1(G45), .C2(new_n244), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n670), .A2(new_n229), .A3(new_n354), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(G107), .B2(new_n229), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT106), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n763), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n660), .A2(new_n711), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n974), .A2(new_n707), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n953), .B(new_n987), .C1(new_n705), .C2(new_n930), .ZN(G393));
  NAND3_X1  g0788(.A1(new_n917), .A2(new_n706), .A3(new_n921), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n912), .A2(new_n711), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n763), .B1(new_n378), .B2(new_n229), .C1(new_n758), .C2(new_n254), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n739), .A2(new_n208), .B1(new_n735), .B2(new_n895), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT109), .Z(new_n993));
  NAND2_X1  g0793(.A1(new_n792), .A2(new_n975), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n743), .A2(new_n348), .B1(new_n717), .B2(new_n748), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT51), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n730), .A2(new_n402), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n354), .B1(new_n733), .B2(new_n217), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(G50), .C2(new_n723), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n993), .A2(new_n994), .A3(new_n996), .A4(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT110), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n741), .A2(new_n728), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n739), .A2(new_n790), .B1(new_n735), .B2(new_n957), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n465), .C2(new_n723), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n743), .A2(new_n724), .B1(new_n717), .B2(new_n740), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT52), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n354), .B1(new_n886), .B2(G116), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1006), .A3(new_n746), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1001), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n708), .B1(new_n1009), .B2(new_n714), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n990), .A2(new_n991), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n989), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n989), .A2(KEYINPUT111), .A3(new_n1011), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n922), .A2(new_n952), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n668), .B1(new_n952), .B2(new_n922), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1019), .ZN(G390));
  AND3_X1   g0820(.A1(new_n698), .A2(new_n700), .A3(new_n801), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT112), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1021), .A2(new_n1022), .A3(G330), .A4(new_n808), .ZN(new_n1023));
  INV_X1    g0823(.A(G330), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT112), .B1(new_n809), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n863), .B1(new_n870), .B2(new_n808), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n850), .B2(new_n862), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n649), .B(new_n774), .C1(new_n681), .C2(new_n638), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n437), .A2(new_n649), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n808), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n863), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n837), .A2(new_n838), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1023), .B(new_n1025), .C1(new_n1027), .C2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n824), .A2(new_n827), .A3(new_n851), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT39), .B1(new_n837), .B2(new_n838), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1035), .A2(new_n1036), .B1(new_n863), .B2(new_n871), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1030), .A2(new_n1032), .A3(new_n1031), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n698), .A2(new_n700), .A3(new_n653), .A4(new_n801), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n808), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1034), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n706), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n709), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G283), .A2(new_n744), .B1(new_n792), .B2(G97), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n213), .B2(new_n722), .C1(new_n446), .C2(new_n717), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G87), .B2(new_n969), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n997), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n779), .B1(G294), .B2(new_n736), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT114), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n264), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n969), .A2(G150), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n264), .B1(new_n1053), .B2(KEYINPUT53), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(KEYINPUT53), .B2(new_n1053), .C1(new_n748), .C2(new_n730), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G132), .B2(new_n718), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT54), .B(G143), .Z(new_n1057));
  AOI22_X1  g0857(.A1(G137), .A2(new_n723), .B1(new_n792), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT113), .ZN(new_n1059));
  INV_X1    g0859(.A(G128), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n743), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1058), .A2(KEYINPUT113), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G125), .C2(new_n736), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1056), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n733), .A2(new_n202), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1052), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n708), .B1(new_n1066), .B2(new_n714), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1045), .B(new_n1067), .C1(new_n975), .C2(new_n800), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1044), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1023), .A2(new_n1025), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n870), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1041), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1021), .A2(G330), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1073), .B(new_n1074), .C1(new_n1075), .C2(new_n808), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n841), .A2(new_n1024), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n845), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1080), .A2(new_n1034), .A3(new_n1042), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n844), .B(new_n624), .C1(new_n1024), .C2(new_n841), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n668), .B1(new_n1043), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1069), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G378));
  NAND2_X1  g0886(.A1(new_n375), .A2(KEYINPUT55), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT55), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1088), .B(new_n363), .C1(new_n373), .C2(new_n374), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n352), .A2(new_n814), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT56), .Z(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n840), .B2(G330), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n828), .A2(new_n829), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT117), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1091), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(KEYINPUT117), .A3(new_n1092), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1032), .A2(KEYINPUT40), .A3(new_n810), .ZN(new_n1106));
  AND4_X1   g0906(.A1(G330), .A2(new_n1098), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n873), .B1(new_n1097), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT119), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n864), .A2(new_n865), .A3(new_n872), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n809), .B1(new_n849), .B2(new_n838), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1106), .B(G330), .C1(new_n1111), .C2(KEYINPUT40), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1095), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n840), .A2(G330), .A3(new_n1105), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1108), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1027), .A2(new_n1033), .A3(new_n1073), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1083), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1079), .ZN(new_n1121));
  OAI211_X1 g0921(.A(KEYINPUT119), .B(new_n873), .C1(new_n1097), .C2(new_n1107), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1116), .A2(new_n1121), .A3(KEYINPUT57), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1080), .B1(new_n1034), .B2(new_n1042), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1110), .B1(new_n1114), .B2(new_n1113), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1126), .A2(new_n1082), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT57), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n668), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1120), .B2(new_n1079), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1132), .A2(KEYINPUT120), .A3(new_n1116), .A4(new_n1122), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1125), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n734), .A2(G58), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT115), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n274), .C1(new_n221), .C2(new_n739), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n354), .B(new_n1137), .C1(G283), .C2(new_n736), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT116), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G97), .A2(new_n723), .B1(new_n718), .B2(G107), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n446), .B2(new_n743), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G68), .B2(new_n886), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1139), .B(new_n1142), .C1(new_n554), .C2(new_n741), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT58), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n717), .A2(new_n1060), .B1(new_n730), .B2(new_n348), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n969), .A2(new_n1057), .B1(new_n792), .B2(G137), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n787), .B2(new_n722), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(G125), .C2(new_n744), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT59), .ZN(new_n1150));
  AOI21_X1  g0950(.A(G41), .B1(new_n736), .B2(G124), .ZN(new_n1151));
  AOI21_X1  g0951(.A(G33), .B1(new_n734), .B2(G159), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n202), .B1(new_n262), .B2(G41), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1145), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n708), .B1(new_n1156), .B2(new_n714), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(G50), .B2(new_n800), .C1(new_n1105), .C2(new_n710), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT118), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1160), .B2(new_n706), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1134), .A2(new_n1161), .ZN(G375));
  NOR2_X1   g0962(.A1(new_n739), .A2(new_n378), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n743), .A2(new_n728), .B1(new_n735), .B2(new_n738), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(G77), .C2(new_n734), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n718), .A2(G283), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n264), .B1(new_n722), .B2(new_n446), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G107), .B2(new_n792), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n965), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n743), .A2(new_n787), .B1(new_n717), .B2(new_n783), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G150), .B2(new_n792), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n723), .A2(new_n1057), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n264), .B1(new_n886), .B2(G50), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1136), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n739), .A2(new_n748), .B1(new_n735), .B2(new_n1060), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT121), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1169), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n708), .B1(new_n1177), .B2(new_n714), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n808), .B2(new_n710), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n208), .B2(new_n799), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1077), .B2(new_n706), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1082), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n932), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1183), .B2(new_n1083), .ZN(G381));
  NAND3_X1  g0984(.A1(new_n1134), .A2(new_n1085), .A3(new_n1161), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(G387), .A2(G390), .A3(G384), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OR3_X1    g0988(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(KEYINPUT122), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT122), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1188), .A2(new_n1192), .A3(new_n1189), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1191), .A2(new_n1193), .ZN(G407));
  INV_X1    g0994(.A(G213), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(G343), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT123), .B1(new_n1186), .B2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n1195), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1186), .A2(KEYINPUT123), .A3(new_n1196), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n1191), .C2(new_n1193), .ZN(G409));
  NOR2_X1   g1000(.A1(KEYINPUT124), .A2(KEYINPUT63), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1085), .B1(new_n1134), .B2(new_n1161), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1116), .A2(new_n706), .A3(new_n1122), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1121), .A2(new_n1160), .A3(new_n932), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1085), .A2(new_n1158), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1196), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT60), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1182), .A2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1082), .A2(new_n1072), .A3(KEYINPUT60), .A4(new_n1076), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1210), .A2(new_n667), .A3(new_n1080), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1181), .ZN(new_n1213));
  INV_X1    g1013(.A(G384), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(G384), .A3(new_n1181), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1203), .A2(new_n1208), .A3(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(KEYINPUT124), .A2(KEYINPUT63), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1202), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G375), .A2(G378), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1208), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1196), .A2(G2897), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1217), .B2(KEYINPUT125), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1217), .A2(KEYINPUT125), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1217), .A2(KEYINPUT125), .A3(new_n1225), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT61), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n931), .A2(new_n932), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n947), .B1(new_n1232), .B2(new_n706), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n909), .A3(G390), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1014), .A2(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT126), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(G393), .B(new_n768), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1233), .A2(G390), .A3(KEYINPUT126), .A4(new_n909), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT127), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT127), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1238), .A2(new_n1240), .A3(new_n1243), .A4(new_n1239), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1234), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(new_n1239), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1236), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1217), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1221), .A2(new_n1222), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1201), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1220), .A2(new_n1231), .A3(new_n1249), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1208), .B1(G375), .B2(G378), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1255), .B2(new_n1250), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1203), .A2(KEYINPUT62), .A3(new_n1208), .A4(new_n1217), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1253), .B1(new_n1261), .B2(new_n1249), .ZN(G405));
  OAI21_X1  g1062(.A(new_n1250), .B1(new_n1186), .B2(new_n1203), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1221), .A2(new_n1185), .A3(new_n1217), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(new_n1249), .ZN(G402));
endmodule


