//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n190), .B(new_n192), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT0), .B(G128), .Z(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n193), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT0), .B(G128), .C1(new_n203), .C2(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  MUX2_X1   g020(.A(new_n199), .B(new_n206), .S(G125), .Z(new_n207));
  INV_X1    g021(.A(G224), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G953), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n207), .B(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n211));
  XNOR2_X1  g025(.A(G110), .B(G122), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT77), .A2(G104), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT77), .A2(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT77), .A2(G104), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT77), .A2(G104), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G107), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n214), .A3(G104), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n219), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n217), .B1(G104), .B2(new_n214), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT66), .A2(G116), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(G119), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n232), .B2(G119), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n239), .A3(G119), .A4(new_n234), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n230), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n229), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(G116), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT66), .A2(G116), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n236), .B1(new_n247), .B2(G119), .ZN(new_n248));
  INV_X1    g062(.A(new_n240), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n251), .A3(new_n240), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n244), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G113), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n232), .A2(G119), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(new_n244), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT79), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n238), .A2(new_n251), .A3(new_n240), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n251), .B1(new_n238), .B2(new_n240), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT5), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT79), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(new_n256), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n243), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n250), .A2(new_n230), .A3(new_n252), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n242), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n220), .A2(new_n221), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n223), .B1(new_n268), .B2(new_n214), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n222), .A2(new_n224), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n267), .B(G101), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(G101), .B1(new_n269), .B2(new_n270), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n266), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n211), .B(new_n213), .C1(new_n264), .C2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT6), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n258), .A2(new_n263), .ZN(new_n277));
  INV_X1    g091(.A(new_n243), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n274), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n212), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT80), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n273), .A2(new_n271), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n277), .A2(new_n278), .B1(new_n266), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n212), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n280), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n213), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n282), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n210), .B1(new_n276), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n285), .B1(new_n284), .B2(new_n212), .ZN(new_n292));
  NOR4_X1   g106(.A1(new_n264), .A2(new_n274), .A3(KEYINPUT80), .A4(new_n213), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n241), .B1(new_n258), .B2(new_n263), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n238), .A2(new_n240), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n257), .B1(new_n296), .B2(KEYINPUT5), .ZN(new_n297));
  OAI22_X1  g111(.A1(new_n295), .A2(new_n229), .B1(new_n243), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n212), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT7), .B1(new_n208), .B2(G953), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n207), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n291), .B1(new_n294), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n188), .B1(new_n290), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n210), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n212), .B1(new_n279), .B2(new_n280), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n292), .A2(new_n293), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n287), .A2(new_n211), .A3(KEYINPUT6), .A4(new_n213), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT6), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n275), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n282), .A2(new_n286), .ZN(new_n315));
  INV_X1    g129(.A(new_n303), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n298), .B2(new_n300), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n187), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n306), .A2(KEYINPUT83), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT83), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n321), .B(new_n188), .C1(new_n290), .C2(new_n305), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT9), .B(G234), .ZN(new_n325));
  OAI21_X1  g139(.A(G221), .B1(new_n325), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G469), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(new_n291), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n273), .A2(new_n206), .A3(new_n271), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n199), .A2(new_n225), .A3(new_n227), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT10), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT11), .ZN(new_n334));
  INV_X1    g148(.A(G134), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(G137), .ZN(new_n336));
  INV_X1    g150(.A(G137), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT11), .A3(G134), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(G137), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G131), .ZN(new_n341));
  INV_X1    g155(.A(G131), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n336), .A2(new_n338), .A3(new_n342), .A4(new_n339), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n199), .A2(new_n225), .A3(new_n227), .A4(KEYINPUT10), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n330), .A2(new_n333), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G953), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G227), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT76), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G140), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n330), .A2(new_n333), .A3(new_n345), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n341), .A2(new_n343), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n330), .A2(new_n333), .A3(new_n358), .A4(new_n345), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n228), .A2(new_n198), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n331), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT12), .B1(new_n362), .B2(new_n357), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT12), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n364), .B(new_n344), .C1(new_n361), .C2(new_n331), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n346), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n354), .A2(new_n360), .B1(new_n366), .B2(new_n353), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n329), .B1(new_n367), .B2(G469), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n352), .B1(new_n360), .B2(new_n346), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n363), .A2(new_n365), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n370), .A2(new_n353), .A3(new_n347), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n328), .B(new_n291), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n327), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(G113), .B(G122), .Z(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(G104), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n348), .A3(G214), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(new_n191), .ZN(new_n381));
  NOR2_X1   g195(.A1(G237), .A2(G953), .ZN(new_n382));
  AOI21_X1  g196(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n378), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT18), .A2(G131), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n191), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(KEYINPUT85), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT73), .A2(G125), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(KEYINPUT73), .A2(G125), .A3(G140), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G146), .ZN(new_n396));
  XNOR2_X1  g210(.A(G125), .B(G140), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n189), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n381), .A2(new_n383), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n385), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n387), .A2(new_n388), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n403), .A2(KEYINPUT86), .A3(new_n386), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n390), .B(new_n399), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G131), .B1(new_n381), .B2(new_n383), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n387), .A2(new_n342), .A3(new_n388), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n394), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n392), .A2(G125), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g225(.A(G146), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n397), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n408), .B(new_n412), .C1(new_n416), .C2(G146), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n377), .B1(new_n405), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n406), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n406), .A2(new_n407), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(new_n419), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n394), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(new_n189), .C1(KEYINPUT16), .C2(new_n410), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n409), .A2(new_n411), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT74), .A3(new_n189), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n385), .B1(new_n403), .B2(new_n378), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n430), .A2(new_n389), .B1(new_n398), .B2(new_n396), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n401), .A2(new_n400), .A3(new_n385), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT86), .B1(new_n403), .B2(new_n386), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n422), .A2(new_n429), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n418), .B1(new_n435), .B2(new_n377), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT88), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n375), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  INV_X1    g254(.A(new_n438), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n422), .A2(new_n429), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n442), .A2(new_n377), .A3(new_n405), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n440), .B(new_n441), .C1(new_n443), .C2(new_n418), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n435), .A2(new_n377), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n291), .B1(new_n446), .B2(new_n443), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT89), .B(G475), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT13), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n196), .B2(G143), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n191), .A2(KEYINPUT13), .A3(G128), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n196), .A2(G143), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT90), .A4(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n455), .B(G134), .C1(KEYINPUT90), .C2(new_n453), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n191), .A2(G128), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n454), .A3(new_n335), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n233), .A2(G122), .A3(new_n234), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n232), .A2(G122), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n214), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n459), .A2(new_n214), .A3(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n456), .B(new_n458), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n214), .A3(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n457), .A2(new_n454), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G134), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n458), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n459), .A2(new_n468), .A3(new_n460), .ZN(new_n469));
  OAI21_X1  g283(.A(G107), .B1(new_n459), .B2(new_n468), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n464), .B(new_n467), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G217), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n325), .A2(new_n473), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n463), .A2(new_n471), .A3(new_n474), .ZN(new_n477));
  AOI21_X1  g291(.A(G902), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT15), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT91), .Z(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT92), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n484));
  INV_X1    g298(.A(new_n478), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(new_n480), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n348), .A2(G952), .ZN(new_n488));
  INV_X1    g302(.A(G234), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n488), .B1(new_n489), .B2(new_n379), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n291), .B(new_n348), .C1(G234), .C2(G237), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT21), .B(G898), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n450), .A2(new_n487), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n373), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n323), .A2(KEYINPUT93), .A3(new_n324), .A4(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n320), .A2(new_n324), .A3(new_n322), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n373), .A2(new_n495), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT75), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n505));
  INV_X1    g319(.A(G119), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(G128), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n507), .B(new_n508), .C1(G119), .C2(new_n196), .ZN(new_n509));
  XNOR2_X1  g323(.A(G119), .B(G128), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT24), .B(G110), .Z(new_n511));
  AOI22_X1  g325(.A1(new_n509), .A2(G110), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n426), .A2(new_n428), .A3(new_n512), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n509), .A2(G110), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n412), .A3(new_n398), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n348), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n513), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n513), .B2(new_n515), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT25), .A3(new_n291), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n515), .ZN(new_n523));
  INV_X1    g337(.A(new_n518), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n515), .A3(new_n518), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n291), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n473), .B1(G234), .B2(new_n291), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n504), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n531), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n522), .B2(new_n529), .ZN(new_n537));
  INV_X1    g351(.A(new_n534), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n537), .A2(KEYINPUT75), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n543));
  XOR2_X1   g357(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n544));
  NAND2_X1  g358(.A1(new_n382), .A2(G210), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT26), .B(G101), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n357), .A2(new_n204), .A3(new_n202), .ZN(new_n550));
  INV_X1    g364(.A(new_n339), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n335), .A2(G137), .ZN(new_n552));
  OAI21_X1  g366(.A(G131), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n195), .A2(new_n553), .A3(new_n343), .A4(new_n197), .ZN(new_n554));
  AND4_X1   g368(.A1(new_n265), .A2(new_n242), .A3(new_n550), .A4(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n265), .A2(new_n242), .B1(new_n550), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n549), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n265), .A2(new_n242), .A3(new_n550), .A4(new_n554), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT28), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n548), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n259), .A2(new_n260), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n241), .B1(new_n562), .B2(new_n230), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n554), .B1(new_n344), .B2(new_n205), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT65), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n550), .A2(new_n565), .A3(new_n566), .A4(new_n554), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n563), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n548), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n573), .A2(new_n574), .A3(new_n555), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n543), .A2(new_n561), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n549), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n266), .A2(new_n564), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(new_n558), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n558), .A2(new_n559), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n543), .B(new_n574), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n567), .B(new_n569), .C1(new_n550), .C2(new_n554), .ZN(new_n583));
  INV_X1    g397(.A(new_n572), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n266), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(new_n576), .A3(new_n548), .A4(new_n558), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n542), .B1(new_n577), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n548), .A3(new_n558), .ZN(new_n590));
  AOI22_X1  g404(.A1(KEYINPUT71), .A2(new_n589), .B1(new_n590), .B2(KEYINPUT31), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n582), .A2(new_n586), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT72), .ZN(new_n593));
  NOR2_X1   g407(.A1(G472), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n588), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT32), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n573), .A2(new_n555), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n574), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT29), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n557), .A2(new_n548), .A3(new_n560), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n579), .A2(new_n558), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT28), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n560), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n548), .A2(KEYINPUT29), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n602), .B(new_n291), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n595), .A2(new_n596), .B1(new_n607), .B2(G472), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n588), .A2(new_n593), .A3(KEYINPUT32), .A4(new_n594), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n541), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n503), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  NAND3_X1  g426(.A1(new_n306), .A2(KEYINPUT94), .A3(new_n319), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n614), .B(new_n188), .C1(new_n290), .C2(new_n305), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n475), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n476), .A2(new_n477), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n476), .B2(new_n477), .ZN(new_n620));
  OAI21_X1  g434(.A(G478), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n479), .A2(new_n291), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n478), .B2(new_n479), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n450), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n494), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n613), .A2(new_n324), .A3(new_n615), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n588), .A2(new_n593), .A3(new_n291), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n595), .ZN(new_n632));
  INV_X1    g446(.A(new_n373), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n632), .A2(new_n633), .A3(new_n541), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT96), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  AND3_X1   g452(.A1(new_n613), .A2(new_n324), .A3(new_n615), .ZN(new_n639));
  INV_X1    g453(.A(new_n487), .ZN(new_n640));
  INV_X1    g454(.A(new_n439), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n436), .A2(new_n375), .A3(new_n438), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n449), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n640), .A2(new_n643), .A3(new_n494), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n639), .A2(new_n634), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NOR2_X1   g461(.A1(new_n524), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n523), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n533), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n532), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n503), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND2_X1  g470(.A1(new_n595), .A2(new_n596), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n607), .A2(G472), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n609), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(new_n613), .A3(new_n324), .A4(new_n615), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n633), .A2(new_n652), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n491), .B1(new_n492), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n640), .A2(new_n643), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n196), .ZN(G30));
  XNOR2_X1  g481(.A(new_n323), .B(KEYINPUT38), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n597), .A2(new_n574), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n291), .B1(new_n603), .B2(new_n548), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT97), .Z(new_n672));
  NAND3_X1  g486(.A1(new_n657), .A2(new_n609), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n663), .B(KEYINPUT39), .Z(new_n674));
  AND2_X1   g488(.A1(new_n373), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n324), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n439), .A2(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n651), .A2(new_n640), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n673), .A2(new_n677), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n668), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT98), .B(G143), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G45));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n624), .B1(new_n445), .B2(new_n449), .ZN(new_n687));
  INV_X1    g501(.A(new_n663), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n686), .A3(new_n688), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n633), .A3(new_n652), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n639), .A2(KEYINPUT100), .A3(new_n659), .A4(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n695));
  INV_X1    g509(.A(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n661), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n695), .B1(new_n660), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  OAI21_X1  g514(.A(new_n291), .B1(new_n369), .B2(new_n371), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n326), .A3(new_n372), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n702), .A2(new_n705), .A3(new_n326), .A4(new_n372), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n659), .A2(new_n540), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n629), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT102), .B1(new_n707), .B2(new_n628), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND4_X1  g528(.A1(new_n613), .A2(new_n324), .A3(new_n615), .A4(new_n644), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n707), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n232), .ZN(G18));
  INV_X1    g531(.A(new_n703), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n613), .A2(new_n324), .A3(new_n718), .A4(new_n615), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n659), .A2(new_n495), .A3(new_n651), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n506), .ZN(G21));
  XOR2_X1   g536(.A(new_n594), .B(KEYINPUT103), .Z(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n574), .A2(new_n605), .B1(new_n590), .B2(KEYINPUT31), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n725), .A2(new_n726), .B1(new_n576), .B2(new_n575), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n729), .B1(new_n631), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n537), .A2(new_n538), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n630), .A2(KEYINPUT105), .A3(G472), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n732), .A4(new_n733), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n640), .A2(new_n679), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n613), .A2(new_n324), .A3(new_n615), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n704), .A2(new_n706), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n740), .A2(new_n494), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND2_X1  g558(.A1(new_n631), .A2(new_n730), .ZN(new_n745));
  INV_X1    g559(.A(new_n729), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n651), .A3(new_n733), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT107), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n731), .A2(new_n749), .A3(new_n651), .A4(new_n733), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n719), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n696), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  AOI21_X1  g568(.A(new_n678), .B1(new_n320), .B2(new_n322), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n367), .A2(G469), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n329), .B(KEYINPUT108), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n372), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n326), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n755), .A2(new_n610), .A3(new_n696), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n609), .A2(KEYINPUT109), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n609), .A2(KEYINPUT109), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n608), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n732), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n678), .B(new_n759), .C1(new_n320), .C2(new_n322), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n692), .A2(new_n762), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NAND4_X1  g586(.A1(new_n755), .A2(new_n610), .A3(new_n664), .A4(new_n760), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n625), .B1(new_n679), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n776), .B2(new_n679), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n679), .A2(new_n779), .A3(new_n625), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n775), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(KEYINPUT113), .B(new_n781), .C1(new_n778), .C2(new_n779), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n652), .B1(new_n631), .B2(new_n595), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n783), .A2(KEYINPUT44), .A3(new_n784), .A4(new_n785), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n755), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(G469), .B1(new_n367), .B2(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT110), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT110), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n793), .B(G469), .C1(new_n367), .C2(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n367), .A2(KEYINPUT45), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n796), .B2(new_n757), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n372), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n326), .A3(new_n674), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n337), .ZN(G39));
  INV_X1    g618(.A(new_n755), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n805), .A2(new_n659), .A3(new_n540), .A4(new_n692), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n801), .A2(KEYINPUT47), .A3(new_n326), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT47), .B1(new_n801), .B2(new_n326), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NOR2_X1   g625(.A1(new_n651), .A2(new_n663), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n758), .A3(new_n326), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n671), .B(KEYINPUT97), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n595), .B2(new_n596), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n813), .B1(new_n815), .B2(new_n609), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n639), .A2(KEYINPUT115), .A3(new_n816), .A4(new_n739), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n673), .A2(new_n760), .A3(new_n812), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n818), .B1(new_n740), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n666), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n753), .A2(new_n699), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n497), .B(new_n501), .C1(new_n610), .C2(new_n653), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n540), .A2(new_n373), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n687), .A2(new_n827), .B1(new_n679), .B2(new_n487), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n626), .A2(KEYINPUT114), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n494), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n826), .A2(new_n595), .A3(new_n830), .A4(new_n631), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n707), .A2(new_n715), .B1(new_n499), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n721), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n712), .A2(new_n825), .A3(new_n743), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n692), .B1(new_n748), .B2(new_n750), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n768), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n643), .A2(new_n487), .A3(new_n663), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n755), .A2(new_n659), .A3(new_n661), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n773), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n771), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n666), .B1(new_n835), .B2(new_n752), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n699), .A4(new_n821), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n824), .A2(new_n834), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n712), .A2(new_n825), .A3(new_n743), .A4(new_n833), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n771), .A2(new_n836), .A3(new_n839), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n841), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n845), .B1(new_n851), .B2(KEYINPUT52), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n852), .A3(new_n843), .A4(new_n824), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n846), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n845), .B1(new_n841), .B2(new_n842), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n850), .A2(new_n856), .A3(new_n843), .A4(new_n824), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n847), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT116), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n858), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n854), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n808), .A2(new_n809), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n702), .A2(new_n372), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n864), .B1(new_n326), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n780), .A2(new_n782), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n738), .A2(new_n491), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n866), .A2(new_n755), .A3(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n805), .A2(new_n490), .A3(new_n703), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n751), .A3(new_n867), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n673), .A2(new_n541), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n870), .A2(new_n679), .A3(new_n624), .A4(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n668), .A2(new_n324), .A3(new_n703), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n874), .A2(KEYINPUT50), .A3(new_n868), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT50), .B1(new_n874), .B2(new_n868), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n871), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n878));
  OR3_X1    g692(.A1(new_n869), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n878), .B1(new_n869), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n868), .A2(new_n752), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n870), .A2(new_n687), .A3(new_n872), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n488), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n870), .A2(new_n767), .A3(new_n867), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT48), .Z(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n879), .A2(new_n880), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n863), .A2(new_n890), .B1(G952), .B2(G953), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n865), .A2(KEYINPUT49), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n865), .A2(KEYINPUT49), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n537), .A2(new_n538), .A3(new_n678), .A4(new_n327), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n892), .A2(new_n778), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n668), .A2(new_n673), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n891), .A2(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n348), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n291), .B1(new_n846), .B2(new_n853), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n309), .A2(new_n313), .A3(new_n307), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n290), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n899), .B1(new_n901), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n904), .B1(new_n901), .B2(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT118), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n904), .C1(new_n901), .C2(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n912), .B2(new_n914), .ZN(G51));
  NAND2_X1  g729(.A1(new_n846), .A2(new_n853), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n854), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n757), .B(KEYINPUT57), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n369), .B2(new_n371), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n900), .A2(new_n794), .A3(new_n795), .A4(new_n792), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n898), .B1(new_n921), .B2(new_n922), .ZN(G54));
  INV_X1    g737(.A(new_n436), .ZN(new_n924));
  AND2_X1   g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n900), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n900), .B2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n898), .ZN(G60));
  OR2_X1    g742(.A1(new_n619), .A2(new_n620), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n622), .Z(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n918), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n899), .ZN(new_n934));
  INV_X1    g748(.A(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n863), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n936), .B2(new_n929), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n916), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n521), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n916), .A2(KEYINPUT122), .A3(new_n940), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT122), .B1(new_n916), .B2(new_n940), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n942), .B(new_n939), .C1(new_n846), .C2(new_n853), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n649), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(new_n949), .A3(new_n899), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT61), .A4(new_n899), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  OAI21_X1  g768(.A(G953), .B1(new_n493), .B2(new_n208), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n834), .B2(G953), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n276), .B(new_n289), .C1(G898), .C2(new_n348), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n571), .A2(new_n572), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(new_n416), .Z(new_n961));
  NAND2_X1  g775(.A1(new_n841), .A2(new_n699), .ZN(new_n962));
  OR3_X1    g776(.A1(new_n962), .A2(new_n683), .A3(KEYINPUT62), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT62), .B1(new_n962), .B2(new_n683), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n828), .A2(new_n829), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n610), .A2(new_n675), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n803), .B1(new_n755), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n963), .A2(new_n810), .A3(new_n964), .A4(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n968), .B2(new_n348), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n959), .B1(new_n969), .B2(KEYINPUT123), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT123), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n662), .A2(G953), .ZN(new_n972));
  INV_X1    g786(.A(new_n802), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n767), .A2(new_n639), .A3(new_n739), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n810), .A2(new_n771), .A3(new_n773), .A4(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n803), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n977), .A2(new_n978), .A3(new_n699), .A4(new_n841), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT126), .B1(new_n803), .B2(new_n962), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n972), .B1(new_n981), .B2(G953), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n971), .B1(new_n982), .B2(new_n961), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n970), .B1(new_n983), .B2(new_n969), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n348), .B1(G227), .B2(G900), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT124), .Z(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(new_n981), .A2(new_n834), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  AOI211_X1 g804(.A(new_n548), .B(new_n598), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n990), .B1(new_n968), .B2(new_n848), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n992), .A2(new_n669), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n599), .B(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n590), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n990), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n846), .B2(new_n857), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n991), .A2(new_n993), .A3(new_n898), .A4(new_n997), .ZN(G57));
endmodule


