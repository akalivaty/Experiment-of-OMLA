//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n221), .A2(new_n222), .A3(new_n207), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n205), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n218), .ZN(new_n232));
  AND3_X1   g0032(.A1(new_n220), .A2(new_n228), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n207), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT69), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n225), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT68), .B1(new_n254), .B2(new_n225), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n225), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(KEYINPUT69), .A3(new_n255), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n249), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n252), .B1(new_n264), .B2(new_n207), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n262), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n267));
  INV_X1    g0067(.A(G150), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n226), .A2(G33), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n267), .B1(new_n268), .B2(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n266), .A2(new_n273), .A3(KEYINPUT70), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n265), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n278), .A2(KEYINPUT9), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(KEYINPUT9), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G223), .B1(G77), .B2(new_n285), .ZN(new_n288));
  INV_X1    g0088(.A(G222), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n286), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT67), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G33), .A3(G41), .ZN(new_n301));
  INV_X1    g0101(.A(new_n225), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n295), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n305), .B2(G226), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n294), .A2(G190), .A3(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n279), .A2(new_n280), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n294), .A2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT74), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n308), .B(new_n310), .C1(new_n311), .C2(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n279), .A2(new_n280), .A3(new_n310), .A4(new_n307), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n279), .A2(new_n280), .A3(new_n311), .A4(new_n307), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n278), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n317), .B(new_n319), .C1(G179), .C2(new_n309), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n312), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n290), .A2(G232), .A3(G1698), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT75), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT75), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n290), .A2(new_n325), .A3(G232), .A4(G1698), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n290), .A2(G226), .A3(new_n286), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n293), .ZN(new_n330));
  INV_X1    g0130(.A(new_n297), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n304), .B2(new_n216), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n322), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  AOI211_X1 g0134(.A(KEYINPUT13), .B(new_n332), .C1(new_n329), .C2(new_n293), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G169), .B1(new_n334), .B2(new_n335), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(KEYINPUT14), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n338), .A2(KEYINPUT14), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n272), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(G77), .B1(G20), .B2(new_n215), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n207), .B2(new_n270), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n266), .A2(KEYINPUT11), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n251), .A2(new_n215), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT12), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n261), .A2(new_n255), .ZN(new_n348));
  INV_X1    g0148(.A(new_n263), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G68), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n345), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT11), .B1(new_n266), .B2(new_n344), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n341), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n330), .A2(new_n333), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT13), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n330), .A2(new_n322), .A3(new_n333), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G190), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(G200), .B1(new_n334), .B2(new_n335), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n354), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT76), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n360), .A2(new_n361), .A3(new_n364), .A4(new_n354), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n356), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n331), .B1(new_n304), .B2(new_n214), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n287), .A2(KEYINPUT77), .A3(G226), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT77), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n290), .A2(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n208), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n290), .A2(G223), .A3(new_n286), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  XOR2_X1   g0173(.A(new_n373), .B(KEYINPUT78), .Z(new_n374));
  NAND4_X1  g0174(.A1(new_n368), .A2(new_n371), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n367), .B1(new_n375), .B2(new_n293), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G179), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n318), .B2(new_n376), .ZN(new_n378));
  XNOR2_X1  g0178(.A(G58), .B(G68), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT7), .B1(new_n285), .B2(new_n226), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n382), .B(G20), .C1(new_n282), .C2(new_n284), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n380), .B1(new_n384), .B2(new_n215), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT16), .B(new_n380), .C1(new_n384), .C2(new_n215), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n348), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n271), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n264), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n390), .B2(new_n251), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n378), .A2(KEYINPUT18), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT18), .B1(new_n378), .B2(new_n393), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n375), .A2(new_n293), .ZN(new_n397));
  OAI21_X1  g0197(.A(G200), .B1(new_n397), .B2(new_n367), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n376), .A2(G190), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(new_n389), .A3(new_n392), .A4(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n350), .A2(G77), .ZN(new_n402));
  XOR2_X1   g0202(.A(new_n402), .B(KEYINPUT73), .Z(new_n403));
  INV_X1    g0203(.A(KEYINPUT72), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT15), .B(G87), .Z(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n404), .B1(new_n406), .B2(new_n272), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(KEYINPUT72), .A3(new_n342), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n390), .A2(new_n269), .B1(G20), .B2(G77), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G77), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n410), .A2(new_n348), .B1(new_n411), .B2(new_n251), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n293), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n285), .A2(G107), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n415), .B1(new_n291), .B2(new_n214), .C1(new_n216), .C2(new_n370), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(KEYINPUT71), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(KEYINPUT71), .B2(new_n416), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n297), .B1(new_n305), .B2(G244), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n413), .B1(new_n420), .B2(G190), .ZN(new_n421));
  INV_X1    g0221(.A(G200), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(new_n420), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n336), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n413), .C1(G169), .C2(new_n420), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n396), .A2(new_n401), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n321), .A2(new_n366), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G45), .ZN(new_n429));
  OAI21_X1  g0229(.A(G250), .B1(new_n429), .B2(G1), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n225), .B1(KEYINPUT67), .B2(new_n298), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(new_n301), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n429), .A2(new_n296), .A3(G1), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT81), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n282), .A2(new_n284), .A3(G238), .A4(new_n286), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(G1698), .ZN(new_n436));
  INV_X1    g0236(.A(G116), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n281), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n293), .ZN(new_n441));
  INV_X1    g0241(.A(new_n430), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n303), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT81), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n429), .A2(G1), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G274), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n434), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G190), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT83), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n446), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(KEYINPUT81), .B1(new_n293), .B2(new_n440), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT83), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(G190), .A4(new_n447), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT84), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n454), .A3(KEYINPUT84), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n282), .A2(new_n284), .A3(new_n226), .A4(G68), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n272), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(KEYINPUT19), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT82), .B(G87), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G97), .A2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n463), .A2(new_n464), .B1(new_n226), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n348), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n406), .A2(new_n251), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n249), .A2(G33), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n250), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n258), .A2(new_n262), .A3(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n467), .B(new_n468), .C1(new_n471), .C2(new_n209), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(G200), .B2(new_n448), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n457), .A2(new_n458), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n467), .A2(new_n468), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n406), .B2(new_n471), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n448), .A2(new_n318), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n452), .A2(new_n336), .A3(new_n447), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n282), .A2(new_n284), .A3(new_n226), .A4(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n290), .A2(new_n483), .A3(new_n226), .A4(G87), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n226), .B2(G107), .ZN(new_n487));
  INV_X1    g0287(.A(G107), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT23), .A3(G20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n438), .A2(new_n226), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT88), .B(KEYINPUT24), .C1(new_n485), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT88), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n482), .B2(new_n484), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n496), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n348), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n290), .A2(G250), .A3(new_n286), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n290), .A2(G257), .A3(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G294), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n293), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT89), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n507), .A3(new_n293), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n445), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n303), .A2(new_n511), .A3(G264), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n433), .B1(new_n510), .B2(new_n509), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n506), .A2(new_n449), .A3(new_n508), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n505), .A2(new_n513), .A3(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n422), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n471), .A2(new_n488), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n250), .A2(G107), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n520), .B(KEYINPUT25), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n500), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n506), .A2(new_n508), .A3(new_n514), .ZN(new_n525));
  INV_X1    g0325(.A(new_n516), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(G169), .B1(new_n526), .B2(G179), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n522), .B1(new_n499), .B2(new_n348), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(new_n286), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n536), .A2(new_n293), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n509), .A2(new_n510), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n446), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n303), .A2(new_n511), .A3(G257), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT80), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n303), .A2(new_n511), .A3(KEYINPUT80), .A4(G257), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(G200), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n250), .A2(G97), .ZN(new_n546));
  OAI21_X1  g0346(.A(G107), .B1(new_n381), .B2(new_n383), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n548), .A2(G97), .A3(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n460), .A2(KEYINPUT6), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT79), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(G107), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n488), .A2(KEYINPUT79), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n549), .A2(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n464), .A2(KEYINPUT6), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n548), .A2(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n488), .A2(KEYINPUT79), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(G107), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n554), .A2(G20), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n269), .A2(G77), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n547), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n546), .B1(new_n562), .B2(new_n348), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n258), .A2(new_n262), .A3(G97), .A4(new_n470), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n536), .A2(new_n293), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n565), .A2(G190), .A3(new_n543), .A4(new_n542), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n545), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n560), .A2(new_n561), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n382), .B1(new_n290), .B2(G20), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n488), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n348), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n546), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n564), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n318), .B1(new_n537), .B2(new_n544), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n565), .A2(new_n336), .A3(new_n543), .A4(new_n542), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n282), .A2(new_n284), .A3(G257), .A4(new_n286), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT85), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n290), .A2(KEYINPUT85), .A3(G257), .A4(new_n286), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n290), .A2(G264), .A3(G1698), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n285), .A2(G303), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n293), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n303), .A2(new_n511), .A3(G270), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n513), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n256), .A2(new_n257), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n250), .A2(G116), .A3(new_n469), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n591), .A2(new_n593), .B1(new_n437), .B2(new_n251), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n254), .A2(new_n225), .B1(G20), .B2(new_n437), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n534), .B(new_n226), .C1(G33), .C2(new_n460), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(KEYINPUT20), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n318), .B1(new_n594), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n590), .A2(new_n602), .A3(KEYINPUT86), .A4(KEYINPUT21), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n595), .A2(KEYINPUT20), .A3(new_n596), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT20), .B1(new_n595), .B2(new_n596), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n348), .A2(new_n592), .B1(G116), .B2(new_n250), .ZN(new_n607));
  OAI21_X1  g0407(.A(G169), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n588), .B1(new_n585), .B2(new_n293), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT86), .B1(new_n610), .B2(KEYINPUT21), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n594), .A2(new_n601), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n614), .A3(G179), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n586), .A2(G190), .A3(new_n589), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n606), .A2(new_n607), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n609), .A2(new_n422), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT87), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n609), .B2(G190), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n590), .A2(G200), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n578), .A2(new_n603), .A3(new_n617), .A4(new_n627), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n428), .A2(new_n480), .A3(new_n529), .A4(new_n628), .ZN(G372));
  AND3_X1   g0429(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n474), .A2(new_n479), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n473), .A2(new_n455), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n630), .A2(new_n633), .A3(new_n634), .A4(new_n479), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n635), .A2(new_n479), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n632), .A2(new_n636), .A3(KEYINPUT90), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n633), .A2(new_n479), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n524), .A3(new_n578), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n528), .A2(new_n527), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n590), .A2(new_n602), .A3(KEYINPUT21), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT86), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n603), .A3(new_n615), .A4(new_n613), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n639), .A2(new_n640), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n427), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT91), .Z(new_n652));
  INV_X1    g0452(.A(new_n362), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n356), .B1(new_n653), .B2(new_n425), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n401), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n396), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n312), .A3(new_n316), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n320), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n659), .ZN(G369));
  NOR3_X1   g0460(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT87), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n625), .B1(new_n623), .B2(new_n624), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n647), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n226), .A2(G13), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n249), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n619), .ZN(new_n673));
  MUX2_X1   g0473(.A(new_n664), .B(new_n647), .S(new_n673), .Z(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n525), .A2(G169), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n526), .A2(G179), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n499), .A2(new_n348), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n678), .B(new_n671), .C1(new_n679), .C2(new_n522), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n528), .A2(new_n672), .ZN(new_n681));
  OAI211_X1 g0481(.A(KEYINPUT92), .B(new_n680), .C1(new_n529), .C2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n678), .B1(new_n679), .B2(new_n522), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n671), .B1(new_n679), .B2(new_n522), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n524), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT92), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n675), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n647), .A2(new_n672), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n683), .B2(new_n687), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n684), .A2(new_n671), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n690), .A2(new_n693), .A3(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n229), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n223), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n698), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G1), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n463), .A2(new_n437), .A3(new_n464), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n650), .A2(new_n672), .ZN(new_n705));
  INV_X1    g0505(.A(new_n479), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n448), .A2(G200), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n707), .B(new_n475), .C1(new_n471), .C2(new_n209), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n456), .B2(new_n455), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n706), .B1(new_n709), .B2(new_n458), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n634), .A3(new_n630), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n641), .A2(new_n630), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n706), .B1(new_n712), .B2(KEYINPUT26), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n649), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(new_n672), .ZN(new_n715));
  MUX2_X1   g0515(.A(new_n705), .B(new_n715), .S(KEYINPUT29), .Z(new_n716));
  NOR2_X1   g0516(.A1(new_n609), .A2(G179), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n565), .A2(new_n543), .A3(new_n542), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n448), .A3(new_n516), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT93), .Z(new_n720));
  INV_X1    g0520(.A(new_n718), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n505), .A2(new_n512), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n448), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n721), .A2(new_n723), .A3(G179), .A4(new_n609), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT30), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n672), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n567), .A2(new_n577), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n663), .A2(new_n647), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n529), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n728), .A2(new_n710), .A3(new_n729), .A4(new_n672), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n730), .B2(KEYINPUT31), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n732), .B(new_n672), .C1(new_n725), .C2(new_n719), .ZN(new_n733));
  OAI21_X1  g0533(.A(G330), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n716), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n704), .B1(new_n736), .B2(G1), .ZN(G364));
  AOI21_X1  g0537(.A(new_n249), .B1(new_n665), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n698), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n675), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G330), .B2(new_n674), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n697), .A2(new_n285), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G355), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G116), .B2(new_n229), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n224), .A2(new_n429), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n285), .A2(new_n229), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n247), .B2(G45), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n225), .B1(G20), .B2(new_n318), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n740), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n226), .A2(G190), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT94), .Z(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT95), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT96), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT96), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n336), .A2(G200), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n768), .A2(KEYINPUT99), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(KEYINPUT99), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n765), .A2(G329), .B1(new_n772), .B2(G283), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n336), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n757), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n285), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n226), .A2(new_n449), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n774), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G322), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n336), .A2(new_n422), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G326), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n757), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT33), .B(G317), .Z(new_n786));
  OAI221_X1 g0586(.A(new_n781), .B1(new_n783), .B2(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n767), .A2(new_n778), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n777), .B(new_n787), .C1(G303), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G294), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n760), .A2(G190), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n773), .B(new_n790), .C1(new_n791), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n764), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n772), .A2(G107), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n793), .A2(G97), .ZN(new_n801));
  INV_X1    g0601(.A(new_n785), .ZN(new_n802));
  INV_X1    g0602(.A(new_n775), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G68), .A2(new_n802), .B1(new_n803), .B2(G77), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n213), .B2(new_n779), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n788), .A2(new_n463), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n290), .B1(new_n783), .B2(new_n207), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n800), .A2(new_n801), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n795), .B1(new_n799), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n756), .B1(new_n810), .B2(new_n753), .ZN(new_n811));
  INV_X1    g0611(.A(new_n752), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n674), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n742), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NOR2_X1   g0615(.A1(new_n425), .A2(new_n671), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n413), .A2(new_n671), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n423), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n425), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n705), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n650), .A2(new_n672), .A3(new_n819), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n740), .B1(new_n823), .B2(new_n734), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n734), .B2(new_n823), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n772), .A2(G87), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n776), .B2(new_n764), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n789), .A2(G107), .ZN(new_n828));
  INV_X1    g0628(.A(G303), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n783), .A2(new_n829), .B1(new_n779), .B2(new_n791), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G116), .B2(new_n803), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n290), .B1(new_n802), .B2(G283), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n801), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n771), .A2(new_n215), .B1(new_n834), .B2(new_n764), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n836), .A2(new_n779), .B1(new_n785), .B2(new_n268), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n783), .A2(new_n838), .B1(new_n775), .B2(new_n796), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(KEYINPUT34), .B1(new_n793), .B2(G58), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n285), .B1(new_n789), .B2(G50), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(KEYINPUT34), .C2(new_n840), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n827), .A2(new_n833), .B1(new_n835), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n753), .ZN(new_n845));
  INV_X1    g0645(.A(new_n740), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n753), .A2(new_n750), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n411), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n845), .B(new_n848), .C1(new_n819), .C2(new_n751), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n825), .A2(new_n849), .ZN(G384));
  NAND2_X1  g0650(.A1(new_n554), .A2(new_n559), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT35), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n554), .A2(KEYINPUT35), .A3(new_n559), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(new_n854), .A3(G116), .A4(new_n227), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT36), .Z(new_n856));
  OAI211_X1 g0656(.A(new_n223), .B(G77), .C1(new_n213), .C2(new_n215), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n207), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n249), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G330), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT17), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n376), .A2(new_n422), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G190), .B2(new_n376), .ZN(new_n864));
  INV_X1    g0664(.A(new_n393), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n400), .A2(KEYINPUT17), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n866), .A2(new_n867), .B1(new_n394), .B2(new_n395), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n387), .A2(new_n266), .A3(new_n388), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n392), .ZN(new_n870));
  INV_X1    g0670(.A(new_n669), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n378), .A2(new_n393), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n393), .A2(new_n871), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n875), .A2(new_n400), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n378), .A2(new_n870), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n879), .A2(new_n400), .A3(new_n872), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n880), .B2(new_n877), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n874), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n363), .A2(new_n365), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n355), .B(new_n671), .C1(new_n885), .C2(new_n341), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n653), .B1(new_n355), .B2(new_n671), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n356), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n726), .A2(KEYINPUT31), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n819), .B(new_n889), .C1(new_n731), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(KEYINPUT101), .A2(KEYINPUT40), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n884), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n726), .ZN(new_n895));
  NOR4_X1   g0695(.A1(new_n628), .A2(new_n480), .A3(new_n529), .A4(new_n671), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n732), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n726), .A2(KEYINPUT31), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n899), .A2(new_n819), .A3(new_n889), .A4(new_n892), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n891), .A2(KEYINPUT101), .ZN(new_n901));
  XNOR2_X1  g0701(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n876), .B1(new_n396), .B2(new_n401), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n875), .A2(new_n400), .A3(new_n876), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n878), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n902), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n900), .A2(new_n901), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n894), .B1(new_n910), .B2(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n899), .A2(new_n427), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT102), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n861), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  INV_X1    g0715(.A(new_n714), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT29), .B1(new_n916), .B2(new_n671), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(KEYINPUT29), .B2(new_n705), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n658), .B1(new_n918), .B2(new_n427), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n915), .B(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n907), .A2(new_n921), .A3(new_n908), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n874), .A2(new_n881), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n921), .B1(new_n925), .B2(new_n908), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n356), .A2(new_n671), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n927), .A2(new_n929), .B1(new_n396), .B2(new_n871), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n642), .A2(new_n648), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n637), .B2(new_n638), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n671), .B1(new_n932), .B2(new_n640), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n816), .B1(new_n933), .B2(new_n819), .ZN(new_n934));
  INV_X1    g0734(.A(new_n889), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n934), .A2(new_n884), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n920), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n249), .B2(new_n665), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n920), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n860), .B1(new_n939), .B2(new_n940), .ZN(G367));
  NOR2_X1   g0741(.A1(new_n240), .A2(new_n747), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n754), .B1(new_n229), .B2(new_n406), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n740), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n472), .A2(new_n671), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n479), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n641), .A2(new_n945), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n947), .B2(KEYINPUT103), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(KEYINPUT103), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n812), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n285), .B1(new_n783), .B2(new_n776), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n791), .A2(new_n785), .B1(new_n779), .B2(new_n829), .ZN(new_n952));
  INV_X1    g0752(.A(new_n768), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n951), .B(new_n952), .C1(new_n953), .C2(G97), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n789), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n788), .B2(new_n437), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G317), .B2(new_n765), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n793), .A2(G107), .B1(G283), .B2(new_n803), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT108), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n765), .A2(G137), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n953), .A2(G77), .B1(G58), .B2(new_n789), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n794), .A2(new_n215), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n290), .B1(new_n785), .B2(new_n796), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G150), .A2(new_n780), .B1(new_n803), .B2(G50), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n836), .B2(new_n783), .ZN(new_n969));
  NOR4_X1   g0769(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n959), .A2(new_n962), .B1(new_n963), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n753), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n971), .B2(new_n973), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n944), .B(new_n950), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n698), .B(KEYINPUT41), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n675), .A2(new_n688), .A3(new_n692), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n688), .B1(new_n675), .B2(new_n692), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n716), .A2(new_n734), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n574), .A2(new_n671), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n567), .A2(new_n577), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT105), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n630), .A2(new_n671), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n984), .B2(new_n985), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT106), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n578), .A2(KEYINPUT105), .A3(new_n983), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT106), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n991), .A2(new_n992), .A3(new_n986), .A4(new_n988), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n680), .B1(new_n529), .B2(new_n681), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT92), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n691), .B1(new_n997), .B2(new_n682), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n994), .B1(new_n998), .B2(new_n694), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n994), .B(KEYINPUT44), .C1(new_n998), .C2(new_n694), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n990), .A2(new_n993), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n693), .A2(new_n695), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n695), .A4(new_n1004), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1003), .A2(new_n1009), .A3(new_n690), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT107), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1001), .A2(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(KEYINPUT107), .A3(new_n690), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n982), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n978), .B1(new_n1015), .B2(new_n735), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n738), .ZN(new_n1017));
  OR3_X1    g0817(.A1(new_n693), .A2(new_n994), .A3(KEYINPUT42), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n577), .B1(new_n994), .B2(new_n684), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n672), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT42), .B1(new_n693), .B2(new_n994), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT104), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n690), .A2(new_n994), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1028), .A2(new_n1031), .A3(new_n1029), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n977), .B1(new_n1017), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(G387));
  AND3_X1   g0838(.A1(new_n716), .A2(new_n734), .A3(new_n981), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n700), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n736), .B2(new_n981), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n743), .A2(new_n702), .B1(new_n488), .B2(new_n697), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n702), .C1(G68), .C2(G77), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n271), .A2(G50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n747), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT110), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1046), .A2(new_n1047), .B1(new_n429), .B2(new_n237), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n846), .B1(new_n1050), .B2(new_n754), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n785), .A2(new_n271), .B1(new_n775), .B2(new_n215), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT111), .Z(new_n1053));
  AOI22_X1  g0853(.A1(new_n765), .A2(G150), .B1(new_n772), .B2(G97), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n793), .A2(new_n405), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n290), .B1(new_n779), .B2(new_n207), .C1(new_n796), .C2(new_n783), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G77), .B2(new_n789), .ZN(new_n1057));
  AND4_X1   g0857(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n783), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1059), .A2(G322), .B1(new_n803), .B2(G303), .ZN(new_n1060));
  INV_X1    g0860(.A(G317), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n776), .B2(new_n785), .C1(new_n1061), .C2(new_n779), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT48), .ZN(new_n1063));
  INV_X1    g0863(.A(G283), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n794), .C1(new_n791), .C2(new_n788), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n285), .B1(new_n437), .B2(new_n768), .C1(new_n764), .C2(new_n784), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1058), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1051), .B1(new_n1070), .B2(new_n975), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n688), .B2(new_n752), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n981), .B2(new_n739), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1041), .A2(new_n1073), .ZN(G393));
  NOR2_X1   g0874(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT107), .B1(new_n1013), .B2(new_n690), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1039), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1013), .A2(new_n690), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1077), .B(new_n698), .C1(new_n1079), .C2(new_n1039), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT114), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n244), .A2(new_n747), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n754), .B1(new_n460), .B2(new_n229), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n740), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1004), .A2(new_n812), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n285), .B1(new_n775), .B2(new_n791), .C1(new_n829), .C2(new_n785), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n783), .A2(new_n1061), .B1(new_n779), .B2(new_n776), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT52), .Z(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(G283), .C2(new_n789), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n765), .A2(G322), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n793), .A2(G116), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n800), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n285), .B1(new_n789), .B2(G68), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n826), .B(new_n1093), .C1(new_n836), .C2(new_n764), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT112), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n793), .A2(G77), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n207), .B2(new_n785), .C1(new_n271), .C2(new_n775), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1098), .A2(KEYINPUT113), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n783), .A2(new_n268), .B1(new_n779), .B2(new_n796), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT51), .Z(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1096), .B(new_n1102), .C1(KEYINPUT113), .C2(new_n1098), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1084), .B(new_n1085), .C1(new_n753), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1079), .B2(new_n739), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1080), .A2(new_n1081), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1081), .B1(new_n1080), .B2(new_n1107), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G390));
  INV_X1    g0911(.A(new_n816), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n935), .B1(new_n822), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n927), .B1(new_n1113), .B2(new_n928), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n819), .C1(new_n731), .C2(new_n733), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1115), .A2(new_n935), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n818), .A2(new_n425), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n714), .A2(new_n672), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n935), .B1(new_n1118), .B2(new_n1112), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n909), .A2(new_n929), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1114), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n899), .A2(G330), .A3(new_n819), .A4(new_n889), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n739), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n846), .B1(new_n271), .B2(new_n847), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n771), .A2(new_n215), .B1(new_n791), .B2(new_n764), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n789), .A2(G87), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n290), .B1(new_n802), .B2(G107), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n779), .A2(new_n437), .B1(new_n775), .B2(new_n460), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G283), .B2(new_n1059), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1129), .A2(new_n1097), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT118), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n285), .B1(new_n780), .B2(G132), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n783), .C1(new_n768), .C2(new_n207), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n765), .B2(G125), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n788), .A2(new_n268), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT54), .B(G143), .Z(new_n1142));
  AOI22_X1  g0942(.A1(G137), .A2(new_n802), .B1(new_n803), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n794), .B2(new_n796), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT117), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1135), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(KEYINPUT118), .B2(new_n1134), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n922), .A2(new_n926), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1127), .B1(new_n975), .B2(new_n1148), .C1(new_n1149), .C2(new_n751), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1126), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n820), .B1(new_n897), .B2(new_n898), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n889), .B1(new_n1153), .B2(G330), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1112), .B(new_n1118), .C1(new_n1115), .C2(new_n935), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1115), .A2(new_n935), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1123), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n822), .A2(new_n1112), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1159), .A2(KEYINPUT115), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT115), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n899), .A2(new_n427), .A3(G330), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n659), .B(new_n1164), .C1(new_n716), .C2(new_n428), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n928), .B1(new_n1160), .B2(new_n889), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1116), .B(new_n1121), .C1(new_n1168), .C2(new_n1149), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n927), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1169), .B1(new_n1172), .B2(new_n1123), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1115), .A2(new_n935), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n891), .A2(new_n861), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1160), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT115), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1159), .A2(KEYINPUT115), .A3(new_n1160), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1165), .B1(new_n1181), .B2(new_n1157), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n700), .B1(new_n1182), .B2(new_n1125), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT116), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1174), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n698), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(KEYINPUT116), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1152), .B1(new_n1185), .B2(new_n1187), .ZN(G378));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT120), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n321), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n278), .A2(new_n669), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n312), .A2(KEYINPUT120), .A3(new_n316), .A4(new_n320), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1194), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1190), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1198), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1189), .A3(new_n1196), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n911), .B2(new_n861), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT40), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n891), .A2(KEYINPUT101), .B1(new_n908), .B2(new_n907), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n900), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1202), .B(G330), .C1(new_n1207), .C2(new_n894), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n937), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1204), .A2(new_n937), .A3(new_n1208), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1203), .A2(new_n750), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n847), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n740), .B1(G50), .B2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G97), .A2(new_n802), .B1(new_n803), .B2(new_n405), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n488), .B2(new_n779), .C1(new_n437), .C2(new_n783), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n966), .B(new_n1218), .C1(G58), .C2(new_n953), .ZN(new_n1219));
  INV_X1    g1019(.A(G41), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n285), .C1(new_n788), .C2(new_n411), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT119), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1219), .B(new_n1222), .C1(new_n1064), .C2(new_n764), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT58), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G50), .B1(new_n281), .B2(new_n1220), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n290), .B2(G41), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1059), .A2(G125), .B1(new_n802), .B2(G132), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G128), .A2(new_n780), .B1(new_n803), .B2(G137), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1142), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1229), .B1(new_n788), .B2(new_n1230), .C1(new_n794), .C2(new_n268), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  AOI211_X1 g1033(.A(G33), .B(G41), .C1(new_n953), .C2(G159), .ZN(new_n1234));
  INV_X1    g1034(.A(G124), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1233), .B(new_n1234), .C1(new_n1235), .C2(new_n764), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1224), .B(new_n1226), .C1(new_n1232), .C2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1216), .B1(new_n1237), .B2(new_n753), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1213), .A2(new_n739), .B1(new_n1214), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1156), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1166), .B1(new_n1173), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1204), .A2(new_n937), .A3(new_n1208), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n937), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(KEYINPUT57), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n698), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1241), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n1245), .B2(new_n1246), .ZN(G375));
  OAI211_X1 g1047(.A(new_n1165), .B(new_n1157), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1167), .A2(new_n978), .A3(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n764), .A2(new_n829), .B1(new_n771), .B2(new_n411), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n789), .A2(G97), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n783), .A2(new_n791), .B1(new_n779), .B2(new_n1064), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G107), .B2(new_n803), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n290), .B1(new_n802), .B2(G116), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1251), .A2(new_n1055), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n764), .A2(new_n1137), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n953), .A2(G58), .B1(G159), .B2(new_n789), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n783), .A2(new_n834), .B1(new_n779), .B2(new_n838), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n290), .B1(new_n1230), .B2(new_n785), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(G150), .C2(new_n803), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1257), .B(new_n1260), .C1(new_n207), .C2(new_n794), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1250), .A2(new_n1255), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n753), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1263), .B(new_n740), .C1(G68), .C2(new_n1215), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n935), .B2(new_n750), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1163), .B2(new_n739), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1266), .ZN(G381));
  INV_X1    g1067(.A(new_n1124), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1169), .A2(new_n1268), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1186), .B2(KEYINPUT116), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1151), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT57), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n698), .A3(new_n1244), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1272), .A2(new_n1276), .A3(new_n1239), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1080), .A2(new_n1107), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT114), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1080), .A2(new_n1081), .A3(new_n1107), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1037), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1041), .A2(new_n814), .A3(new_n1073), .ZN(new_n1282));
  OR3_X1    g1082(.A1(G381), .A2(G384), .A3(new_n1282), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1277), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT121), .Z(G407));
  OAI211_X1 g1085(.A(G407), .B(G213), .C1(G343), .C2(new_n1277), .ZN(G409));
  INV_X1    g1086(.A(KEYINPUT125), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G375), .A2(G378), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n670), .A2(G213), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1241), .B(new_n978), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n739), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1214), .A2(new_n1238), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1290), .B1(new_n1272), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1248), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1240), .A2(KEYINPUT60), .A3(new_n1165), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n698), .A4(new_n1167), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(G384), .A3(new_n1266), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G384), .B1(new_n1299), .B2(new_n1266), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1288), .A2(new_n1295), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT63), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1288), .A2(new_n1295), .A3(new_n1306), .A4(new_n1303), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1272), .B1(new_n1239), .B2(new_n1276), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1289), .B1(G378), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT122), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT122), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1288), .A2(new_n1295), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1290), .A2(G2897), .ZN(new_n1316));
  XOR2_X1   g1116(.A(new_n1316), .B(KEYINPUT123), .Z(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1299), .A2(new_n1266), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1300), .A3(new_n1317), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1313), .A2(new_n1315), .A3(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1308), .A2(new_n1309), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1035), .B1(new_n738), .B2(new_n1016), .ZN(new_n1327));
  OAI22_X1  g1127(.A1(new_n1108), .A2(new_n1109), .B1(new_n1327), .B2(new_n977), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(new_n1281), .A3(KEYINPUT124), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G393), .A2(G396), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1282), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1328), .A2(new_n1281), .A3(KEYINPUT124), .A4(new_n1331), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1326), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1304), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1304), .A2(new_n1338), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1324), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1336), .A2(KEYINPUT61), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1287), .B1(new_n1337), .B2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1335), .B1(new_n1346), .B2(new_n1325), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1342), .A2(new_n1335), .A3(new_n1309), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1348), .B1(new_n1340), .B2(new_n1339), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1347), .A2(KEYINPUT125), .A3(new_n1349), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1345), .A2(new_n1350), .ZN(G405));
  NAND2_X1  g1151(.A1(new_n1288), .A2(new_n1277), .ZN(new_n1352));
  XOR2_X1   g1152(.A(new_n1352), .B(new_n1303), .Z(new_n1353));
  NAND3_X1  g1153(.A1(new_n1353), .A2(KEYINPUT126), .A3(new_n1335), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1335), .B(KEYINPUT126), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1354), .B1(new_n1355), .B2(new_n1353), .ZN(G402));
endmodule


