

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731;

  INV_X1 U371 ( .A(n705), .ZN(n349) );
  NAND2_X1 U372 ( .A1(n429), .A2(n430), .ZN(n512) );
  XNOR2_X1 U373 ( .A(G128), .B(KEYINPUT77), .ZN(n427) );
  AND2_X2 U374 ( .A1(n350), .A2(n349), .ZN(n364) );
  XNOR2_X1 U375 ( .A(n403), .B(n351), .ZN(n350) );
  INV_X1 U376 ( .A(n361), .ZN(n351) );
  NOR2_X2 U377 ( .A1(G902), .A2(n686), .ZN(n450) );
  XOR2_X1 U378 ( .A(G113), .B(G104), .Z(n508) );
  NOR2_X2 U379 ( .A1(n591), .A2(n570), .ZN(n571) );
  XNOR2_X2 U380 ( .A(n380), .B(KEYINPUT0), .ZN(n592) );
  XNOR2_X2 U381 ( .A(n605), .B(n604), .ZN(n675) );
  NOR2_X1 U382 ( .A1(n644), .A2(n645), .ZN(n641) );
  XNOR2_X1 U383 ( .A(n608), .B(n607), .ZN(n719) );
  NAND2_X1 U384 ( .A1(n400), .A2(n398), .ZN(n608) );
  NAND2_X1 U385 ( .A1(n588), .A2(n585), .ZN(n424) );
  XNOR2_X1 U386 ( .A(KEYINPUT31), .B(n593), .ZN(n631) );
  XNOR2_X1 U387 ( .A(n576), .B(KEYINPUT22), .ZN(n583) );
  XNOR2_X1 U388 ( .A(n539), .B(KEYINPUT106), .ZN(n627) );
  XNOR2_X1 U389 ( .A(n408), .B(n356), .ZN(n644) );
  XNOR2_X1 U390 ( .A(n491), .B(n490), .ZN(n548) );
  XNOR2_X1 U391 ( .A(n435), .B(n434), .ZN(n511) );
  XNOR2_X1 U392 ( .A(n586), .B(KEYINPUT64), .ZN(n423) );
  XNOR2_X1 U393 ( .A(G119), .B(KEYINPUT5), .ZN(n436) );
  INV_X2 U394 ( .A(G953), .ZN(n723) );
  XNOR2_X1 U395 ( .A(n352), .B(n353), .ZN(n383) );
  NAND2_X1 U396 ( .A1(n394), .A2(n404), .ZN(n352) );
  XOR2_X1 U397 ( .A(n452), .B(KEYINPUT62), .Z(n353) );
  XNOR2_X2 U398 ( .A(n448), .B(n447), .ZN(n717) );
  XNOR2_X2 U399 ( .A(n415), .B(n416), .ZN(n711) );
  XOR2_X1 U400 ( .A(KEYINPUT4), .B(G146), .Z(n514) );
  XNOR2_X1 U401 ( .A(n514), .B(G131), .ZN(n431) );
  NOR2_X1 U402 ( .A1(n608), .A2(n379), .ZN(n378) );
  XNOR2_X1 U403 ( .A(n388), .B(KEYINPUT70), .ZN(n433) );
  INV_X1 U404 ( .A(KEYINPUT3), .ZN(n388) );
  NOR2_X1 U405 ( .A1(n637), .A2(n355), .ZN(n371) );
  XNOR2_X1 U406 ( .A(n374), .B(n373), .ZN(n716) );
  INV_X1 U407 ( .A(KEYINPUT10), .ZN(n373) );
  XNOR2_X1 U408 ( .A(G140), .B(G125), .ZN(n374) );
  XOR2_X1 U409 ( .A(KEYINPUT96), .B(KEYINPUT9), .Z(n497) );
  XNOR2_X1 U410 ( .A(n411), .B(n410), .ZN(n499) );
  INV_X1 U411 ( .A(KEYINPUT8), .ZN(n410) );
  NAND2_X1 U412 ( .A1(n723), .A2(G234), .ZN(n411) );
  INV_X1 U413 ( .A(G143), .ZN(n426) );
  XOR2_X1 U414 ( .A(KEYINPUT92), .B(G122), .Z(n486) );
  XNOR2_X1 U415 ( .A(G143), .B(G131), .ZN(n485) );
  XOR2_X1 U416 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n483) );
  XNOR2_X1 U417 ( .A(n514), .B(n515), .ZN(n387) );
  XNOR2_X1 U418 ( .A(n386), .B(n385), .ZN(n384) );
  XNOR2_X1 U419 ( .A(KEYINPUT17), .B(KEYINPUT75), .ZN(n386) );
  XNOR2_X1 U420 ( .A(G125), .B(KEYINPUT18), .ZN(n385) );
  XNOR2_X1 U421 ( .A(n511), .B(n402), .ZN(n401) );
  XNOR2_X1 U422 ( .A(n439), .B(n440), .ZN(n402) );
  XNOR2_X1 U423 ( .A(n470), .B(n367), .ZN(n366) );
  INV_X1 U424 ( .A(G128), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n407), .B(n527), .ZN(n563) );
  NOR2_X1 U426 ( .A1(n551), .A2(n657), .ZN(n407) );
  NAND2_X1 U427 ( .A1(n425), .A2(n627), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n541), .B(KEYINPUT19), .ZN(n568) );
  NAND2_X1 U429 ( .A1(n414), .A2(n412), .ZN(n576) );
  INV_X1 U430 ( .A(n592), .ZN(n414) );
  XNOR2_X1 U431 ( .A(n528), .B(KEYINPUT99), .ZN(n539) );
  OR2_X1 U432 ( .A1(n701), .A2(G902), .ZN(n408) );
  INV_X1 U433 ( .A(G472), .ZN(n395) );
  AND2_X1 U434 ( .A1(G953), .A2(G902), .ZN(n458) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n481) );
  INV_X1 U436 ( .A(KEYINPUT85), .ZN(n434) );
  NOR2_X1 U437 ( .A1(n639), .A2(n399), .ZN(n398) );
  XNOR2_X1 U438 ( .A(n369), .B(n359), .ZN(n400) );
  INV_X1 U439 ( .A(n638), .ZN(n399) );
  XNOR2_X1 U440 ( .A(G101), .B(G104), .ZN(n441) );
  XOR2_X1 U441 ( .A(G110), .B(G107), .Z(n442) );
  INV_X1 U442 ( .A(KEYINPUT89), .ZN(n446) );
  OR2_X1 U443 ( .A1(G237), .A2(G902), .ZN(n518) );
  XNOR2_X1 U444 ( .A(G902), .B(KEYINPUT15), .ZN(n611) );
  NOR2_X1 U445 ( .A1(n548), .A2(n547), .ZN(n505) );
  INV_X1 U446 ( .A(n645), .ZN(n413) );
  XOR2_X1 U447 ( .A(KEYINPUT7), .B(KEYINPUT95), .Z(n493) );
  XNOR2_X1 U448 ( .A(KEYINPUT94), .B(KEYINPUT98), .ZN(n492) );
  XNOR2_X1 U449 ( .A(n498), .B(n363), .ZN(n501) );
  XNOR2_X1 U450 ( .A(G116), .B(KEYINPUT97), .ZN(n496) );
  XNOR2_X1 U451 ( .A(n489), .B(n488), .ZN(n694) );
  XNOR2_X1 U452 ( .A(n711), .B(n417), .ZN(n680) );
  INV_X1 U453 ( .A(n512), .ZN(n513) );
  XNOR2_X1 U454 ( .A(n387), .B(n384), .ZN(n516) );
  OR2_X1 U455 ( .A1(n719), .A2(n675), .ZN(n376) );
  INV_X1 U456 ( .A(n372), .ZN(n558) );
  XNOR2_X1 U457 ( .A(n396), .B(KEYINPUT72), .ZN(n551) );
  XNOR2_X1 U458 ( .A(n504), .B(G478), .ZN(n538) );
  NOR2_X1 U459 ( .A1(n699), .A2(G902), .ZN(n504) );
  XNOR2_X1 U460 ( .A(n409), .B(n472), .ZN(n701) );
  XNOR2_X1 U461 ( .A(n471), .B(n480), .ZN(n409) );
  XNOR2_X1 U462 ( .A(n469), .B(n366), .ZN(n471) );
  INV_X1 U463 ( .A(G475), .ZN(n393) );
  INV_X1 U464 ( .A(G210), .ZN(n391) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n729) );
  INV_X1 U466 ( .A(KEYINPUT40), .ZN(n405) );
  NOR2_X1 U467 ( .A1(n537), .A2(n580), .ZN(n637) );
  XNOR2_X1 U468 ( .A(n372), .B(KEYINPUT110), .ZN(n534) );
  NOR2_X1 U469 ( .A1(n543), .A2(n542), .ZN(n625) );
  AND2_X1 U470 ( .A1(n420), .A2(n644), .ZN(n620) );
  XNOR2_X1 U471 ( .A(n579), .B(KEYINPUT65), .ZN(n420) );
  OR2_X1 U472 ( .A1(n583), .A2(n578), .ZN(n579) );
  INV_X1 U473 ( .A(n705), .ZN(n382) );
  AND2_X1 U474 ( .A1(G210), .A2(n518), .ZN(n354) );
  OR2_X1 U475 ( .A1(n556), .A2(n555), .ZN(n355) );
  XOR2_X1 U476 ( .A(KEYINPUT91), .B(n476), .Z(n356) );
  AND2_X2 U477 ( .A1(n404), .A2(n419), .ZN(n357) );
  XOR2_X1 U478 ( .A(n486), .B(n485), .Z(n358) );
  NAND2_X1 U479 ( .A1(n706), .A2(n378), .ZN(n419) );
  XOR2_X1 U480 ( .A(n557), .B(KEYINPUT48), .Z(n359) );
  XNOR2_X1 U481 ( .A(KEYINPUT66), .B(n613), .ZN(n360) );
  XOR2_X1 U482 ( .A(n696), .B(n695), .Z(n361) );
  INV_X1 U483 ( .A(KEYINPUT2), .ZN(n379) );
  AND2_X1 U484 ( .A1(n723), .A2(n379), .ZN(n362) );
  NAND2_X1 U485 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U486 ( .A(n507), .ZN(n363) );
  AND2_X1 U487 ( .A1(n575), .A2(n413), .ZN(n412) );
  INV_X1 U488 ( .A(n675), .ZN(n706) );
  XNOR2_X1 U489 ( .A(n364), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U490 ( .A(n510), .B(n509), .ZN(n415) );
  NAND2_X1 U491 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U492 ( .A(n365), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U493 ( .A1(n685), .A2(n705), .ZN(n365) );
  XNOR2_X2 U494 ( .A(n536), .B(KEYINPUT1), .ZN(n640) );
  XNOR2_X2 U495 ( .A(n450), .B(n451), .ZN(n536) );
  NAND2_X1 U496 ( .A1(n368), .A2(n573), .ZN(n574) );
  XNOR2_X1 U497 ( .A(n572), .B(KEYINPUT34), .ZN(n368) );
  XNOR2_X2 U498 ( .A(n512), .B(G134), .ZN(n495) );
  XNOR2_X1 U499 ( .A(n529), .B(KEYINPUT46), .ZN(n370) );
  NAND2_X1 U500 ( .A1(n389), .A2(n723), .ZN(n377) );
  NAND2_X1 U501 ( .A1(n377), .A2(n375), .ZN(n676) );
  NAND2_X1 U502 ( .A1(n376), .A2(n362), .ZN(n375) );
  NAND2_X1 U503 ( .A1(n568), .A2(n569), .ZN(n380) );
  XNOR2_X1 U504 ( .A(n381), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U505 ( .A(n592), .ZN(n594) );
  XNOR2_X2 U506 ( .A(n495), .B(n431), .ZN(n448) );
  NOR2_X2 U507 ( .A1(n421), .A2(n620), .ZN(n587) );
  NOR2_X1 U508 ( .A1(n389), .A2(n391), .ZN(n390) );
  NOR2_X1 U509 ( .A1(n389), .A2(n393), .ZN(n392) );
  NOR2_X1 U510 ( .A1(n389), .A2(n395), .ZN(n394) );
  INV_X1 U511 ( .A(n419), .ZN(n389) );
  NAND2_X1 U512 ( .A1(n390), .A2(n404), .ZN(n684) );
  NAND2_X1 U513 ( .A1(n392), .A2(n404), .ZN(n403) );
  NAND2_X1 U514 ( .A1(n357), .A2(G478), .ZN(n698) );
  NAND2_X1 U515 ( .A1(n357), .A2(G469), .ZN(n691) );
  NAND2_X1 U516 ( .A1(n357), .A2(G217), .ZN(n702) );
  NAND2_X1 U517 ( .A1(n397), .A2(n526), .ZN(n396) );
  XNOR2_X1 U518 ( .A(n525), .B(n524), .ZN(n397) );
  XNOR2_X1 U519 ( .A(n448), .B(n401), .ZN(n452) );
  NAND2_X2 U520 ( .A1(n418), .A2(n360), .ZN(n404) );
  NAND2_X1 U521 ( .A1(n563), .A2(n539), .ZN(n406) );
  INV_X1 U522 ( .A(n511), .ZN(n416) );
  XNOR2_X1 U523 ( .A(n516), .B(n513), .ZN(n417) );
  NAND2_X1 U524 ( .A1(n609), .A2(n610), .ZN(n418) );
  NAND2_X1 U525 ( .A1(n731), .A2(n422), .ZN(n421) );
  INV_X1 U526 ( .A(n728), .ZN(n422) );
  XNOR2_X2 U527 ( .A(n424), .B(n423), .ZN(n731) );
  XNOR2_X1 U528 ( .A(n684), .B(n683), .ZN(n685) );
  AND2_X1 U529 ( .A1(n584), .A2(n533), .ZN(n425) );
  INV_X1 U530 ( .A(KEYINPUT83), .ZN(n557) );
  INV_X1 U531 ( .A(n532), .ZN(n533) );
  INV_X1 U532 ( .A(n438), .ZN(n439) );
  INV_X1 U533 ( .A(KEYINPUT23), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n468), .B(n446), .ZN(n447) );
  XNOR2_X1 U535 ( .A(n487), .B(n358), .ZN(n488) );
  INV_X1 U536 ( .A(n538), .ZN(n547) );
  XNOR2_X1 U537 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U538 ( .A(n503), .B(n502), .ZN(n699) );
  NOR2_X1 U539 ( .A1(G952), .A2(n723), .ZN(n705) );
  NAND2_X1 U540 ( .A1(n427), .A2(n426), .ZN(n430) );
  INV_X1 U541 ( .A(n427), .ZN(n428) );
  NAND2_X1 U542 ( .A1(n428), .A2(G143), .ZN(n429) );
  XNOR2_X1 U543 ( .A(G116), .B(G101), .ZN(n432) );
  XNOR2_X1 U544 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U545 ( .A(G113), .B(G137), .Z(n437) );
  XNOR2_X1 U546 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U547 ( .A1(n481), .A2(G210), .ZN(n440) );
  XNOR2_X1 U548 ( .A(KEYINPUT69), .B(G469), .ZN(n451) );
  XNOR2_X1 U549 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U550 ( .A(G140), .B(n443), .Z(n445) );
  NAND2_X1 U551 ( .A1(G227), .A2(n723), .ZN(n444) );
  XNOR2_X1 U552 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U553 ( .A(G137), .B(KEYINPUT67), .Z(n468) );
  XNOR2_X1 U554 ( .A(n449), .B(n717), .ZN(n686) );
  NOR2_X1 U555 ( .A1(n452), .A2(G902), .ZN(n453) );
  XNOR2_X2 U556 ( .A(n453), .B(G472), .ZN(n531) );
  XNOR2_X1 U557 ( .A(KEYINPUT104), .B(n531), .ZN(n577) );
  NAND2_X1 U558 ( .A1(n611), .A2(G234), .ZN(n454) );
  XNOR2_X1 U559 ( .A(n454), .B(KEYINPUT20), .ZN(n473) );
  NAND2_X1 U560 ( .A1(G221), .A2(n473), .ZN(n455) );
  XNOR2_X1 U561 ( .A(KEYINPUT21), .B(n455), .ZN(n645) );
  NAND2_X1 U562 ( .A1(G234), .A2(G237), .ZN(n456) );
  XNOR2_X1 U563 ( .A(n456), .B(KEYINPUT14), .ZN(n459) );
  NAND2_X1 U564 ( .A1(G952), .A2(n459), .ZN(n670) );
  NOR2_X1 U565 ( .A1(G953), .A2(n670), .ZN(n457) );
  XNOR2_X1 U566 ( .A(KEYINPUT87), .B(n457), .ZN(n567) );
  INV_X1 U567 ( .A(n567), .ZN(n462) );
  NAND2_X1 U568 ( .A1(n459), .A2(n458), .ZN(n564) );
  XOR2_X1 U569 ( .A(KEYINPUT107), .B(n564), .Z(n460) );
  NOR2_X1 U570 ( .A1(G900), .A2(n460), .ZN(n461) );
  NOR2_X1 U571 ( .A1(n462), .A2(n461), .ZN(n523) );
  NOR2_X1 U572 ( .A1(n645), .A2(n523), .ZN(n463) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(n463), .ZN(n477) );
  XNOR2_X1 U574 ( .A(G146), .B(n716), .ZN(n480) );
  NAND2_X1 U575 ( .A1(n499), .A2(G221), .ZN(n467) );
  XOR2_X1 U576 ( .A(KEYINPUT74), .B(KEYINPUT24), .Z(n465) );
  XOR2_X2 U577 ( .A(G119), .B(G110), .Z(n506) );
  XNOR2_X1 U578 ( .A(n506), .B(KEYINPUT90), .ZN(n464) );
  XNOR2_X1 U579 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U580 ( .A(n467), .B(n466), .ZN(n472) );
  INV_X1 U581 ( .A(n468), .ZN(n469) );
  XOR2_X1 U582 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n475) );
  NAND2_X1 U583 ( .A1(n473), .A2(G217), .ZN(n474) );
  XNOR2_X1 U584 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U585 ( .A1(n477), .A2(n644), .ZN(n532) );
  NOR2_X1 U586 ( .A1(n577), .A2(n532), .ZN(n478) );
  XNOR2_X1 U587 ( .A(KEYINPUT28), .B(n478), .ZN(n479) );
  NAND2_X1 U588 ( .A1(n536), .A2(n479), .ZN(n543) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(G475), .ZN(n491) );
  XNOR2_X1 U590 ( .A(n480), .B(n508), .ZN(n489) );
  NAND2_X1 U591 ( .A1(G214), .A2(n481), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U593 ( .A(n484), .B(KEYINPUT93), .Z(n487) );
  NOR2_X1 U594 ( .A1(G902), .A2(n694), .ZN(n490) );
  XNOR2_X1 U595 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U596 ( .A(n495), .B(n494), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U598 ( .A(G122), .B(G107), .Z(n507) );
  NAND2_X1 U599 ( .A1(n499), .A2(G217), .ZN(n500) );
  XNOR2_X1 U600 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U601 ( .A(KEYINPUT101), .B(n505), .Z(n575) );
  INV_X1 U602 ( .A(n575), .ZN(n660) );
  XOR2_X1 U603 ( .A(KEYINPUT16), .B(n506), .Z(n510) );
  XNOR2_X1 U604 ( .A(n508), .B(n507), .ZN(n509) );
  NAND2_X1 U605 ( .A1(G224), .A2(n723), .ZN(n515) );
  NAND2_X1 U606 ( .A1(n680), .A2(n611), .ZN(n517) );
  XNOR2_X2 U607 ( .A(n517), .B(n354), .ZN(n562) );
  XNOR2_X1 U608 ( .A(n562), .B(KEYINPUT38), .ZN(n657) );
  NAND2_X1 U609 ( .A1(G214), .A2(n518), .ZN(n519) );
  XNOR2_X1 U610 ( .A(KEYINPUT86), .B(n519), .ZN(n530) );
  INV_X1 U611 ( .A(n530), .ZN(n658) );
  NOR2_X1 U612 ( .A1(n657), .A2(n658), .ZN(n520) );
  XNOR2_X1 U613 ( .A(n520), .B(KEYINPUT109), .ZN(n661) );
  NOR2_X1 U614 ( .A1(n660), .A2(n661), .ZN(n521) );
  XNOR2_X1 U615 ( .A(KEYINPUT41), .B(n521), .ZN(n671) );
  NOR2_X1 U616 ( .A1(n543), .A2(n671), .ZN(n522) );
  XNOR2_X1 U617 ( .A(n522), .B(KEYINPUT42), .ZN(n730) );
  NAND2_X1 U618 ( .A1(n536), .A2(n641), .ZN(n596) );
  NOR2_X1 U619 ( .A1(n596), .A2(n523), .ZN(n526) );
  NOR2_X1 U620 ( .A1(n577), .A2(n658), .ZN(n525) );
  XNOR2_X1 U621 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n524) );
  XNOR2_X1 U622 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n527) );
  NAND2_X1 U623 ( .A1(n548), .A2(n538), .ZN(n528) );
  NOR2_X1 U624 ( .A1(n730), .A2(n729), .ZN(n529) );
  NAND2_X1 U625 ( .A1(n562), .A2(n530), .ZN(n541) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n531), .Z(n570) );
  INV_X1 U627 ( .A(n570), .ZN(n584) );
  NOR2_X1 U628 ( .A1(n541), .A2(n534), .ZN(n535) );
  XOR2_X1 U629 ( .A(KEYINPUT36), .B(n535), .Z(n537) );
  INV_X1 U630 ( .A(n640), .ZN(n589) );
  XNOR2_X1 U631 ( .A(KEYINPUT84), .B(n589), .ZN(n580) );
  NOR2_X1 U632 ( .A1(n548), .A2(n538), .ZN(n630) );
  NOR2_X1 U633 ( .A1(n539), .A2(n630), .ZN(n662) );
  NAND2_X1 U634 ( .A1(n662), .A2(KEYINPUT47), .ZN(n540) );
  XNOR2_X1 U635 ( .A(n540), .B(KEYINPUT78), .ZN(n546) );
  INV_X1 U636 ( .A(n568), .ZN(n542) );
  INV_X1 U637 ( .A(n625), .ZN(n544) );
  NAND2_X1 U638 ( .A1(n544), .A2(KEYINPUT47), .ZN(n545) );
  NAND2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n556) );
  NAND2_X1 U640 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U641 ( .A(KEYINPUT105), .B(n549), .ZN(n573) );
  INV_X1 U642 ( .A(n573), .ZN(n550) );
  NOR2_X1 U643 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n562), .A2(n552), .ZN(n624) );
  XOR2_X1 U645 ( .A(n662), .B(KEYINPUT79), .Z(n598) );
  NOR2_X1 U646 ( .A1(n598), .A2(KEYINPUT47), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n625), .A2(n553), .ZN(n554) );
  NAND2_X1 U648 ( .A1(n624), .A2(n554), .ZN(n555) );
  NAND2_X1 U649 ( .A1(n589), .A2(n558), .ZN(n559) );
  NOR2_X1 U650 ( .A1(n658), .A2(n559), .ZN(n560) );
  XNOR2_X1 U651 ( .A(n560), .B(KEYINPUT43), .ZN(n561) );
  NOR2_X1 U652 ( .A1(n562), .A2(n561), .ZN(n639) );
  NAND2_X1 U653 ( .A1(n563), .A2(n630), .ZN(n638) );
  NOR2_X1 U654 ( .A1(G898), .A2(n564), .ZN(n565) );
  XOR2_X1 U655 ( .A(KEYINPUT88), .B(n565), .Z(n566) );
  NAND2_X1 U656 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n641), .A2(n640), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n571), .B(KEYINPUT33), .ZN(n672) );
  NOR2_X1 U659 ( .A1(n592), .A2(n672), .ZN(n572) );
  XNOR2_X1 U660 ( .A(n574), .B(KEYINPUT35), .ZN(n728) );
  NAND2_X1 U661 ( .A1(n589), .A2(n577), .ZN(n578) );
  INV_X1 U662 ( .A(n580), .ZN(n581) );
  NAND2_X1 U663 ( .A1(n644), .A2(n581), .ZN(n582) );
  XNOR2_X1 U664 ( .A(KEYINPUT103), .B(n582), .ZN(n585) );
  NOR2_X2 U665 ( .A1(n584), .A2(n583), .ZN(n588) );
  XNOR2_X1 U666 ( .A(KEYINPUT32), .B(KEYINPUT76), .ZN(n586) );
  XNOR2_X1 U667 ( .A(n587), .B(KEYINPUT44), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U669 ( .A1(n644), .A2(n590), .ZN(n614) );
  NOR2_X1 U670 ( .A1(n531), .A2(n591), .ZN(n652) );
  NAND2_X1 U671 ( .A1(n652), .A2(n594), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n531), .A2(n594), .ZN(n595) );
  NOR2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n616) );
  NOR2_X1 U674 ( .A1(n631), .A2(n616), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n599), .B(KEYINPUT100), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n614), .A2(n600), .ZN(n601) );
  XNOR2_X1 U678 ( .A(KEYINPUT102), .B(n601), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n605) );
  XOR2_X1 U680 ( .A(KEYINPUT82), .B(KEYINPUT45), .Z(n604) );
  NOR2_X2 U681 ( .A1(n675), .A2(n611), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n606), .B(KEYINPUT80), .ZN(n610) );
  INV_X1 U683 ( .A(KEYINPUT81), .ZN(n607) );
  INV_X1 U684 ( .A(n719), .ZN(n609) );
  INV_X1 U685 ( .A(n611), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  XOR2_X1 U687 ( .A(G101), .B(n614), .Z(G3) );
  NAND2_X1 U688 ( .A1(n627), .A2(n616), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n615), .B(G104), .ZN(G6) );
  XOR2_X1 U690 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n618) );
  NAND2_X1 U691 ( .A1(n616), .A2(n630), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U693 ( .A(G107), .B(n619), .ZN(G9) );
  INV_X1 U694 ( .A(n620), .ZN(n621) );
  XNOR2_X1 U695 ( .A(G110), .B(n621), .ZN(G12) );
  XOR2_X1 U696 ( .A(G128), .B(KEYINPUT29), .Z(n623) );
  NAND2_X1 U697 ( .A1(n625), .A2(n630), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(G30) );
  XNOR2_X1 U699 ( .A(G143), .B(n624), .ZN(G45) );
  NAND2_X1 U700 ( .A1(n627), .A2(n625), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(G146), .ZN(G48) );
  XOR2_X1 U702 ( .A(G113), .B(KEYINPUT111), .Z(n629) );
  NAND2_X1 U703 ( .A1(n631), .A2(n627), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(G15) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n632), .B(KEYINPUT112), .ZN(n633) );
  XNOR2_X1 U707 ( .A(G116), .B(n633), .ZN(G18) );
  XOR2_X1 U708 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n635) );
  XNOR2_X1 U709 ( .A(G125), .B(KEYINPUT37), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(G27) );
  XNOR2_X1 U712 ( .A(G134), .B(n638), .ZN(G36) );
  XOR2_X1 U713 ( .A(G140), .B(n639), .Z(G42) );
  NOR2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U715 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT49), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT115), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n648), .A2(n531), .ZN(n649) );
  NOR2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(KEYINPUT51), .ZN(n654) );
  XNOR2_X1 U724 ( .A(KEYINPUT117), .B(n654), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n671), .A2(n655), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n656), .B(KEYINPUT118), .ZN(n667) );
  AND2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n672), .A2(n665), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n668), .B(KEYINPUT52), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U737 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U738 ( .A(KEYINPUT53), .B(n678), .ZN(n679) );
  XNOR2_X1 U739 ( .A(KEYINPUT119), .B(n679), .ZN(G75) );
  INV_X1 U740 ( .A(n680), .ZN(n682) );
  XOR2_X1 U741 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n681) );
  BUF_X1 U742 ( .A(n686), .Z(n690) );
  XOR2_X1 U743 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n688) );
  XNOR2_X1 U744 ( .A(KEYINPUT121), .B(KEYINPUT120), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U746 ( .A(n690), .B(n689), .Z(n692) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U748 ( .A1(n705), .A2(n693), .ZN(G54) );
  XOR2_X1 U749 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n696) );
  XNOR2_X1 U750 ( .A(n694), .B(KEYINPUT123), .ZN(n695) );
  XNOR2_X1 U751 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U752 ( .A1(n705), .A2(n700), .ZN(G63) );
  XNOR2_X1 U753 ( .A(n701), .B(KEYINPUT124), .ZN(n703) );
  XNOR2_X1 U754 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U755 ( .A1(n705), .A2(n704), .ZN(G66) );
  NAND2_X1 U756 ( .A1(n723), .A2(n706), .ZN(n710) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U758 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U759 ( .A1(n708), .A2(G898), .ZN(n709) );
  NAND2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n715) );
  XOR2_X1 U761 ( .A(n711), .B(KEYINPUT125), .Z(n713) );
  NOR2_X1 U762 ( .A1(G898), .A2(n723), .ZN(n712) );
  NOR2_X1 U763 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(G69) );
  XNOR2_X1 U765 ( .A(KEYINPUT126), .B(n716), .ZN(n718) );
  XNOR2_X1 U766 ( .A(n718), .B(n717), .ZN(n721) );
  XNOR2_X1 U767 ( .A(n719), .B(n721), .ZN(n720) );
  NAND2_X1 U768 ( .A1(n720), .A2(n723), .ZN(n726) );
  XNOR2_X1 U769 ( .A(n721), .B(G227), .ZN(n722) );
  NOR2_X1 U770 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U771 ( .A1(G900), .A2(n724), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U773 ( .A(KEYINPUT127), .B(n727), .ZN(G72) );
  XOR2_X1 U774 ( .A(n728), .B(G122), .Z(G24) );
  XOR2_X1 U775 ( .A(n729), .B(G131), .Z(G33) );
  XOR2_X1 U776 ( .A(G137), .B(n730), .Z(G39) );
  XNOR2_X1 U777 ( .A(n731), .B(G119), .ZN(G21) );
endmodule

