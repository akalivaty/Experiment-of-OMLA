//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT75), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G137), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G128), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G119), .B(G128), .ZN(new_n203));
  INV_X1    g017(.A(G110), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT24), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n202), .A2(G110), .B1(new_n203), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT16), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(G140), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n214), .A2(G146), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(G146), .B1(new_n214), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n209), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT74), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n209), .B(KEYINPUT74), .C1(new_n218), .C2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n198), .A2(new_n200), .A3(new_n204), .A4(new_n201), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n203), .B2(new_n208), .ZN(new_n226));
  XNOR2_X1  g040(.A(G125), .B(G140), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n214), .A2(new_n217), .A3(G146), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT76), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT76), .ZN(new_n234));
  AOI211_X1 g048(.A(new_n234), .B(new_n231), .C1(new_n222), .C2(new_n223), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n195), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n231), .B1(new_n222), .B2(new_n223), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n195), .B1(new_n237), .B2(KEYINPUT76), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n188), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n239), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n190), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n214), .A2(new_n217), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n228), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n230), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT74), .B1(new_n247), .B2(new_n209), .ZN(new_n248));
  INV_X1    g062(.A(new_n223), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n232), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n234), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n237), .A2(KEYINPUT76), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n238), .B1(new_n253), .B2(new_n195), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n189), .A2(G902), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n244), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G137), .ZN(new_n264));
  INV_X1    g078(.A(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G134), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n263), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n264), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n269), .B2(new_n264), .ZN(new_n272));
  OAI21_X1  g086(.A(G131), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT67), .B(KEYINPUT11), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT68), .B(G134), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G137), .ZN(new_n277));
  INV_X1    g091(.A(G131), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(G137), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .A4(new_n271), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT69), .B(G131), .C1(new_n270), .C2(new_n272), .ZN(new_n282));
  INV_X1    g096(.A(G143), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G146), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n283), .A3(G146), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n228), .A2(KEYINPUT64), .A3(G143), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT64), .B1(new_n228), .B2(G143), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n285), .B(new_n287), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  NOR2_X1   g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n228), .A2(G143), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n228), .A3(G143), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n295), .A2(new_n297), .B1(new_n283), .B2(G146), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n290), .A2(new_n293), .B1(new_n298), .B2(new_n291), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n281), .A2(new_n282), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n197), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT2), .B(G113), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OR3_X1    g121(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n307), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n306), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT71), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n276), .A2(G137), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n264), .A2(G134), .ZN(new_n314));
  OAI21_X1  g128(.A(G131), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n280), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n294), .A2(KEYINPUT1), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n290), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n298), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n300), .A2(new_n312), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n312), .B1(new_n300), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT28), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(G237), .A2(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G210), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT27), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G101), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n327), .A2(KEYINPUT29), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n335), .A2(new_n188), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n316), .B2(new_n322), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n300), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n300), .A3(KEYINPUT72), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n312), .ZN(new_n344));
  AOI211_X1 g158(.A(KEYINPUT70), .B(KEYINPUT30), .C1(new_n300), .C2(new_n323), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT70), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n300), .A2(new_n323), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n337), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n332), .B1(new_n349), .B2(new_n324), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n327), .A2(new_n334), .ZN(new_n352));
  INV_X1    g166(.A(new_n332), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n336), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n324), .A2(new_n332), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT73), .B(KEYINPUT31), .Z(new_n359));
  NOR2_X1   g173(.A1(new_n348), .A2(new_n345), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n338), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT72), .B1(new_n338), .B2(new_n300), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n344), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n358), .B(new_n359), .C1(new_n360), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n347), .A2(new_n337), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n347), .A2(new_n346), .A3(new_n337), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n312), .B1(new_n341), .B2(new_n342), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n357), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT31), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n356), .B(new_n364), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n373), .A2(G472), .A3(G902), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n355), .A2(G472), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(G472), .A2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(new_n356), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n371), .B1(new_n349), .B2(new_n358), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n373), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n258), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT9), .B(G234), .ZN(new_n382));
  OAI21_X1  g196(.A(G221), .B1(new_n382), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(G107), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n386), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n388), .A2(G104), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n385), .A2(G107), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n296), .B1(G143), .B2(new_n228), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n283), .A2(KEYINPUT66), .A3(G146), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n284), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n318), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n321), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT79), .B1(new_n401), .B2(KEYINPUT10), .ZN(new_n402));
  INV_X1    g216(.A(new_n396), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n295), .A2(new_n297), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n404), .A2(new_n284), .A3(new_n320), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n404), .A2(new_n284), .B1(G128), .B2(new_n317), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n290), .A2(new_n293), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n386), .A2(new_n389), .A3(new_n391), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(G101), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n404), .A2(new_n284), .A3(new_n291), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(G101), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT78), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n299), .A2(new_n420), .A3(new_n421), .A4(new_n414), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n402), .A2(new_n410), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n281), .A2(new_n282), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT80), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n392), .A2(new_n395), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n392), .B2(new_n395), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n396), .A2(KEYINPUT80), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n392), .A2(new_n395), .A3(new_n426), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT81), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n409), .B1(new_n319), .B2(new_n321), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n423), .B(new_n424), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT82), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n424), .A4(new_n423), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n424), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n430), .A2(new_n431), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n407), .B1(new_n448), .B2(new_n322), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT12), .Z(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G110), .B(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n191), .A2(G227), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n453), .B(new_n454), .Z(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT77), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n423), .B1(new_n436), .B2(new_n437), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n447), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT84), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n461), .A3(new_n447), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n455), .B1(new_n440), .B2(new_n445), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n452), .A2(new_n457), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G469), .B1(new_n465), .B2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n451), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n460), .A2(new_n462), .B1(new_n440), .B2(new_n445), .ZN(new_n468));
  INV_X1    g282(.A(new_n455), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G469), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n188), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n384), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G214), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G110), .B(G122), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT8), .Z(new_n477));
  AND3_X1   g291(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT5), .ZN(new_n478));
  OAI21_X1  g292(.A(G113), .B1(new_n301), .B2(KEYINPUT5), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n448), .B(new_n309), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n481));
  OR3_X1    g295(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n481), .B1(new_n478), .B2(new_n479), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n309), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n396), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n477), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n411), .A2(new_n415), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G125), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n319), .A2(new_n321), .A3(new_n212), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n191), .A2(G224), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n488), .B2(new_n489), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n484), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n433), .A2(new_n495), .ZN(new_n496));
  AND4_X1   g310(.A1(new_n421), .A2(new_n308), .A3(new_n414), .A4(new_n311), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n498), .A3(new_n476), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n476), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n484), .B1(new_n429), .B2(new_n432), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n497), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT6), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT6), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n505), .B(new_n501), .C1(new_n502), .C2(new_n497), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n488), .A2(new_n489), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(new_n490), .Z(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G210), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n500), .A2(new_n509), .A3(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n475), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n385), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n218), .A2(new_n219), .ZN(new_n519));
  OR2_X1    g333(.A1(KEYINPUT86), .A2(G143), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(G214), .A3(new_n328), .ZN(new_n521));
  INV_X1    g335(.A(G237), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n191), .A3(G214), .ZN(new_n523));
  NOR2_X1   g337(.A1(KEYINPUT86), .A2(G143), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT17), .A3(G131), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n520), .B1(G214), .B2(new_n328), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n523), .A2(new_n524), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n521), .A2(new_n525), .A3(new_n278), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n519), .B(new_n527), .C1(new_n532), .C2(KEYINPUT17), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT18), .A2(G131), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n521), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n227), .B(new_n228), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n537));
  INV_X1    g351(.A(new_n534), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT87), .B(new_n534), .C1(new_n521), .C2(new_n525), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n535), .B(new_n536), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n518), .B1(new_n542), .B2(KEYINPUT93), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n533), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(KEYINPUT94), .A3(new_n545), .ZN(new_n549));
  INV_X1    g363(.A(new_n518), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n516), .B1(new_n553), .B2(new_n188), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT19), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT88), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n210), .A2(G125), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n215), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n211), .A2(new_n213), .B1(KEYINPUT88), .B2(new_n555), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n228), .C1(new_n559), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT89), .ZN(new_n561));
  INV_X1    g375(.A(new_n556), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n555), .A2(KEYINPUT88), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n562), .B1(new_n227), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n228), .A4(new_n558), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n561), .A2(new_n532), .A3(new_n230), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n541), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT90), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n541), .A3(KEYINPUT90), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n550), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT91), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n570), .A2(new_n574), .A3(new_n550), .A4(new_n571), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n552), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G475), .A2(G902), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n551), .B1(new_n572), .B2(KEYINPUT91), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n575), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n578), .B1(new_n581), .B2(KEYINPUT20), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT20), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n576), .A2(new_n579), .A3(new_n583), .A4(new_n577), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n554), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n199), .B2(G143), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n199), .A2(G143), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n265), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n588), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT95), .B1(new_n592), .B2(new_n586), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(G128), .B(G143), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n276), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G122), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G116), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n302), .A2(G122), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n388), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n276), .B(new_n595), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n388), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n598), .B1(new_n599), .B2(KEYINPUT14), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n599), .A2(KEYINPUT14), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT96), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n599), .A2(new_n608), .A3(KEYINPUT14), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n603), .B(new_n604), .C1(new_n388), .C2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n382), .A2(new_n187), .A3(G953), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n602), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n602), .B2(new_n611), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OR3_X1    g429(.A1(new_n615), .A2(KEYINPUT97), .A3(G902), .ZN(new_n616));
  INV_X1    g430(.A(G478), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(KEYINPUT15), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n188), .B1(new_n613), .B2(new_n614), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT97), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n616), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n619), .A2(new_n618), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n191), .A2(G952), .ZN(new_n624));
  INV_X1    g438(.A(G234), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n522), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n188), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT21), .B(G898), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n585), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n381), .A2(new_n473), .A3(new_n515), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  INV_X1    g448(.A(new_n379), .ZN(new_n635));
  INV_X1    g449(.A(G472), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n372), .B2(new_n188), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n635), .A2(new_n637), .A3(new_n258), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n473), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT98), .Z(new_n640));
  INV_X1    g454(.A(new_n630), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n515), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n615), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(G478), .A3(new_n188), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n642), .A2(new_n585), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n385), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n553), .A2(new_n188), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(G475), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n576), .A2(new_n583), .A3(new_n577), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n583), .B1(new_n576), .B2(new_n577), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n656), .B(new_n623), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n654), .B1(new_n660), .B2(new_n630), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n578), .A2(KEYINPUT20), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n554), .B1(new_n662), .B2(new_n657), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n663), .A2(KEYINPUT100), .A3(new_n641), .A4(new_n623), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n661), .A2(new_n515), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n640), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT35), .B(G107), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  AOI21_X1  g483(.A(KEYINPUT25), .B1(new_n254), .B2(new_n188), .ZN(new_n670));
  INV_X1    g484(.A(new_n243), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n189), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n673));
  INV_X1    g487(.A(new_n255), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n237), .B(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT36), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n195), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n678), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n674), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n672), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT103), .B1(new_n244), .B2(new_n681), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n585), .A2(new_n683), .A3(new_n631), .A4(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n635), .A2(new_n637), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n473), .A2(new_n515), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  NAND2_X1  g503(.A1(new_n372), .A2(new_n374), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n355), .A2(G472), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n380), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n683), .A2(new_n515), .A3(new_n684), .ZN(new_n693));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n627), .B1(new_n628), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n660), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n473), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  XOR2_X1   g514(.A(new_n695), .B(KEYINPUT39), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n473), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n703));
  INV_X1    g517(.A(new_n514), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n511), .B1(new_n500), .B2(new_n509), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT38), .Z(new_n707));
  OAI21_X1  g521(.A(new_n353), .B1(new_n325), .B2(new_n326), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT104), .Z(new_n709));
  OAI21_X1  g523(.A(new_n188), .B1(new_n709), .B2(new_n370), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G472), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n380), .A3(new_n690), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n582), .A2(new_n584), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n656), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n623), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n244), .A2(new_n681), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n474), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n713), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n703), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G143), .ZN(G45));
  NOR3_X1   g536(.A1(new_n585), .A2(new_n648), .A3(new_n695), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n692), .A2(new_n723), .A3(new_n693), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n466), .A2(new_n472), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n383), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT105), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n683), .A2(new_n684), .A3(new_n515), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n380), .B2(new_n375), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n473), .A4(new_n723), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT106), .B(G146), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G48));
  INV_X1    g548(.A(new_n462), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n461), .B1(new_n458), .B2(new_n447), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n446), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n737), .A2(new_n455), .B1(new_n451), .B2(new_n464), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(G902), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n383), .A3(new_n472), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n381), .A3(new_n649), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND3_X1  g557(.A1(new_n665), .A2(new_n740), .A3(new_n381), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NAND4_X1  g559(.A1(new_n739), .A2(new_n383), .A3(new_n472), .A4(new_n515), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n692), .A3(new_n685), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  NOR3_X1   g563(.A1(new_n716), .A2(new_n475), .A3(new_n706), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n376), .B(KEYINPUT107), .Z(new_n751));
  NAND2_X1  g565(.A1(new_n372), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n637), .A3(new_n258), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n740), .A3(new_n641), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  NAND2_X1  g570(.A1(new_n372), .A2(new_n188), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n757), .A2(G472), .B1(new_n372), .B2(new_n751), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n648), .B1(new_n714), .B2(new_n656), .ZN(new_n759));
  INV_X1    g573(.A(new_n717), .ZN(new_n760));
  INV_X1    g574(.A(new_n695), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n746), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n212), .ZN(G27));
  NAND3_X1  g578(.A1(new_n706), .A2(new_n383), .A3(new_n474), .ZN(new_n765));
  NAND2_X1  g579(.A1(G469), .A2(G902), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT108), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n465), .B2(G469), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n769), .B2(new_n472), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n381), .A2(new_n770), .A3(new_n723), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT109), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n381), .A2(new_n770), .A3(new_n774), .A4(new_n723), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n771), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT110), .B1(new_n777), .B2(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n772), .A2(KEYINPUT110), .A3(new_n773), .A4(new_n775), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n278), .ZN(G33));
  NAND3_X1  g596(.A1(new_n381), .A2(new_n770), .A3(new_n696), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n585), .A2(new_n647), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT111), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT43), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n686), .A2(new_n717), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n706), .A2(new_n474), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT112), .Z(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n465), .A2(KEYINPUT45), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n471), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n465), .A2(KEYINPUT45), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n768), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT46), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n472), .B1(new_n798), .B2(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n383), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n701), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT47), .B(new_n383), .C1(new_n799), .C2(new_n800), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n692), .A2(new_n257), .A3(new_n792), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n723), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT113), .B(G140), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G42));
  INV_X1    g627(.A(new_n740), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n792), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n712), .A2(new_n626), .A3(new_n258), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n585), .A3(new_n648), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n757), .A2(G472), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n760), .A3(new_n752), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n815), .A2(new_n627), .A3(new_n787), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n824));
  OR3_X1    g638(.A1(new_n814), .A2(new_n474), .A3(new_n707), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n787), .A2(new_n627), .A3(new_n754), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n787), .A2(new_n627), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n814), .A2(new_n474), .A3(new_n707), .ZN(new_n829));
  NOR2_X1   g643(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n828), .A2(new_n754), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n823), .A2(KEYINPUT118), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n822), .A2(new_n821), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n831), .A3(new_n827), .A4(new_n817), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n826), .A2(new_n793), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n739), .A2(new_n472), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(new_n384), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n809), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n832), .A2(new_n836), .A3(new_n840), .A4(KEYINPUT51), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n815), .A2(new_n759), .A3(new_n816), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n842), .B(new_n624), .C1(new_n826), .C2(new_n746), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n822), .A2(new_n381), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n834), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT51), .B1(new_n849), .B2(new_n840), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n744), .A2(new_n633), .A3(new_n687), .A4(new_n741), .ZN(new_n852));
  INV_X1    g666(.A(new_n759), .ZN(new_n853));
  INV_X1    g667(.A(new_n623), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n715), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n642), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n473), .A3(new_n856), .A4(new_n638), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n755), .A2(new_n748), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n821), .A2(new_n723), .A3(new_n770), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n783), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n663), .A2(new_n854), .A3(new_n761), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n683), .A2(new_n684), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(new_n792), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n473), .A3(new_n692), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(KEYINPUT114), .A3(new_n473), .A4(new_n692), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n779), .A2(new_n859), .A3(new_n780), .A4(new_n869), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n697), .A2(new_n726), .B1(new_n762), .B2(new_n746), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n769), .A2(new_n472), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n760), .A2(new_n384), .A3(new_n695), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT115), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n712), .A3(new_n750), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n732), .A2(new_n872), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n871), .B1(new_n731), .B2(new_n727), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(KEYINPUT52), .A3(new_n879), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n870), .A2(KEYINPUT53), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n859), .A2(new_n869), .A3(new_n779), .A4(new_n780), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT52), .B1(new_n883), .B2(new_n879), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND4_X1   g704(.A1(KEYINPUT52), .A2(new_n732), .A3(new_n872), .A4(new_n879), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n882), .A2(new_n891), .A3(KEYINPUT116), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n887), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n886), .B1(new_n893), .B2(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n891), .B1(KEYINPUT116), .B2(new_n882), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n880), .A2(new_n889), .A3(new_n881), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n870), .B(KEYINPUT53), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  INV_X1    g713(.A(new_n885), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n887), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n898), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n851), .A2(new_n895), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(G952), .B2(G953), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n838), .B(KEYINPUT49), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n712), .A2(new_n258), .ZN(new_n907));
  NOR4_X1   g721(.A1(new_n707), .A2(new_n384), .A3(new_n475), .A4(new_n785), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(G75));
  NOR2_X1   g724(.A1(new_n191), .A2(G952), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n504), .A2(new_n506), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n508), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n188), .B1(new_n898), .B2(new_n901), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G210), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(KEYINPUT119), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n914), .A2(KEYINPUT120), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n916), .B(new_n919), .C1(KEYINPUT119), .C2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n911), .B1(new_n921), .B2(new_n923), .ZN(G51));
  AND3_X1   g738(.A1(new_n898), .A2(new_n902), .A3(new_n901), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n902), .B1(new_n898), .B2(new_n901), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n767), .B(KEYINPUT57), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n470), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n915), .A2(new_n797), .A3(new_n796), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n911), .B1(new_n929), .B2(new_n930), .ZN(G54));
  AND2_X1   g745(.A1(KEYINPUT58), .A2(G475), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n915), .A2(new_n576), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n576), .B1(new_n915), .B2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n911), .ZN(G60));
  INV_X1    g749(.A(new_n911), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n644), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n936), .B1(new_n927), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n938), .B1(new_n895), .B2(new_n903), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n644), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n870), .B1(new_n896), .B2(new_n897), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n899), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n902), .B1(new_n946), .B2(new_n886), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n939), .B1(new_n947), .B2(new_n925), .ZN(new_n948));
  INV_X1    g762(.A(new_n644), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(KEYINPUT121), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n941), .B1(new_n944), .B2(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(new_n898), .A2(new_n901), .ZN(new_n952));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT122), .Z(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT60), .Z(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n254), .B(KEYINPUT123), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n911), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  INV_X1    g773(.A(new_n955), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n898), .B2(new_n901), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n679), .A2(new_n680), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n958), .A2(KEYINPUT124), .A3(new_n959), .A4(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n966));
  INV_X1    g780(.A(new_n957), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n936), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n952), .A2(new_n962), .A3(new_n955), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n965), .B(new_n966), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n964), .A2(new_n970), .ZN(G66));
  INV_X1    g785(.A(new_n859), .ZN(new_n972));
  NAND2_X1  g786(.A1(G224), .A2(G953), .ZN(new_n973));
  OAI22_X1  g787(.A1(new_n972), .A2(G953), .B1(new_n629), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n912), .B1(G898), .B2(new_n191), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n974), .B(new_n975), .Z(G69));
  NAND2_X1  g790(.A1(new_n368), .A2(new_n343), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n564), .A2(new_n558), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(G900), .A2(G953), .ZN(new_n980));
  INV_X1    g794(.A(new_n781), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n883), .A2(new_n783), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n750), .A2(new_n381), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n803), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n804), .A2(new_n981), .A3(new_n811), .A4(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n979), .B(new_n980), .C1(new_n985), .C2(G953), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n883), .A2(new_n721), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT62), .Z(new_n988));
  INV_X1    g802(.A(new_n702), .ZN(new_n989));
  INV_X1    g803(.A(new_n792), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(new_n381), .A3(new_n990), .A4(new_n855), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n804), .A2(new_n811), .ZN(new_n993));
  AOI21_X1  g807(.A(G953), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n986), .B1(new_n994), .B2(new_n979), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n986), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g813(.A(new_n986), .B1(new_n997), .B2(new_n996), .C1(new_n994), .C2(new_n979), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(new_n349), .A2(new_n324), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n332), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n992), .A2(new_n859), .A3(new_n993), .ZN(new_n1004));
  XOR2_X1   g818(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1005));
  NOR2_X1   g819(.A1(new_n636), .A2(new_n188), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n985), .B2(new_n972), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n349), .A2(new_n324), .A3(new_n353), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT127), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AND4_X1   g826(.A1(new_n894), .A2(new_n1010), .A3(new_n1003), .A4(new_n1007), .ZN(new_n1013));
  NOR4_X1   g827(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .A4(new_n911), .ZN(G57));
endmodule


