//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT94), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT94), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT14), .A3(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(KEYINPUT14), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT15), .A4(new_n211), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n203), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n203), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G1gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT95), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(G1gat), .B2(new_n221), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n219), .A2(new_n227), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT13), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT96), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT96), .ZN(new_n235));
  AOI211_X1 g034(.A(new_n235), .B(new_n232), .C1(new_n228), .C2(new_n229), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OR3_X1    g036(.A1(new_n216), .A2(KEYINPUT17), .A3(new_n218), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT17), .B1(new_n216), .B2(new_n218), .ZN(new_n239));
  INV_X1    g038(.A(new_n227), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n231), .A3(new_n229), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n229), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT93), .B1(new_n237), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT11), .ZN(new_n250));
  INV_X1    g049(.A(G169gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT92), .B(KEYINPUT12), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(KEYINPUT93), .B(new_n254), .C1(new_n237), .C2(new_n246), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n259));
  XNOR2_X1  g058(.A(G183gat), .B(G211gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G71gat), .A2(G78gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT98), .ZN(new_n264));
  NAND2_X1  g063(.A1(G71gat), .A2(G78gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT97), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G64gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT99), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT100), .Z(new_n271));
  AOI21_X1  g070(.A(new_n267), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(G71gat), .A2(G78gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n268), .B1(new_n273), .B2(new_n265), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT21), .ZN(new_n278));
  INV_X1    g077(.A(G127gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n227), .B1(KEYINPUT21), .B2(new_n277), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT101), .B(G155gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n282), .A2(new_n285), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n262), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n288), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(new_n286), .A3(new_n261), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G99gat), .A2(G106gat), .ZN(new_n293));
  INV_X1    g092(.A(G85gat), .ZN(new_n294));
  INV_X1    g093(.A(G92gat), .ZN(new_n295));
  AOI22_X1  g094(.A1(KEYINPUT8), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n294), .B2(new_n295), .ZN(new_n298));
  NAND4_X1  g097(.A1(KEYINPUT102), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G99gat), .B(G106gat), .Z(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n238), .A2(new_n239), .A3(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n300), .A2(new_n301), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n300), .A2(new_n301), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n219), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n307), .A2(KEYINPUT103), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT103), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G190gat), .B(G218gat), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n313), .ZN(new_n315));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT105), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT105), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n314), .A2(new_n321), .A3(new_n315), .A4(new_n318), .ZN(new_n322));
  INV_X1    g121(.A(new_n314), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT104), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT104), .B1(new_n311), .B2(new_n313), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n318), .B1(new_n314), .B2(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n320), .A2(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n292), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n251), .A2(new_n329), .A3(KEYINPUT23), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(G169gat), .B2(G176gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT65), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT66), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G190gat), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n338), .A2(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n334), .B(new_n336), .C1(new_n345), .C2(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n353), .A2(KEYINPUT25), .A3(new_n333), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n349), .A2(KEYINPUT25), .B1(new_n354), .B2(new_n335), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT67), .B(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT27), .B(G183gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT28), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT27), .ZN(new_n360));
  NOR2_X1   g159(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n356), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n363), .B2(KEYINPUT28), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n251), .A2(new_n329), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT26), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n335), .B1(new_n365), .B2(KEYINPUT26), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n346), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n279), .A2(G134gat), .ZN(new_n373));
  INV_X1    g172(.A(G134gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G127gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT68), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n279), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G113gat), .B(G120gat), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n377), .B(new_n378), .C1(KEYINPUT1), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G120gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G113gat), .ZN(new_n382));
  INV_X1    g181(.A(G113gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G120gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT69), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G127gat), .B(G134gat), .ZN(new_n387));
  AND2_X1   g186(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n388));
  NOR2_X1   g187(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n381), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n386), .A2(new_n387), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n380), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n380), .A2(new_n392), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n355), .A2(new_n395), .A3(new_n371), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT34), .ZN(new_n398));
  AND2_X1   g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT64), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n394), .B2(new_n396), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n398), .ZN(new_n403));
  INV_X1    g202(.A(new_n400), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n394), .A2(new_n396), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT32), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n402), .A2(new_n398), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n406), .A3(new_n401), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n412), .A2(KEYINPUT71), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(KEYINPUT71), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n405), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(G15gat), .B(G43gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT72), .ZN(new_n417));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n408), .A2(new_n410), .A3(new_n415), .A4(new_n419), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT36), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT36), .B1(new_n421), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n349), .A2(KEYINPUT25), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n354), .A2(new_n335), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT66), .B(G183gat), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n361), .B1(new_n431), .B2(KEYINPUT27), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n432), .B2(new_n356), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n369), .B1(new_n433), .B2(new_n359), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n426), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n355), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT29), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT76), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n355), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT75), .B1(new_n355), .B2(new_n371), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT76), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n438), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n372), .A2(new_n439), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G211gat), .B(G218gat), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G197gat), .B(G204gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(G211gat), .A2(G218gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT22), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT74), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n454), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(new_n449), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n457), .B(KEYINPUT73), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n450), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n448), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n435), .A2(new_n439), .A3(new_n436), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n372), .A2(new_n441), .A3(new_n438), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n467), .B2(new_n461), .ZN(new_n468));
  AOI211_X1 g267(.A(KEYINPUT77), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G8gat), .B(G36gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT78), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n473), .B(G64gat), .Z(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(new_n295), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n475), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n463), .A2(new_n477), .A3(new_n470), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n479));
  OR3_X1    g278(.A1(new_n471), .A2(KEYINPUT30), .A3(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT0), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(G57gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(new_n294), .ZN(new_n485));
  XNOR2_X1  g284(.A(G141gat), .B(G148gat), .ZN(new_n486));
  INV_X1    g285(.A(G162gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT80), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G162gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(G155gat), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n486), .B1(new_n491), .B2(KEYINPUT2), .ZN(new_n492));
  XNOR2_X1  g291(.A(G155gat), .B(G162gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G148gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G141gat), .ZN(new_n496));
  INV_X1    g295(.A(G141gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G148gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n500));
  INV_X1    g299(.A(G155gat), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n487), .ZN(new_n502));
  NAND2_X1  g301(.A1(G155gat), .A2(G162gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT79), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n494), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n395), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n493), .A2(new_n492), .B1(new_n502), .B2(new_n504), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n508), .A2(new_n393), .A3(KEYINPUT82), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT82), .B1(new_n508), .B2(new_n393), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G225gat), .A2(G233gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n515));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n509), .B2(new_n510), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT3), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n508), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n506), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n508), .A2(new_n519), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n395), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n393), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n512), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n514), .B(new_n515), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  OR3_X1    g326(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n516), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n515), .A2(new_n513), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n528), .A2(new_n523), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n485), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT6), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n527), .A2(new_n485), .A3(new_n531), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(new_n532), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT84), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n527), .A2(new_n531), .ZN(new_n538));
  INV_X1    g337(.A(new_n485), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n527), .A2(new_n485), .A3(new_n531), .ZN(new_n541));
  AND4_X1   g340(.A1(KEYINPUT84), .A2(new_n540), .A3(new_n536), .A4(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n533), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n481), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n508), .A2(KEYINPUT29), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n461), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n506), .A2(KEYINPUT3), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT86), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT29), .B1(new_n508), .B2(new_n519), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(new_n461), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(KEYINPUT86), .A3(new_n547), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G228gat), .ZN(new_n555));
  INV_X1    g354(.A(G233gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n457), .A2(new_n449), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n459), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n441), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n508), .B1(new_n561), .B2(new_n519), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n551), .A2(new_n461), .B1(new_n555), .B2(new_n556), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G50gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G78gat), .B(G106gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT85), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n558), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n571), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n558), .B2(new_n565), .ZN(new_n576));
  AOI211_X1 g375(.A(new_n567), .B(new_n564), .C1(new_n554), .C2(new_n557), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n574), .A2(new_n578), .A3(KEYINPUT87), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT87), .B1(new_n574), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n425), .B1(new_n544), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n463), .A2(new_n583), .A3(new_n470), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n448), .A2(new_n461), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n467), .A2(new_n462), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT37), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n584), .A2(new_n587), .A3(new_n588), .A4(new_n475), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT90), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n475), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n583), .B1(new_n463), .B2(new_n470), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT38), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n540), .A2(new_n536), .A3(new_n541), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n594), .A2(new_n478), .A3(new_n533), .ZN(new_n595));
  INV_X1    g394(.A(new_n586), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n448), .B2(new_n461), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT38), .B1(new_n597), .B2(KEYINPUT37), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n598), .A2(new_n599), .A3(new_n475), .A4(new_n584), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n590), .A2(new_n593), .A3(new_n595), .A4(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n574), .A2(new_n578), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n511), .A2(new_n513), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT89), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT89), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n528), .A2(new_n523), .A3(new_n529), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n606), .B2(new_n513), .ZN(new_n607));
  OAI211_X1 g406(.A(KEYINPUT39), .B(new_n604), .C1(new_n607), .C2(new_n603), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n606), .A2(new_n513), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n539), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT40), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n532), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n611), .A3(KEYINPUT40), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n613), .A2(new_n479), .A3(new_n480), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n601), .A2(new_n602), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n582), .A2(new_n616), .ZN(new_n617));
  AND4_X1   g416(.A1(new_n574), .A2(new_n578), .A3(new_n421), .A4(new_n422), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n481), .A2(new_n543), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT35), .ZN(new_n620));
  AND2_X1   g419(.A1(KEYINPUT91), .A2(KEYINPUT35), .ZN(new_n621));
  NOR2_X1   g420(.A1(KEYINPUT91), .A2(KEYINPUT35), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n621), .B(new_n622), .C1(new_n594), .C2(new_n533), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n481), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n258), .B(new_n328), .C1(new_n617), .C2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n269), .A2(new_n271), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n306), .B(new_n275), .C1(new_n627), .C2(new_n267), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n302), .B1(new_n272), .B2(new_n276), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n329), .ZN(new_n635));
  INV_X1    g434(.A(G204gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n628), .A2(new_n639), .A3(new_n629), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n277), .A2(KEYINPUT10), .A3(new_n306), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n632), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI211_X1 g443(.A(KEYINPUT106), .B(new_n632), .C1(new_n640), .C2(new_n641), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n633), .B(new_n638), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n642), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n633), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n637), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n626), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n543), .B(KEYINPUT107), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  INV_X1    g456(.A(new_n481), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n222), .A2(new_n220), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR4_X1   g463(.A1(new_n659), .A2(KEYINPUT42), .A3(new_n660), .A4(new_n661), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT108), .B1(new_n659), .B2(G8gat), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n659), .A2(KEYINPUT108), .A3(G8gat), .ZN(new_n667));
  OAI22_X1  g466(.A1(new_n664), .A2(new_n665), .B1(new_n666), .B2(new_n667), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n425), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n652), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n421), .A2(new_n422), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n653), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n671), .B1(new_n669), .B2(new_n674), .ZN(G1326gat));
  INV_X1    g474(.A(new_n581), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  AOI21_X1  g478(.A(new_n327), .B1(new_n617), .B2(new_n625), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n258), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n292), .A2(new_n650), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n685), .A2(KEYINPUT110), .A3(new_n654), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT110), .B1(new_n685), .B2(new_n654), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(G29gat), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n258), .B1(new_n617), .B2(new_n625), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n292), .A2(new_n327), .A3(new_n650), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n205), .A3(new_n655), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n688), .A2(new_n696), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n693), .A2(G36gat), .A3(new_n481), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n685), .B2(new_n481), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  OAI21_X1  g500(.A(G43gat), .B1(new_n685), .B2(new_n670), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n693), .A2(G43gat), .A3(new_n672), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1330gat));
  OAI21_X1  g507(.A(G50gat), .B1(new_n685), .B2(new_n602), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n676), .B1(new_n694), .B2(KEYINPUT111), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711));
  AOI21_X1  g510(.A(G50gat), .B1(new_n693), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n709), .A2(KEYINPUT48), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n682), .A2(new_n581), .A3(new_n683), .A4(new_n684), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n715), .A2(G50gat), .B1(new_n710), .B2(new_n712), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g516(.A(new_n651), .B1(new_n617), .B2(new_n625), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n328), .A2(new_n683), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n655), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g522(.A(new_n481), .B(KEYINPUT112), .Z(new_n724));
  NOR2_X1   g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  AOI21_X1  g528(.A(G71gat), .B1(new_n721), .B2(new_n673), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n425), .A2(G71gat), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g532(.A1(new_n721), .A2(new_n581), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n292), .A2(new_n683), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n651), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n682), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n654), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT114), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n327), .B(new_n737), .C1(new_n617), .C2(new_n625), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(KEYINPUT51), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n680), .A2(new_n736), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(KEYINPUT114), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n617), .A2(new_n625), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n320), .A2(new_n322), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n324), .A2(new_n326), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n751), .A4(new_n736), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT113), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n680), .A2(new_n754), .A3(KEYINPUT51), .A4(new_n736), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n650), .B1(new_n747), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n655), .A2(new_n294), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n740), .B1(new_n757), .B2(new_n758), .ZN(G1336gat));
  AND2_X1   g558(.A1(new_n682), .A2(new_n738), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n295), .B1(new_n760), .B2(new_n658), .ZN(new_n761));
  INV_X1    g560(.A(new_n724), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n295), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n651), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n742), .A2(KEYINPUT51), .ZN(new_n765));
  INV_X1    g564(.A(new_n752), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT115), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G92gat), .B1(new_n739), .B2(new_n724), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n774));
  OAI211_X1 g573(.A(new_n773), .B(new_n774), .C1(new_n757), .C2(new_n763), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n739), .B2(new_n670), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n672), .A2(G99gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n757), .B2(new_n778), .ZN(G1338gat));
  INV_X1    g578(.A(G106gat), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n760), .B2(new_n581), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n602), .A2(G106gat), .A3(new_n651), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT53), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n783), .B1(new_n747), .B2(new_n756), .ZN(new_n787));
  INV_X1    g586(.A(new_n602), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n681), .B1(new_n748), .B2(new_n751), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT44), .B(new_n327), .C1(new_n617), .C2(new_n625), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n788), .B(new_n738), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT53), .B1(new_n791), .B2(G106gat), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT117), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n743), .A2(new_n746), .B1(new_n753), .B2(new_n755), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(KEYINPUT117), .C1(new_n794), .C2(new_n784), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n786), .B1(new_n793), .B2(new_n796), .ZN(G1339gat));
  NOR2_X1   g596(.A1(new_n230), .A2(new_n233), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT119), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n231), .B1(new_n241), .B2(new_n229), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n252), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n237), .A2(new_n246), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n254), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n803), .A3(new_n650), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n640), .A2(new_n641), .A3(new_n632), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT54), .B(new_n805), .C1(new_n644), .C2(new_n645), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n638), .B1(new_n642), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT118), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n805), .A2(KEYINPUT54), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n647), .A2(KEYINPUT106), .ZN(new_n813));
  INV_X1    g612(.A(new_n645), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n808), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n811), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n806), .A2(new_n818), .A3(new_n808), .A4(KEYINPUT55), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n810), .A2(new_n646), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n804), .B1(new_n820), .B2(new_n258), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n327), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n810), .A2(new_n646), .A3(new_n819), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n801), .A2(new_n803), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n751), .A2(new_n823), .A3(new_n824), .A4(new_n817), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n292), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n328), .A2(new_n650), .A3(new_n683), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n655), .A3(new_n724), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n581), .A3(new_n672), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n258), .ZN(new_n832));
  INV_X1    g631(.A(new_n618), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n383), .A3(new_n683), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(G1340gat));
  OAI21_X1  g635(.A(G120gat), .B1(new_n831), .B2(new_n651), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n381), .A3(new_n650), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1341gat));
  AOI21_X1  g638(.A(G127gat), .B1(new_n834), .B2(new_n292), .ZN(new_n840));
  INV_X1    g639(.A(new_n292), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n279), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n830), .B2(new_n842), .ZN(G1342gat));
  OAI21_X1  g642(.A(G134gat), .B1(new_n831), .B2(new_n327), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n828), .A2(new_n655), .A3(new_n481), .A4(new_n751), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(G134gat), .A3(new_n833), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n847), .B2(new_n845), .ZN(new_n850));
  OAI221_X1 g649(.A(new_n844), .B1(new_n845), .B2(new_n847), .C1(new_n849), .C2(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n828), .A2(new_n852), .A3(new_n788), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n762), .A2(new_n654), .A3(new_n425), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n815), .B2(new_n816), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n810), .A2(new_n646), .A3(new_n819), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n804), .B1(new_n857), .B2(new_n258), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n327), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n292), .B1(new_n859), .B2(new_n825), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n827), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n676), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n853), .B(new_n854), .C1(new_n864), .C2(new_n852), .ZN(new_n865));
  OAI21_X1  g664(.A(G141gat), .B1(new_n865), .B2(new_n258), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n829), .A2(new_n602), .A3(new_n425), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n258), .A2(G141gat), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n867), .A2(new_n868), .B1(KEYINPUT123), .B2(KEYINPUT58), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n870), .B(new_n872), .ZN(G1344gat));
  NAND3_X1  g672(.A1(new_n867), .A2(new_n495), .A3(new_n650), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n581), .B1(new_n860), .B2(new_n827), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n852), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT124), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n828), .A2(KEYINPUT57), .A3(new_n788), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n880), .A3(new_n852), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n650), .A3(new_n854), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n875), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n875), .B(G148gat), .C1(new_n865), .C2(new_n651), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n874), .B1(new_n884), .B2(new_n886), .ZN(G1345gat));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n292), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n501), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n292), .A2(G155gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n865), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n889), .B(new_n893), .C1(new_n865), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1346gat));
  NOR2_X1   g694(.A1(new_n865), .A2(new_n327), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n488), .A2(new_n490), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n425), .A2(new_n602), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n897), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n896), .A2(new_n897), .B1(new_n846), .B2(new_n899), .ZN(G1347gat));
  AND2_X1   g699(.A1(new_n828), .A2(new_n654), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n901), .A2(new_n618), .A3(new_n762), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n251), .A3(new_n683), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n901), .A2(new_n658), .A3(new_n676), .A4(new_n673), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n258), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n902), .B2(new_n650), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n904), .A2(new_n329), .A3(new_n651), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  NAND3_X1  g708(.A1(new_n902), .A2(new_n358), .A3(new_n292), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n431), .B1(new_n904), .B2(new_n841), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n902), .A2(new_n357), .A3(new_n751), .ZN(new_n914));
  OAI21_X1  g713(.A(G190gat), .B1(new_n904), .B2(new_n327), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n655), .A2(new_n481), .A3(new_n425), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n882), .A2(new_n683), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G197gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n762), .A3(new_n898), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n922), .A2(G197gat), .A3(new_n258), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n921), .A2(new_n926), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1352gat));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n901), .A2(new_n636), .A3(new_n762), .A4(new_n898), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT127), .B1(new_n930), .B2(new_n651), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n930), .A2(KEYINPUT127), .A3(new_n651), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n933), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(KEYINPUT62), .A3(new_n931), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n882), .A2(new_n650), .A3(new_n919), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(G1353gat));
  OR3_X1    g738(.A1(new_n922), .A2(G211gat), .A3(new_n841), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n882), .A2(new_n292), .A3(new_n919), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1354gat));
  NOR2_X1   g743(.A1(new_n922), .A2(new_n327), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(G218gat), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n882), .A2(new_n919), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n751), .A2(G218gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(G1355gat));
endmodule


