

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n976), .A2(n701), .ZN(n704) );
  BUF_X1 U549 ( .A(n725), .Z(n737) );
  NAND2_X1 U550 ( .A1(n878), .A2(G137), .ZN(n532) );
  INV_X1 U551 ( .A(KEYINPUT29), .ZN(n718) );
  NAND2_X1 U552 ( .A1(n736), .A2(n735), .ZN(n748) );
  NAND2_X1 U553 ( .A1(n691), .A2(n690), .ZN(n725) );
  INV_X1 U554 ( .A(KEYINPUT17), .ZN(n530) );
  NOR2_X1 U555 ( .A1(G651), .A2(n621), .ZN(n641) );
  NOR2_X1 U556 ( .A1(n535), .A2(n534), .ZN(n537) );
  NOR2_X2 U557 ( .A1(n541), .A2(n540), .ZN(G160) );
  XNOR2_X1 U558 ( .A(KEYINPUT78), .B(KEYINPUT7), .ZN(n529) );
  NOR2_X1 U559 ( .A1(G543), .A2(G651), .ZN(n513) );
  XNOR2_X1 U560 ( .A(n513), .B(KEYINPUT64), .ZN(n642) );
  NAND2_X1 U561 ( .A1(G89), .A2(n642), .ZN(n514) );
  XNOR2_X1 U562 ( .A(n514), .B(KEYINPUT4), .ZN(n516) );
  XOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .Z(n621) );
  XNOR2_X1 U564 ( .A(G651), .B(KEYINPUT67), .ZN(n519) );
  NOR2_X1 U565 ( .A1(n621), .A2(n519), .ZN(n639) );
  NAND2_X1 U566 ( .A1(G76), .A2(n639), .ZN(n515) );
  NAND2_X1 U567 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U568 ( .A(n517), .B(KEYINPUT5), .ZN(n527) );
  XNOR2_X1 U569 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n641), .A2(G51), .ZN(n518) );
  XNOR2_X1 U571 ( .A(n518), .B(KEYINPUT76), .ZN(n523) );
  NOR2_X1 U572 ( .A1(G543), .A2(n519), .ZN(n520) );
  XOR2_X1 U573 ( .A(KEYINPUT68), .B(n520), .Z(n521) );
  XNOR2_X1 U574 ( .A(KEYINPUT1), .B(n521), .ZN(n645) );
  NAND2_X1 U575 ( .A1(G63), .A2(n645), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U577 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n529), .B(n528), .ZN(G168) );
  XOR2_X1 U580 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  XNOR2_X2 U582 ( .A(n531), .B(n530), .ZN(n878) );
  XOR2_X1 U583 ( .A(n532), .B(KEYINPUT66), .Z(n535) );
  INV_X1 U584 ( .A(G2105), .ZN(n538) );
  AND2_X1 U585 ( .A1(n538), .A2(G2104), .ZN(n879) );
  NAND2_X1 U586 ( .A1(G101), .A2(n879), .ZN(n533) );
  XNOR2_X1 U587 ( .A(KEYINPUT23), .B(n533), .ZN(n534) );
  AND2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n874) );
  NAND2_X1 U589 ( .A1(n874), .A2(G113), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n541) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n538), .ZN(n875) );
  NAND2_X1 U592 ( .A1(G125), .A2(n875), .ZN(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT65), .B(n539), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n641), .A2(G52), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G64), .A2(n645), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U597 ( .A1(G77), .A2(n639), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G90), .A2(n642), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U600 ( .A(KEYINPUT9), .B(n546), .ZN(n547) );
  XNOR2_X1 U601 ( .A(KEYINPUT69), .B(n547), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(G171) );
  XOR2_X1 U603 ( .A(KEYINPUT109), .B(G2435), .Z(n551) );
  XNOR2_X1 U604 ( .A(G2430), .B(G2438), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n551), .B(n550), .ZN(n558) );
  XOR2_X1 U606 ( .A(G2446), .B(G2454), .Z(n553) );
  XNOR2_X1 U607 ( .A(G2451), .B(G2443), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U609 ( .A(n554), .B(G2427), .Z(n556) );
  XNOR2_X1 U610 ( .A(G1348), .B(G1341), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U612 ( .A(n558), .B(n557), .ZN(n559) );
  AND2_X1 U613 ( .A1(n559), .A2(G14), .ZN(G401) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  NAND2_X1 U617 ( .A1(n641), .A2(G53), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G65), .A2(n645), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G78), .A2(n639), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G91), .A2(n642), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n713) );
  INV_X1 U624 ( .A(n713), .ZN(G299) );
  NAND2_X1 U625 ( .A1(G94), .A2(G452), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT70), .B(n566), .Z(G173) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n832) );
  NAND2_X1 U630 ( .A1(n832), .A2(G567), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n645), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n569), .Z(n577) );
  NAND2_X1 U634 ( .A1(G68), .A2(n639), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT71), .B(KEYINPUT12), .Z(n571) );
  NAND2_X1 U636 ( .A1(G81), .A2(n642), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT13), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(n575), .Z(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n641), .A2(G43), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n976) );
  INV_X1 U644 ( .A(G860), .ZN(n595) );
  OR2_X1 U645 ( .A1(n976), .A2(n595), .ZN(G153) );
  XNOR2_X1 U646 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT74), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G54), .A2(n641), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n639), .A2(G79), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G66), .A2(n645), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G92), .A2(n642), .ZN(n583) );
  XNOR2_X1 U654 ( .A(KEYINPUT75), .B(n583), .ZN(n584) );
  NOR2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U657 ( .A(n588), .B(KEYINPUT15), .ZN(n963) );
  OR2_X1 U658 ( .A1(G868), .A2(n963), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(G284) );
  INV_X1 U660 ( .A(G868), .ZN(n591) );
  NOR2_X1 U661 ( .A1(G286), .A2(n591), .ZN(n592) );
  XOR2_X1 U662 ( .A(KEYINPUT79), .B(n592), .Z(n594) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n596), .A2(n963), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT16), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n598) );
  XNOR2_X1 U669 ( .A(n599), .B(n598), .ZN(G148) );
  NOR2_X1 U670 ( .A1(G868), .A2(n976), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n963), .A2(G868), .ZN(n600) );
  NOR2_X1 U672 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U674 ( .A1(G123), .A2(n875), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n879), .A2(G99), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G111), .A2(n874), .ZN(n607) );
  NAND2_X1 U679 ( .A1(G135), .A2(n878), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n911) );
  XNOR2_X1 U682 ( .A(n911), .B(G2096), .ZN(n611) );
  INV_X1 U683 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U685 ( .A1(n963), .A2(G559), .ZN(n661) );
  XNOR2_X1 U686 ( .A(n976), .B(n661), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n612), .A2(G860), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n641), .A2(G55), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G93), .A2(n642), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G80), .A2(n639), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT82), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G67), .A2(n645), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n654) );
  XNOR2_X1 U696 ( .A(n620), .B(n654), .ZN(G145) );
  NAND2_X1 U697 ( .A1(G87), .A2(n621), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n645), .A2(n624), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n641), .A2(G49), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U703 ( .A1(G75), .A2(n639), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G88), .A2(n642), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n641), .A2(G50), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G62), .A2(n645), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(G166) );
  AND2_X1 U710 ( .A1(G60), .A2(n645), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G72), .A2(n639), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G47), .A2(n641), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G85), .A2(n642), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G73), .A2(n639), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n641), .A2(G48), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G86), .A2(n642), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G61), .A2(n645), .ZN(n646) );
  XNOR2_X1 U723 ( .A(KEYINPUT83), .B(n646), .ZN(n647) );
  NOR2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(G305) );
  NOR2_X1 U726 ( .A1(G868), .A2(n654), .ZN(n651) );
  XOR2_X1 U727 ( .A(n651), .B(KEYINPUT86), .Z(n664) );
  XNOR2_X1 U728 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n653) );
  XNOR2_X1 U729 ( .A(G288), .B(KEYINPUT19), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(n658) );
  XNOR2_X1 U731 ( .A(G166), .B(n654), .ZN(n656) );
  XNOR2_X1 U732 ( .A(G290), .B(n713), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(G305), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n976), .B(n660), .ZN(n901) );
  XOR2_X1 U737 ( .A(n901), .B(n661), .Z(n662) );
  NAND2_X1 U738 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(G295) );
  INV_X1 U740 ( .A(G2072), .ZN(n922) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XOR2_X1 U744 ( .A(KEYINPUT21), .B(n667), .Z(n668) );
  NOR2_X1 U745 ( .A1(n922), .A2(n668), .ZN(n669) );
  XNOR2_X1 U746 ( .A(KEYINPUT87), .B(n669), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U750 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U751 ( .A1(G96), .A2(n672), .ZN(n836) );
  NAND2_X1 U752 ( .A1(G2106), .A2(n836), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n673), .B(KEYINPUT88), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U755 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G108), .A2(n675), .ZN(n837) );
  NAND2_X1 U757 ( .A1(G567), .A2(n837), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U759 ( .A(KEYINPUT89), .B(n678), .ZN(G319) );
  INV_X1 U760 ( .A(G319), .ZN(n680) );
  NAND2_X1 U761 ( .A1(G661), .A2(G483), .ZN(n679) );
  NOR2_X1 U762 ( .A1(n680), .A2(n679), .ZN(n835) );
  NAND2_X1 U763 ( .A1(n835), .A2(G36), .ZN(n681) );
  XNOR2_X1 U764 ( .A(KEYINPUT90), .B(n681), .ZN(G176) );
  NAND2_X1 U765 ( .A1(n878), .A2(G138), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G114), .A2(n874), .ZN(n682) );
  XOR2_X1 U767 ( .A(KEYINPUT91), .B(n682), .Z(n683) );
  NAND2_X1 U768 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U769 ( .A1(G102), .A2(n879), .ZN(n686) );
  NAND2_X1 U770 ( .A1(G126), .A2(n875), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U772 ( .A1(n688), .A2(n687), .ZN(G164) );
  XOR2_X1 U773 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  XNOR2_X1 U774 ( .A(G1986), .B(G290), .ZN(n968) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n690) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n690), .A2(n689), .ZN(n827) );
  NAND2_X1 U778 ( .A1(n968), .A2(n827), .ZN(n814) );
  INV_X1 U779 ( .A(n689), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n725), .A2(n922), .ZN(n693) );
  XNOR2_X1 U781 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U782 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U783 ( .A1(n737), .A2(G1956), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U785 ( .A(KEYINPUT99), .B(n696), .ZN(n712) );
  NOR2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n697) );
  XOR2_X1 U787 ( .A(n697), .B(KEYINPUT28), .Z(n717) );
  INV_X1 U788 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U789 ( .A1(n725), .A2(n942), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n698), .B(KEYINPUT26), .ZN(n700) );
  AND2_X1 U791 ( .A1(n725), .A2(G1341), .ZN(n699) );
  OR2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U793 ( .A1(n704), .A2(n963), .ZN(n703) );
  INV_X1 U794 ( .A(KEYINPUT100), .ZN(n702) );
  XNOR2_X1 U795 ( .A(n703), .B(n702), .ZN(n711) );
  NAND2_X1 U796 ( .A1(n704), .A2(n963), .ZN(n709) );
  INV_X1 U797 ( .A(n737), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n705), .A2(G1348), .ZN(n707) );
  NOR2_X1 U799 ( .A1(G2067), .A2(n737), .ZN(n706) );
  NOR2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U806 ( .A(n719), .B(n718), .ZN(n723) );
  XNOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .ZN(n941) );
  NOR2_X1 U808 ( .A1(n737), .A2(n941), .ZN(n721) );
  AND2_X1 U809 ( .A1(n737), .A2(G1961), .ZN(n720) );
  NOR2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U811 ( .A1(G171), .A2(n724), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n736) );
  INV_X1 U813 ( .A(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U814 ( .A1(G171), .A2(n724), .ZN(n732) );
  INV_X1 U815 ( .A(KEYINPUT101), .ZN(n727) );
  NAND2_X1 U816 ( .A1(G8), .A2(n725), .ZN(n778) );
  NOR2_X1 U817 ( .A1(G1966), .A2(n778), .ZN(n750) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n737), .ZN(n747) );
  NOR2_X1 U819 ( .A1(n750), .A2(n747), .ZN(n726) );
  XNOR2_X1 U820 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U821 ( .A1(G8), .A2(n728), .ZN(n729) );
  XNOR2_X1 U822 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n730), .A2(G168), .ZN(n731) );
  NOR2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U825 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n748), .A2(G286), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n778), .ZN(n739) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n737), .ZN(n738) );
  NOR2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U830 ( .A1(n740), .A2(G303), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U832 ( .A(n743), .B(KEYINPUT102), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n744), .A2(G8), .ZN(n746) );
  XOR2_X1 U834 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n745) );
  XNOR2_X1 U835 ( .A(n746), .B(n745), .ZN(n770) );
  NAND2_X1 U836 ( .A1(G8), .A2(n747), .ZN(n752) );
  INV_X1 U837 ( .A(n748), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n771) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G288), .A2(G1976), .ZN(n753) );
  XOR2_X1 U842 ( .A(KEYINPUT105), .B(n753), .Z(n970) );
  AND2_X1 U843 ( .A1(n754), .A2(n970), .ZN(n756) );
  AND2_X1 U844 ( .A1(n771), .A2(n756), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n770), .A2(n755), .ZN(n767) );
  INV_X1 U846 ( .A(n778), .ZN(n761) );
  INV_X1 U847 ( .A(n756), .ZN(n759) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n762) );
  NOR2_X1 U849 ( .A1(G303), .A2(G1971), .ZN(n757) );
  OR2_X1 U850 ( .A1(n762), .A2(n757), .ZN(n972) );
  XOR2_X1 U851 ( .A(KEYINPUT104), .B(n972), .Z(n758) );
  OR2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n760) );
  OR2_X1 U853 ( .A1(n778), .A2(n760), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U855 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  AND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U858 ( .A(n768), .B(KEYINPUT106), .ZN(n769) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n960) );
  NAND2_X1 U860 ( .A1(n769), .A2(n960), .ZN(n782) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n774) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  AND2_X1 U865 ( .A1(n775), .A2(n778), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U867 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n812) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G140), .A2(n878), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G104), .A2(n879), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n786), .B(n785), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G116), .A2(n874), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G128), .A2(n875), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U881 ( .A(KEYINPUT36), .B(n792), .Z(n897) );
  XOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .Z(n793) );
  XOR2_X1 U883 ( .A(KEYINPUT93), .B(n793), .Z(n823) );
  AND2_X1 U884 ( .A1(n897), .A2(n823), .ZN(n918) );
  NAND2_X1 U885 ( .A1(n827), .A2(n918), .ZN(n821) );
  XOR2_X1 U886 ( .A(KEYINPUT97), .B(KEYINPUT38), .Z(n795) );
  NAND2_X1 U887 ( .A1(G105), .A2(n879), .ZN(n794) );
  XNOR2_X1 U888 ( .A(n795), .B(n794), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G141), .A2(n878), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G129), .A2(n875), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n874), .A2(G117), .ZN(n798) );
  XOR2_X1 U893 ( .A(KEYINPUT96), .B(n798), .Z(n799) );
  NOR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n890) );
  AND2_X1 U896 ( .A1(n890), .A2(G1996), .ZN(n912) );
  NAND2_X1 U897 ( .A1(G131), .A2(n878), .ZN(n804) );
  NAND2_X1 U898 ( .A1(G119), .A2(n875), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G95), .A2(n879), .ZN(n805) );
  XNOR2_X1 U901 ( .A(KEYINPUT95), .B(n805), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n874), .A2(G107), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n889) );
  AND2_X1 U905 ( .A1(n889), .A2(G1991), .ZN(n914) );
  OR2_X1 U906 ( .A1(n912), .A2(n914), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n810), .A2(n827), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n821), .A2(n815), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n830) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n890), .ZN(n928) );
  INV_X1 U912 ( .A(n815), .ZN(n818) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n889), .ZN(n913) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n913), .A2(n816), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n928), .A2(n819), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n823), .A2(n897), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n824), .B(KEYINPUT107), .ZN(n934) );
  NAND2_X1 U922 ( .A1(n825), .A2(n934), .ZN(n826) );
  XNOR2_X1 U923 ( .A(KEYINPUT108), .B(n826), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n831), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U929 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U939 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U941 ( .A(KEYINPUT110), .B(G2090), .Z(n841) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U944 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U947 ( .A(G2078), .B(G2084), .Z(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(G227) );
  XNOR2_X1 U949 ( .A(G1976), .B(G2474), .ZN(n857) );
  XOR2_X1 U950 ( .A(G1971), .B(G1956), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1961), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U953 ( .A(G1981), .B(G1966), .Z(n851) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U955 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U956 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U957 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G124), .A2(n875), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n879), .A2(G100), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G112), .A2(n874), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G136), .A2(n878), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G139), .A2(n878), .ZN(n866) );
  NAND2_X1 U969 ( .A1(G103), .A2(n879), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n875), .A2(G127), .ZN(n867) );
  XNOR2_X1 U972 ( .A(KEYINPUT113), .B(n867), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n874), .A2(G115), .ZN(n868) );
  XOR2_X1 U974 ( .A(KEYINPUT114), .B(n868), .Z(n869) );
  NOR2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U976 ( .A(n871), .B(KEYINPUT47), .ZN(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n921) );
  NAND2_X1 U978 ( .A1(G118), .A2(n874), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G130), .A2(n875), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G142), .A2(n878), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G106), .A2(n879), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n882), .Z(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n921), .B(n885), .ZN(n896) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n887) );
  XNOR2_X1 U988 ( .A(n911), .B(KEYINPUT115), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U990 ( .A(G160), .B(n888), .ZN(n894) );
  XNOR2_X1 U991 ( .A(G162), .B(n889), .ZN(n892) );
  XOR2_X1 U992 ( .A(G164), .B(n890), .Z(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(n900) );
  XNOR2_X1 U998 ( .A(KEYINPUT116), .B(n900), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n963), .B(G286), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n903), .B(G171), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n904), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT49), .B(n905), .Z(n906) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n906), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n907), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n908) );
  XOR2_X1 U1008 ( .A(KEYINPUT117), .B(n908), .Z(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(G160), .B(G2084), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n933) );
  XNOR2_X1 U1018 ( .A(n921), .B(KEYINPUT118), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n923), .B(n922), .ZN(n925) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n926), .ZN(n931) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n929), .Z(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n936), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n937), .A2(G29), .ZN(n1017) );
  XOR2_X1 U1031 ( .A(G25), .B(G1991), .Z(n938) );
  NAND2_X1 U1032 ( .A1(n938), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(G2072), .B(G33), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n946) );
  XOR2_X1 U1036 ( .A(n941), .B(G27), .Z(n944) );
  XOR2_X1 U1037 ( .A(n942), .B(G32), .Z(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1041 ( .A(KEYINPUT53), .B(n949), .Z(n953) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n950), .B(G34), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G2084), .B(n951), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(G35), .B(G2090), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n956), .B(KEYINPUT120), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(G29), .A2(n957), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(KEYINPUT55), .B(n958), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n959), .A2(G11), .ZN(n1015) );
  XNOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .ZN(n985) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G168), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(KEYINPUT57), .B(n962), .ZN(n983) );
  XNOR2_X1 U1056 ( .A(G1348), .B(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G171), .B(G1961), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT121), .B(n966), .ZN(n980) );
  XNOR2_X1 U1060 ( .A(G1956), .B(G299), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n975) );
  NAND2_X1 U1062 ( .A1(G303), .A2(G1971), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n973), .B(KEYINPUT122), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G1341), .B(n976), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(KEYINPUT123), .B(n981), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n1013) );
  INV_X1 U1073 ( .A(G16), .ZN(n1011) );
  XOR2_X1 U1074 ( .A(G1986), .B(G24), .Z(n989) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G23), .B(G1976), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(n991), .B(n990), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G21), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G5), .B(G1961), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n1008) );
  XOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .Z(n996) );
  XNOR2_X1 U1086 ( .A(G4), .B(n996), .ZN(n1004) );
  XOR2_X1 U1087 ( .A(G1981), .B(G6), .Z(n999) );
  XOR2_X1 U1088 ( .A(G20), .B(KEYINPUT124), .Z(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(G1956), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(G19), .B(G1341), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT125), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT126), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

