//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT75), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT75), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(G146), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n192), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G128), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G119), .B(G128), .ZN(new_n207));
  INV_X1    g021(.A(G110), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT24), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n206), .A2(G110), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n195), .A2(new_n199), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT76), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n195), .A2(new_n213), .A3(new_n216), .A4(new_n199), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT77), .ZN(new_n219));
  OR3_X1    g033(.A1(new_n206), .A2(new_n219), .A3(G110), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n206), .B2(G110), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n212), .A2(new_n207), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT65), .B(G146), .ZN(new_n224));
  XNOR2_X1  g038(.A(G125), .B(G140), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n218), .A2(KEYINPUT78), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT78), .B1(new_n218), .B2(new_n228), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G137), .ZN(new_n231));
  INV_X1    g045(.A(G953), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(G221), .A3(G234), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n231), .B(new_n233), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n229), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n218), .A2(new_n228), .A3(new_n234), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT25), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G217), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(G234), .B2(new_n237), .ZN(new_n241));
  INV_X1    g055(.A(new_n230), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n218), .A2(KEYINPUT78), .A3(new_n228), .ZN(new_n243));
  INV_X1    g057(.A(new_n234), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n246));
  INV_X1    g060(.A(new_n238), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n241), .A3(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n245), .A2(new_n236), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n241), .A2(G902), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT2), .A2(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT2), .A2(G113), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT2), .A3(G113), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G116), .B(G119), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n201), .A2(G116), .ZN(new_n262));
  INV_X1    g076(.A(G116), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G119), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n261), .B1(new_n269), .B2(new_n259), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(KEYINPUT64), .A2(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT64), .A2(G143), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(G146), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n196), .A2(KEYINPUT65), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G146), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n278), .A3(G143), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n272), .A2(new_n275), .A3(new_n279), .A4(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(G146), .B1(new_n273), .B2(new_n274), .ZN(new_n281));
  AOI21_X1  g095(.A(G143), .B1(new_n276), .B2(new_n278), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n204), .B1(new_n279), .B2(new_n271), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G134), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G137), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(G137), .ZN(new_n289));
  OAI21_X1  g103(.A(G131), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT11), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n286), .B2(G137), .ZN(new_n292));
  INV_X1    g106(.A(G137), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT11), .A3(G134), .ZN(new_n294));
  INV_X1    g108(.A(G131), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n292), .A2(new_n294), .A3(new_n295), .A4(new_n287), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n292), .A2(new_n294), .A3(new_n287), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G131), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n296), .ZN(new_n301));
  AND2_X1   g115(.A1(KEYINPUT0), .A2(G128), .ZN(new_n302));
  NOR2_X1   g116(.A1(KEYINPUT0), .A2(G128), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n281), .B2(new_n282), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n275), .A2(new_n279), .A3(new_n302), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n298), .A2(KEYINPUT30), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n301), .A2(KEYINPUT66), .A3(new_n305), .A4(new_n306), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n310), .A2(new_n311), .B1(new_n285), .B2(new_n297), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n270), .B(new_n308), .C1(new_n312), .C2(KEYINPUT30), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT26), .B(G101), .ZN(new_n314));
  INV_X1    g128(.A(G237), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n232), .A3(G210), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n314), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n270), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n298), .A2(new_n320), .A3(new_n307), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n313), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT31), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n313), .A2(KEYINPUT31), .A3(new_n319), .A4(new_n321), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n321), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(KEYINPUT28), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT71), .B1(new_n312), .B2(new_n320), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n275), .A2(new_n279), .ZN(new_n330));
  AND2_X1   g144(.A1(KEYINPUT64), .A2(G143), .ZN(new_n331));
  NOR2_X1   g145(.A1(KEYINPUT64), .A2(G143), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n196), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n224), .B2(G143), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n330), .A2(new_n302), .B1(new_n334), .B2(new_n304), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT66), .B1(new_n335), .B2(new_n301), .ZN(new_n336));
  INV_X1    g150(.A(new_n311), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n298), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n270), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n329), .A2(new_n340), .A3(new_n321), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n328), .B1(new_n341), .B2(KEYINPUT28), .ZN(new_n342));
  OAI22_X1  g156(.A1(new_n324), .A2(new_n326), .B1(new_n342), .B2(new_n319), .ZN(new_n343));
  NOR2_X1   g157(.A1(G472), .A2(G902), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT32), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(KEYINPUT28), .ZN(new_n346));
  INV_X1    g160(.A(new_n328), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n319), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n322), .A2(new_n323), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n325), .ZN(new_n351));
  INV_X1    g165(.A(new_n344), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT74), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n310), .A2(new_n311), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n320), .B1(new_n358), .B2(new_n298), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n327), .B1(new_n359), .B2(new_n339), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n360), .B2(new_n329), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n349), .B1(new_n361), .B2(new_n328), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n350), .A2(new_n325), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT74), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n345), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n320), .B1(new_n298), .B2(new_n307), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n327), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n370), .B2(KEYINPUT28), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n368), .B(KEYINPUT28), .C1(new_n327), .C2(new_n369), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n347), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n319), .A2(KEYINPUT29), .ZN(new_n375));
  AOI21_X1  g189(.A(G902), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n342), .A2(KEYINPUT72), .A3(new_n319), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n313), .A2(new_n321), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n378), .B2(new_n349), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT72), .B1(new_n342), .B2(new_n319), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G472), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n253), .B1(new_n367), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n315), .A2(new_n232), .A3(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n273), .A2(new_n274), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(new_n385), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G131), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n195), .A2(new_n199), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n388), .B(G131), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(KEYINPUT17), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT89), .B(G104), .Z(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n226), .B1(new_n196), .B2(new_n225), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT18), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n295), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n388), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n390), .B2(KEYINPUT18), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n394), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n225), .B(KEYINPUT19), .Z(new_n405));
  INV_X1    g219(.A(new_n224), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n227), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n393), .B2(KEYINPUT88), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n388), .A2(G131), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n390), .A2(new_n409), .A3(KEYINPUT88), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n402), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n404), .B1(new_n411), .B2(new_n397), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  NOR2_X1   g227(.A1(G475), .A2(G902), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT90), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n412), .A2(new_n417), .A3(new_n413), .A4(new_n414), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n414), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT20), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n404), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n397), .B1(new_n394), .B2(new_n403), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n237), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G475), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n331), .A2(new_n332), .A3(new_n204), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT92), .A3(KEYINPUT13), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n204), .A2(G143), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(KEYINPUT13), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n273), .A2(G128), .A3(new_n274), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT13), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(G134), .B(new_n428), .C1(new_n430), .C2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n286), .A3(new_n429), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n436), .A2(KEYINPUT93), .ZN(new_n437));
  INV_X1    g251(.A(G107), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n263), .A2(G122), .ZN(new_n439));
  INV_X1    g253(.A(G122), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G116), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT91), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT91), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n440), .A2(G116), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n263), .A2(G122), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT91), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(G107), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n436), .A2(KEYINPUT93), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n435), .A2(new_n437), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT95), .ZN(new_n454));
  AOI21_X1  g268(.A(G107), .B1(new_n448), .B2(new_n449), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n286), .B1(new_n432), .B2(new_n429), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n455), .B1(new_n457), .B2(new_n436), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n446), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n439), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n447), .B1(new_n460), .B2(new_n446), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n438), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n454), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n436), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n444), .B1(new_n468), .B2(new_n456), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n469), .A2(KEYINPUT95), .A3(new_n465), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n453), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT9), .B(G234), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT79), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n240), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n474), .B(new_n453), .C1(new_n467), .C2(new_n470), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(KEYINPUT96), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT96), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n479), .A3(new_n475), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n237), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT97), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n478), .A2(KEYINPUT97), .A3(new_n237), .A4(new_n480), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G478), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT98), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n481), .B2(new_n482), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n487), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n483), .B2(new_n484), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT98), .B1(new_n494), .B2(new_n490), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n426), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT80), .Z(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT82), .B(G104), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT83), .B1(new_n500), .B2(G107), .ZN(new_n501));
  INV_X1    g315(.A(G104), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT82), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G104), .ZN(new_n505));
  AND4_X1   g319(.A1(KEYINPUT83), .A2(new_n503), .A3(new_n505), .A4(G107), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT3), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n438), .A3(G104), .ZN(new_n509));
  AOI21_X1  g323(.A(G107), .B1(new_n503), .B2(new_n505), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g325(.A(G101), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n503), .A2(new_n505), .A3(G107), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT83), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n500), .A2(KEYINPUT83), .A3(G107), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G101), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT3), .B1(new_n500), .B2(G107), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n509), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(G101), .C1(new_n507), .C2(new_n511), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n335), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n301), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n438), .A2(G104), .ZN(new_n526));
  OAI21_X1  g340(.A(G101), .B1(new_n510), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n204), .B1(new_n333), .B2(KEYINPUT1), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n280), .B1(new_n330), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n520), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT10), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n520), .A2(new_n285), .A3(KEYINPUT10), .A4(new_n527), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n524), .A2(new_n525), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n525), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n520), .A2(new_n527), .A3(new_n529), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n285), .B1(new_n520), .B2(new_n527), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n535), .A2(new_n536), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G110), .B(G140), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT81), .ZN(new_n544));
  INV_X1    g358(.A(G227), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n544), .B(new_n546), .Z(new_n547));
  OAI221_X1 g361(.A(new_n537), .B1(new_n535), .B2(new_n536), .C1(new_n538), .C2(new_n539), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n534), .A2(new_n542), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n521), .A2(new_n335), .A3(new_n523), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n532), .A2(new_n533), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n301), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n547), .B1(new_n552), .B2(new_n534), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI211_X1 g369(.A(KEYINPUT85), .B(new_n547), .C1(new_n552), .C2(new_n534), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n499), .B(new_n237), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n534), .A2(new_n542), .A3(new_n548), .ZN(new_n558));
  INV_X1    g372(.A(new_n547), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(new_n547), .A3(new_n534), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(G469), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n499), .A2(new_n237), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n498), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G214), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G210), .B1(G237), .B2(G902), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n521), .A2(new_n270), .A3(new_n523), .ZN(new_n570));
  INV_X1    g384(.A(new_n261), .ZN(new_n571));
  OAI21_X1  g385(.A(G113), .B1(new_n262), .B2(KEYINPUT5), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n269), .B2(KEYINPUT5), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT5), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n266), .B2(new_n268), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT86), .B1(new_n577), .B2(new_n572), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n575), .A2(new_n520), .A3(new_n527), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G122), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n570), .A2(new_n579), .A3(new_n581), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n586), .A3(new_n582), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n285), .A2(new_n189), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n305), .A2(G125), .A3(new_n306), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G224), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(G953), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n585), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n588), .A2(new_n589), .B1(KEYINPUT87), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n592), .A2(new_n595), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n265), .A2(new_n576), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n261), .B1(new_n572), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n520), .A2(new_n527), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n581), .B(KEYINPUT8), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n573), .A2(new_n574), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n578), .A3(new_n261), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n520), .A2(new_n527), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n602), .B(new_n603), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  OAI221_X1 g421(.A(new_n597), .B1(KEYINPUT87), .B2(new_n595), .C1(new_n588), .C2(new_n589), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n599), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n609), .B2(new_n584), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n569), .B1(new_n594), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n594), .A2(new_n610), .A3(new_n569), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n568), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(G234), .A2(G237), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(G952), .A3(new_n232), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT99), .Z(new_n617));
  AND3_X1   g431(.A1(new_n615), .A2(G902), .A3(G953), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT21), .B(G898), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n566), .A2(new_n614), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n384), .A2(new_n496), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n478), .A2(new_n627), .A3(new_n480), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n476), .A2(KEYINPUT33), .A3(new_n477), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(G478), .A3(new_n237), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n481), .A2(new_n486), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n426), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n594), .A2(new_n610), .A3(new_n569), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n622), .B(new_n567), .C1(new_n634), .C2(new_n611), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n626), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n421), .A2(new_n425), .B1(new_n631), .B2(new_n630), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n614), .A2(new_n637), .A3(KEYINPUT101), .A4(new_n622), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(G902), .B1(new_n362), .B2(new_n363), .ZN(new_n640));
  NAND2_X1  g454(.A1(KEYINPUT100), .A2(G472), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n642), .A2(new_n643), .A3(new_n253), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n639), .A2(new_n566), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n420), .A2(new_n415), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(new_n425), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n492), .A2(new_n495), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n623), .A3(new_n644), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n642), .A2(new_n643), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n242), .B(new_n243), .C1(KEYINPUT36), .C2(new_n244), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n244), .A2(KEYINPUT36), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n658), .B1(new_n229), .B2(new_n230), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n251), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n249), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n656), .B1(new_n249), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n623), .A2(new_n496), .A3(new_n655), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT103), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  OAI21_X1  g481(.A(new_n567), .B1(new_n634), .B2(new_n611), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n662), .A3(new_n661), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n353), .B1(new_n351), .B2(new_n352), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n365), .B1(new_n343), .B2(new_n354), .ZN(new_n671));
  AOI211_X1 g485(.A(KEYINPUT74), .B(new_n355), .C1(new_n362), .C2(new_n363), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(G472), .ZN(new_n674));
  INV_X1    g488(.A(new_n381), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n377), .A3(new_n379), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n674), .B1(new_n676), .B2(new_n376), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n669), .B(new_n566), .C1(new_n673), .C2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n618), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n617), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n492), .A2(new_n495), .A3(new_n649), .A4(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT104), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n683), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n663), .A2(new_n566), .A3(new_n614), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n367), .A2(new_n383), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n685), .A2(new_n687), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  NAND2_X1  g506(.A1(new_n492), .A2(new_n495), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n421), .A2(new_n425), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n634), .A2(new_n611), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n567), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n681), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n566), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n249), .A2(new_n660), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n237), .B1(new_n370), .B2(new_n319), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n349), .B1(new_n313), .B2(new_n321), .ZN(new_n705));
  OAI21_X1  g519(.A(G472), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n670), .B(new_n706), .C1(new_n671), .C2(new_n672), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n699), .A2(new_n702), .A3(new_n703), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(new_n387), .Z(G45));
  AOI21_X1  g524(.A(new_n686), .B1(new_n383), .B2(new_n367), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n633), .A2(new_n681), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  INV_X1    g529(.A(new_n639), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n237), .B1(new_n555), .B2(new_n556), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G469), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n718), .A2(new_n497), .A3(new_n557), .ZN(new_n719));
  INV_X1    g533(.A(new_n253), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n719), .B(new_n720), .C1(new_n673), .C2(new_n677), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n715), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n639), .A2(new_n384), .A3(KEYINPUT106), .A4(new_n719), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  INV_X1    g540(.A(new_n635), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n384), .A2(new_n727), .A3(new_n651), .A4(new_n719), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NAND2_X1  g543(.A1(new_n718), .A2(new_n557), .ZN(new_n730));
  INV_X1    g544(.A(new_n497), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n730), .A2(new_n668), .A3(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n661), .A2(new_n662), .A3(new_n621), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n689), .A2(new_n732), .A3(new_n733), .A4(new_n496), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  AND4_X1   g549(.A1(new_n426), .A2(new_n492), .A3(new_n614), .A4(new_n495), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n349), .B1(new_n371), .B2(new_n373), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n363), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n344), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n720), .B(new_n739), .C1(new_n640), .C2(new_n674), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n730), .A2(new_n621), .A3(new_n731), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n736), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND2_X1  g558(.A1(new_n719), .A2(new_n614), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n739), .B(new_n703), .C1(new_n640), .C2(new_n674), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n712), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n189), .ZN(G27));
  INV_X1    g564(.A(new_n712), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n561), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n552), .A2(KEYINPUT107), .A3(new_n547), .A4(new_n534), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n560), .A4(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n564), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n557), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n634), .A2(new_n611), .A3(new_n568), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n497), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n751), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n345), .B2(new_n364), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n343), .A2(new_n354), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n352), .B1(new_n362), .B2(new_n363), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n763), .B(new_n764), .C1(KEYINPUT32), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n383), .A3(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n767), .A2(KEYINPUT109), .A3(new_n720), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT109), .B1(new_n767), .B2(new_n720), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n761), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(new_n761), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n720), .B1(new_n673), .B2(new_n677), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n759), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n712), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n771), .A2(new_n773), .B1(new_n760), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n295), .ZN(G33));
  NOR3_X1   g592(.A1(new_n774), .A2(new_n683), .A3(new_n759), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n286), .ZN(G36));
  NAND2_X1  g594(.A1(new_n694), .A2(KEYINPUT111), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n426), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n632), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n426), .A2(KEYINPUT43), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n784), .A2(KEYINPUT43), .B1(new_n632), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n703), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n655), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n758), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n786), .A2(new_n788), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n790), .B1(KEYINPUT44), .B2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(KEYINPUT45), .A2(new_n753), .A3(new_n560), .A4(new_n754), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT45), .B1(new_n560), .B2(new_n561), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(new_n499), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(new_n563), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n557), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n796), .A2(new_n797), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n497), .A3(new_n700), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT112), .B(G137), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G39));
  OAI21_X1  g619(.A(new_n497), .B1(new_n799), .B2(new_n800), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT47), .B(new_n497), .C1(new_n799), .C2(new_n800), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n673), .A2(new_n677), .ZN(new_n811));
  INV_X1    g625(.A(new_n758), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n751), .A2(new_n812), .A3(new_n720), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  INV_X1    g629(.A(new_n498), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n720), .A2(new_n567), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n698), .A2(new_n784), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n730), .B(KEYINPUT49), .Z(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n708), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n617), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n786), .A2(new_n821), .A3(new_n741), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n812), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n730), .A2(new_n816), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n823), .B1(new_n810), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n698), .A2(new_n567), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n719), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n822), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n826), .B1(new_n822), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n786), .A2(new_n821), .A3(new_n719), .A4(new_n758), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n746), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n719), .A2(new_n758), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n834), .A2(new_n253), .A3(new_n707), .A4(new_n617), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n426), .A2(new_n632), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n825), .A2(KEYINPUT51), .A3(new_n831), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n767), .A2(new_n720), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT109), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n767), .A2(KEYINPUT109), .A3(new_n720), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n832), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT48), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n232), .A2(G952), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT119), .Z(new_n846));
  NOR2_X1   g660(.A1(new_n822), .A2(new_n745), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n846), .B(new_n847), .C1(new_n637), .C2(new_n835), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n838), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n776), .A2(new_n760), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n841), .A2(new_n842), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n772), .B1(new_n851), .B2(new_n761), .ZN(new_n852));
  INV_X1    g666(.A(new_n773), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n488), .A2(new_n855), .A3(new_n491), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT113), .B1(new_n494), .B2(new_n490), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n648), .A2(new_n425), .A3(new_n682), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n661), .A2(new_n859), .A3(new_n662), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n858), .A2(new_n860), .A3(new_n566), .A4(new_n758), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n861), .A2(new_n811), .B1(new_n748), .B2(new_n759), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n779), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n693), .A2(new_n694), .A3(new_n727), .A4(new_n566), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n655), .A2(new_n663), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n774), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n727), .A2(new_n495), .A3(new_n492), .A4(new_n649), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n721), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n856), .A2(new_n694), .A3(new_n857), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n633), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n644), .A3(new_n623), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n734), .A2(new_n872), .A3(new_n743), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n724), .A2(new_n863), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n682), .A2(new_n497), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n756), .B2(new_n557), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n707), .A2(new_n787), .A3(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n711), .A2(new_n712), .B1(new_n877), .B2(new_n736), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  INV_X1    g693(.A(new_n749), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n691), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n691), .A2(new_n880), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT52), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n854), .A2(new_n874), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT115), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n688), .B1(new_n711), .B2(new_n685), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n811), .A2(new_n683), .A3(new_n686), .A4(KEYINPUT104), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n880), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n749), .B1(new_n684), .B2(new_n690), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n877), .A2(new_n736), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n713), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT52), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n728), .A2(new_n624), .A3(new_n664), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n734), .A2(new_n872), .A3(new_n743), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n881), .A2(new_n724), .A3(new_n901), .A4(new_n863), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n777), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n898), .A2(new_n903), .A3(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n884), .A2(new_n905), .A3(new_n885), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n887), .A2(new_n888), .A3(new_n904), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n898), .B2(new_n903), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n884), .A2(new_n885), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT54), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n837), .A2(new_n831), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT117), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n837), .A2(new_n831), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n825), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(KEYINPUT116), .B(new_n823), .C1(new_n810), .C2(new_n824), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n912), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT118), .B(new_n912), .C1(new_n917), .C2(new_n921), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n849), .B(new_n911), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n820), .B1(new_n926), .B2(new_n927), .ZN(G75));
  NAND3_X1  g742(.A1(new_n887), .A2(new_n904), .A3(new_n906), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n585), .A2(new_n587), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n593), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT55), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n232), .A2(G952), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G51));
  NAND2_X1  g752(.A1(new_n904), .A2(new_n906), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n905), .B1(new_n884), .B2(new_n885), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT54), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n907), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n563), .B(KEYINPUT57), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n556), .B2(new_n555), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n929), .A2(G902), .A3(new_n795), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n937), .B1(new_n945), .B2(new_n948), .ZN(G54));
  INV_X1    g763(.A(new_n412), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n929), .A2(G902), .ZN(new_n951));
  NAND2_X1  g765(.A1(KEYINPUT58), .A2(G475), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n937), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n951), .A2(new_n950), .A3(new_n952), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(G60));
  XOR2_X1   g771(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n958));
  NOR2_X1   g772(.A1(new_n486), .A2(new_n237), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n628), .A2(new_n629), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n942), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n964), .A3(new_n954), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n911), .A2(new_n960), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n628), .A2(new_n629), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n941), .B2(new_n907), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT122), .B1(new_n969), .B2(new_n937), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n965), .A2(new_n968), .A3(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n929), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n250), .B(KEYINPUT123), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n929), .A2(new_n659), .A3(new_n657), .A4(new_n974), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n954), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n977), .A2(KEYINPUT61), .A3(new_n954), .A4(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n619), .B2(new_n591), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n901), .A2(new_n724), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n932), .B1(G898), .B2(new_n232), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  OAI21_X1  g803(.A(new_n308), .B1(new_n312), .B2(KEYINPUT30), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n405), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  OAI211_X1 g806(.A(G900), .B(G953), .C1(new_n992), .C2(new_n545), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n545), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n713), .B1(new_n893), .B2(new_n894), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT124), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT124), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n892), .A2(new_n998), .A3(new_n895), .A4(new_n713), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n803), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT125), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n802), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n736), .A3(new_n851), .ZN(new_n1004));
  INV_X1    g818(.A(new_n779), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1004), .A2(new_n814), .A3(new_n854), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1002), .A2(KEYINPUT126), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(KEYINPUT126), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n991), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n709), .B1(new_n997), .B2(new_n999), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT62), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n701), .A2(new_n812), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n384), .A2(new_n871), .A3(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n814), .B(new_n1016), .C1(new_n802), .C2(new_n792), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n991), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1011), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n994), .B1(new_n1021), .B2(new_n232), .ZN(G72));
  OR2_X1    g836(.A1(new_n908), .A2(new_n909), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n378), .A2(new_n319), .ZN(new_n1024));
  XNOR2_X1  g838(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n674), .A2(new_n237), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1025), .B(new_n1026), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1024), .A2(new_n705), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n937), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n985), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1028), .B1(new_n1018), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n705), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1010), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(new_n986), .A3(new_n1008), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n1027), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1034), .B1(new_n1037), .B2(new_n1024), .ZN(G57));
endmodule


