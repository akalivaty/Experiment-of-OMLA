//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT88), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(new_n191), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G953), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT68), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G953), .ZN(new_n203));
  INV_X1    g017(.A(G237), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n201), .A2(new_n203), .A3(G214), .A4(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT86), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT68), .B(G953), .ZN(new_n208));
  INV_X1    g022(.A(new_n206), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n208), .A2(G214), .A3(new_n204), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT18), .A2(G131), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n210), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT18), .A3(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT87), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n207), .B2(new_n210), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT87), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT18), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n213), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n207), .A2(new_n210), .A3(new_n217), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(new_n218), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n194), .A2(KEYINPUT19), .A3(new_n195), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n192), .A2(KEYINPUT19), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n197), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT16), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n188), .A3(G125), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n192), .B2(new_n228), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n230), .A2(new_n197), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n187), .B1(new_n221), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G113), .B(G122), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT90), .B(G104), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n235), .B(new_n236), .Z(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n199), .A2(new_n212), .ZN(new_n239));
  AND4_X1   g053(.A1(new_n219), .A2(new_n214), .A3(KEYINPUT18), .A4(G131), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n219), .B1(new_n218), .B2(KEYINPUT18), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n227), .B(new_n231), .C1(new_n223), .C2(new_n218), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(KEYINPUT89), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n234), .A2(new_n238), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n218), .A2(KEYINPUT17), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n230), .A2(new_n197), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n231), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n214), .A2(G131), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(new_n222), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT92), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n218), .A2(KEYINPUT17), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(KEYINPUT91), .A3(new_n248), .A4(new_n231), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT92), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n251), .A2(new_n257), .A3(new_n252), .A4(new_n222), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n250), .A2(new_n254), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n237), .A3(new_n242), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n245), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT93), .ZN(new_n262));
  NOR2_X1   g076(.A1(G475), .A2(G902), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n263), .B(KEYINPUT94), .Z(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT93), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n245), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n264), .A2(KEYINPUT20), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n268), .A2(KEYINPUT20), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n259), .A2(new_n242), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n238), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n260), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G475), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G116), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G122), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT95), .B1(new_n279), .B2(KEYINPUT14), .ZN(new_n280));
  INV_X1    g094(.A(G122), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G116), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT95), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT14), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n278), .A4(G122), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n279), .A2(KEYINPUT14), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n280), .A2(new_n282), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G107), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n282), .A2(new_n279), .ZN(new_n289));
  INV_X1    g103(.A(G107), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G128), .ZN(new_n293));
  INV_X1    g107(.A(G128), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G143), .ZN(new_n295));
  INV_X1    g109(.A(G134), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n293), .B2(new_n295), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n288), .B(new_n291), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n289), .B(new_n290), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT13), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n295), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n293), .A2(new_n302), .ZN(new_n305));
  OAI21_X1  g119(.A(G134), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n306), .A3(new_n297), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT72), .B(G217), .Z(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(G953), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n300), .A2(new_n307), .A3(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n274), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n316), .A2(KEYINPUT97), .ZN(new_n317));
  OAI21_X1  g131(.A(G478), .B1(KEYINPUT96), .B2(KEYINPUT15), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(KEYINPUT96), .B2(KEYINPUT15), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n316), .B(KEYINPUT97), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n274), .B(new_n208), .C1(G234), .C2(G237), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT21), .B(G898), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT98), .B(G952), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G953), .ZN(new_n327));
  INV_X1    g141(.A(G234), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(new_n204), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(new_n330), .B(KEYINPUT99), .Z(new_n331));
  AND2_X1   g145(.A1(new_n322), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G221), .B1(new_n310), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G469), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(new_n274), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n208), .A2(G227), .ZN(new_n337));
  XOR2_X1   g151(.A(G110), .B(G140), .Z(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G104), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(new_n340), .B2(G107), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n290), .A3(G104), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(G107), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G101), .ZN(new_n346));
  INV_X1    g160(.A(G101), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n341), .A2(new_n343), .A3(new_n347), .A4(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n346), .A2(KEYINPUT76), .A3(KEYINPUT4), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n197), .A2(G143), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n292), .A2(G146), .ZN(new_n355));
  AND2_X1   g169(.A1(KEYINPUT0), .A2(G128), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n292), .A2(G146), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT64), .B1(new_n197), .B2(G143), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT64), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n292), .A3(G146), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(KEYINPUT0), .A2(G128), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n358), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n345), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT77), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n345), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n367), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n353), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n340), .A2(G107), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n290), .A2(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(G101), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n348), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n294), .A2(KEYINPUT1), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n354), .A3(new_n355), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n294), .B1(new_n354), .B2(KEYINPUT1), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n354), .A2(new_n355), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n381), .A2(new_n382), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n379), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n381), .B1(new_n363), .B2(new_n384), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n378), .A2(new_n389), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n388), .A2(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT11), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n296), .B2(G137), .ZN(new_n394));
  INV_X1    g208(.A(G137), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT11), .A3(G134), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n296), .A2(G137), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G131), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n394), .A2(new_n396), .A3(new_n217), .A4(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n374), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n374), .B2(new_n392), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n339), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n374), .A2(new_n392), .A3(new_n402), .ZN(new_n406));
  INV_X1    g220(.A(new_n339), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n363), .A2(new_n384), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n381), .A3(new_n378), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n388), .A2(KEYINPUT79), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n379), .A2(new_n390), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n402), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT12), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT12), .B1(new_n410), .B2(new_n413), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n406), .B(new_n407), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n336), .B1(new_n417), .B2(new_n335), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n406), .B1(new_n414), .B2(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n339), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n406), .A2(new_n407), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n421), .A2(KEYINPUT80), .ZN(new_n422));
  INV_X1    g236(.A(new_n404), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n421), .B2(KEYINPUT80), .ZN(new_n424));
  OAI211_X1 g238(.A(G469), .B(new_n420), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n334), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n277), .A2(new_n332), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G472), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n274), .ZN(new_n429));
  INV_X1    g243(.A(G113), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT2), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G113), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n434), .A2(KEYINPUT66), .ZN(new_n435));
  XNOR2_X1  g249(.A(G116), .B(G119), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(KEYINPUT66), .B2(new_n434), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT67), .ZN(new_n438));
  INV_X1    g252(.A(G119), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G116), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n278), .A2(G119), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT2), .B(G113), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT67), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n435), .A2(new_n437), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n361), .B1(new_n292), .B2(G146), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n197), .A2(KEYINPUT64), .A3(G143), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n354), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n357), .B1(new_n450), .B2(new_n365), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n401), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n395), .A2(KEYINPUT65), .A3(G134), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n296), .B2(G137), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n395), .A2(G134), .ZN(new_n456));
  OAI211_X1 g270(.A(G131), .B(new_n453), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n457), .A2(new_n400), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n390), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n452), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n452), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n447), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n452), .A2(new_n459), .A3(new_n446), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT26), .B(G101), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n208), .A2(G210), .A3(new_n204), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT27), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT27), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n208), .A2(new_n468), .A3(G210), .A4(new_n204), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n469), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n464), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n463), .A2(KEYINPUT31), .A3(new_n464), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n464), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n452), .A2(new_n459), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n447), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n459), .A2(new_n452), .A3(new_n446), .A4(KEYINPUT28), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n471), .A2(KEYINPUT69), .A3(new_n472), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n429), .B1(new_n479), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(KEYINPUT71), .A3(new_n464), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n494), .A3(new_n447), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(KEYINPUT28), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n473), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n481), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n464), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n482), .A2(KEYINPUT30), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n452), .A2(new_n459), .A3(new_n460), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n500), .B1(new_n503), .B2(new_n447), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n474), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n497), .B1(new_n485), .B2(new_n489), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n499), .B(new_n274), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n492), .A2(KEYINPUT32), .B1(G472), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n490), .B1(new_n477), .B2(new_n478), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n429), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT70), .B(new_n509), .C1(new_n510), .C2(new_n429), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n294), .A2(G119), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n439), .A2(G128), .B1(KEYINPUT73), .B2(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(KEYINPUT73), .B2(KEYINPUT23), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT74), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n521), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n517), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(KEYINPUT23), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G110), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n439), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n532), .A3(new_n249), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n529), .A2(new_n531), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n523), .A2(new_n525), .ZN(new_n535));
  INV_X1    g349(.A(G110), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n231), .A2(new_n198), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n208), .A2(G221), .A3(G234), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT22), .B(G137), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n533), .B(new_n542), .C1(new_n537), .C2(new_n538), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n274), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT25), .A4(new_n274), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n309), .B1(G234), .B2(new_n274), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G902), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT75), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n544), .A2(new_n545), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n550), .A2(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n515), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G122), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n444), .A2(new_n445), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n435), .A2(new_n437), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n560), .A2(new_n561), .B1(new_n370), .B2(new_n372), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n353), .A2(new_n562), .A3(KEYINPUT81), .ZN(new_n563));
  OAI21_X1  g377(.A(G113), .B1(new_n440), .B2(KEYINPUT5), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(KEYINPUT5), .B2(new_n436), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n444), .B2(new_n445), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n379), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT81), .B1(new_n353), .B2(new_n562), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n559), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n353), .A2(new_n562), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT81), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(new_n558), .A3(new_n567), .A4(new_n563), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT82), .A4(KEYINPUT6), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n570), .A2(KEYINPUT6), .A3(new_n574), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n559), .C1(new_n568), .C2(new_n569), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT82), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n575), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n408), .A2(new_n190), .A3(new_n381), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n190), .B2(new_n451), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n200), .A2(G224), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT84), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n582), .B(KEYINPUT83), .C1(new_n190), .C2(new_n451), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(KEYINPUT7), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n589), .B(new_n590), .C1(KEYINPUT83), .C2(new_n582), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n558), .B(KEYINPUT8), .ZN(new_n592));
  INV_X1    g406(.A(new_n567), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n566), .A2(new_n379), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n583), .A2(new_n590), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n597), .B2(new_n574), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n587), .A2(new_n588), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n570), .A2(KEYINPUT6), .A3(new_n574), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n579), .A3(new_n578), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n585), .B1(new_n601), .B2(new_n575), .ZN(new_n602));
  INV_X1    g416(.A(new_n598), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT84), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G210), .B1(G237), .B2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n599), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n587), .A2(new_n605), .A3(new_n598), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G214), .B1(G237), .B2(G902), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT85), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT85), .ZN(new_n612));
  INV_X1    g426(.A(new_n610), .ZN(new_n613));
  AOI211_X1 g427(.A(new_n612), .B(new_n613), .C1(new_n607), .C2(new_n608), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n427), .B(new_n557), .C1(new_n611), .C2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n426), .A2(new_n555), .ZN(new_n618));
  INV_X1    g432(.A(new_n492), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n510), .B2(G902), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n617), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n621), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n623), .A2(KEYINPUT100), .A3(new_n555), .A4(new_n426), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n606), .B1(new_n602), .B2(new_n603), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n613), .B1(new_n608), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n300), .A2(new_n307), .A3(KEYINPUT103), .A4(new_n311), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n313), .A2(KEYINPUT33), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n314), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G478), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(G902), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT101), .B(KEYINPUT33), .Z(new_n636));
  AOI21_X1  g450(.A(new_n635), .B1(new_n315), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n636), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT102), .B(new_n638), .C1(new_n313), .C2(new_n314), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n632), .B(new_n634), .C1(new_n637), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT104), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n316), .A2(new_n633), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n640), .B2(KEYINPUT104), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n268), .A2(KEYINPUT20), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n261), .A2(new_n269), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n276), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n627), .A2(new_n650), .A3(new_n331), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n625), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT34), .B(G104), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  AND3_X1   g468(.A1(new_n245), .A2(new_n266), .A3(new_n260), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n266), .B1(new_n245), .B2(new_n260), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g471(.A1(KEYINPUT20), .A2(new_n268), .B1(new_n657), .B2(new_n269), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n658), .A2(new_n276), .A3(new_n322), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n627), .A2(new_n659), .A3(new_n331), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n625), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT35), .B(G107), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NAND2_X1  g477(.A1(new_n550), .A2(new_n551), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n543), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n539), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n553), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n621), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n427), .B(new_n670), .C1(new_n611), .C2(new_n614), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  AND3_X1   g487(.A1(new_n515), .A2(new_n426), .A3(new_n668), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n329), .B(KEYINPUT105), .Z(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n323), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR4_X1   g492(.A1(new_n658), .A2(new_n276), .A3(new_n322), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n674), .A2(new_n627), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XNOR2_X1  g495(.A(new_n609), .B(KEYINPUT38), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n322), .B1(new_n648), .B2(new_n649), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n678), .B(KEYINPUT39), .Z(new_n684));
  AND2_X1   g498(.A1(new_n426), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n489), .A2(new_n493), .A3(new_n495), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n687), .A2(KEYINPUT106), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n475), .B1(new_n687), .B2(KEYINPUT106), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n274), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI22_X1  g504(.A1(G472), .A2(new_n690), .B1(new_n492), .B2(KEYINPUT32), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n513), .A3(new_n514), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n692), .A2(new_n610), .A3(new_n669), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n682), .A2(new_n683), .A3(new_n686), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n292), .ZN(G45));
  OR2_X1    g509(.A1(new_n640), .A2(KEYINPUT104), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n641), .A3(new_n643), .ZN(new_n697));
  INV_X1    g511(.A(new_n678), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n697), .B(new_n698), .C1(new_n270), .C2(new_n276), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n674), .A2(new_n700), .A3(new_n627), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NAND2_X1  g516(.A1(new_n417), .A2(new_n335), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n417), .A2(new_n335), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n704), .A2(new_n705), .A3(new_n334), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n515), .A2(new_n555), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n651), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT41), .B(G113), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NOR2_X1   g524(.A1(new_n660), .A2(new_n707), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n278), .ZN(G18));
  NAND4_X1  g526(.A1(new_n277), .A2(new_n515), .A3(new_n332), .A4(new_n668), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n605), .B1(new_n587), .B2(new_n598), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n602), .A2(new_n606), .A3(new_n603), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n610), .B(new_n706), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT107), .B(G119), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G21));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n620), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(KEYINPUT108), .B(G472), .C1(new_n510), .C2(G902), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n496), .A2(new_n481), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n489), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n479), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n428), .A3(new_n274), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n723), .A2(new_n555), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n331), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n704), .A2(new_n705), .A3(new_n729), .A4(new_n334), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n627), .A3(new_n683), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  AND3_X1   g546(.A1(new_n723), .A2(new_n668), .A3(new_n727), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n700), .A2(new_n733), .A3(new_n627), .A4(new_n706), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  INV_X1    g549(.A(new_n336), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n703), .A2(new_n425), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n333), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT109), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n426), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n610), .A3(new_n608), .A4(new_n607), .ZN(new_n743));
  INV_X1    g557(.A(new_n555), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n511), .B2(new_n508), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n700), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT42), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n607), .A2(new_n610), .A3(new_n608), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n699), .A2(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n557), .A3(new_n742), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n217), .ZN(G33));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n607), .A2(new_n610), .A3(new_n608), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n426), .B(KEYINPUT109), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n754), .A2(new_n556), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n753), .B1(new_n756), .B2(new_n679), .ZN(new_n757));
  INV_X1    g571(.A(new_n679), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n743), .A2(new_n758), .A3(KEYINPUT110), .A4(new_n556), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n296), .ZN(G36));
  OAI21_X1  g575(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n335), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n736), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n704), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n333), .A3(new_n684), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT111), .Z(new_n771));
  NAND2_X1  g585(.A1(new_n277), .A2(new_n697), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n621), .A3(new_n668), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n771), .A2(new_n748), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NAND2_X1  g594(.A1(new_n769), .A2(new_n333), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n769), .A2(KEYINPUT47), .A3(new_n333), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n754), .A2(new_n515), .A3(new_n555), .A4(new_n699), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NOR2_X1   g602(.A1(new_n704), .A2(new_n705), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT112), .Z(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n613), .B(new_n334), .C1(new_n791), .C2(KEYINPUT49), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(KEYINPUT49), .B2(new_n791), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n692), .A2(new_n744), .ZN(new_n794));
  OR4_X1    g608(.A1(new_n682), .A2(new_n793), .A3(new_n772), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n329), .ZN(new_n797));
  INV_X1    g611(.A(new_n706), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n754), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n799), .A3(new_n277), .A4(new_n645), .ZN(new_n800));
  INV_X1    g614(.A(new_n675), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n774), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT118), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n799), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(KEYINPUT120), .A3(new_n733), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT120), .B1(new_n804), .B2(new_n733), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n800), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n803), .A2(new_n728), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n783), .B2(new_n784), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n790), .A2(new_n334), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n785), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n809), .B(new_n748), .C1(new_n810), .C2(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n682), .A2(new_n610), .A3(new_n798), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n809), .A2(KEYINPUT50), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT50), .B1(new_n809), .B2(new_n815), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n796), .B1(new_n808), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n804), .A2(new_n745), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT48), .Z(new_n822));
  NAND3_X1  g636(.A1(new_n809), .A2(new_n627), .A3(new_n706), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n797), .A2(new_n799), .A3(new_n650), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n327), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n783), .A2(new_n784), .A3(new_n811), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n809), .A2(new_n748), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT51), .ZN(new_n829));
  INV_X1    g643(.A(new_n818), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n816), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(new_n808), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n808), .A2(new_n832), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n820), .B(new_n826), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n674), .B(new_n627), .C1(new_n700), .C2(new_n679), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n738), .A2(new_n668), .A3(new_n678), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n627), .A2(new_n838), .A3(new_n683), .A4(new_n692), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n734), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n837), .A2(KEYINPUT52), .A3(new_n734), .A4(new_n839), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT114), .B1(new_n842), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n625), .A2(new_n729), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n270), .A2(new_n276), .A3(new_n322), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n650), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n847), .B(new_n850), .C1(new_n611), .C2(new_n614), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n851), .A2(new_n615), .A3(new_n671), .ZN(new_n852));
  INV_X1    g666(.A(new_n707), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n613), .B(new_n729), .C1(new_n608), .C2(new_n626), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n853), .B(new_n854), .C1(new_n650), .C2(new_n659), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n717), .A3(new_n731), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n700), .A2(new_n733), .A3(new_n742), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n322), .A2(new_n698), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n658), .A2(new_n276), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n674), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n754), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n751), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n757), .A2(new_n759), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n852), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n836), .B1(new_n846), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n707), .B1(new_n660), .B2(new_n651), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n627), .A2(new_n683), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n730), .A2(new_n555), .A3(new_n723), .A4(new_n727), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n869), .A2(new_n870), .B1(new_n713), .B2(new_n716), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n857), .A2(new_n860), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n748), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n747), .A3(new_n874), .A4(new_n750), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n760), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n876), .B(new_n852), .C1(new_n845), .C2(new_n844), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(KEYINPUT115), .A3(new_n836), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n843), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n842), .A2(new_n880), .A3(new_n843), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n876), .A2(new_n852), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT116), .B1(new_n883), .B2(new_n836), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n881), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n864), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT53), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n879), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n883), .A2(new_n836), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n836), .B2(new_n877), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n891), .B2(new_n894), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n835), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n795), .B1(new_n898), .B2(new_n899), .ZN(G75));
  AOI21_X1  g714(.A(new_n274), .B1(new_n879), .B2(new_n889), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(G210), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n581), .B(new_n585), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n902), .B2(new_n903), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n208), .A2(G952), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  AOI211_X1 g723(.A(new_n274), .B(new_n765), .C1(new_n879), .C2(new_n889), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n336), .B(KEYINPUT57), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n879), .A2(new_n890), .A3(new_n889), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n890), .B1(new_n879), .B2(new_n889), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n405), .A2(new_n416), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n916), .B2(new_n908), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n918));
  INV_X1    g732(.A(new_n908), .ZN(new_n919));
  INV_X1    g733(.A(new_n915), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n865), .A2(new_n866), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT115), .B1(new_n877), .B2(new_n836), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n887), .B1(new_n886), .B2(KEYINPUT53), .ZN(new_n923));
  NOR4_X1   g737(.A1(new_n864), .A2(new_n885), .A3(KEYINPUT116), .A4(new_n836), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n921), .A2(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n891), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n920), .B1(new_n927), .B2(new_n911), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n918), .B(new_n919), .C1(new_n928), .C2(new_n910), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n917), .A2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  INV_X1    g745(.A(new_n657), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n908), .ZN(G60));
  INV_X1    g749(.A(new_n637), .ZN(new_n936));
  INV_X1    g750(.A(new_n639), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n936), .A2(new_n937), .B1(new_n631), .B2(new_n629), .ZN(new_n938));
  XOR2_X1   g752(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n633), .A2(new_n274), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n927), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n919), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n896), .B2(new_n897), .ZN(new_n944));
  INV_X1    g758(.A(new_n938), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(G63));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT60), .Z(new_n948));
  NAND3_X1  g762(.A1(new_n925), .A2(new_n666), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n925), .A2(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n919), .B(new_n949), .C1(new_n950), .C2(new_n554), .ZN(new_n951));
  XOR2_X1   g765(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G66));
  INV_X1    g767(.A(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n324), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n852), .A2(new_n872), .ZN(new_n956));
  INV_X1    g770(.A(new_n208), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n601), .B(new_n575), .C1(G898), .C2(new_n208), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  NAND2_X1  g774(.A1(new_n225), .A2(new_n226), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n503), .B(new_n961), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n957), .A2(G900), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n771), .A2(new_n627), .A3(new_n683), .A4(new_n745), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n837), .A2(new_n734), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n751), .B(new_n965), .C1(new_n785), .C2(new_n786), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n779), .A2(new_n964), .A3(new_n863), .A4(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n962), .B(new_n963), .C1(new_n967), .C2(new_n957), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n850), .A2(new_n748), .A3(new_n557), .A4(new_n685), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n779), .A2(new_n787), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n694), .A2(new_n965), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(new_n973), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT125), .Z(new_n977));
  AOI21_X1  g791(.A(new_n957), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n968), .B1(new_n978), .B2(new_n962), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n208), .B1(G227), .B2(G900), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n968), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n979), .B(new_n982), .Z(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n967), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n956), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n504), .A2(new_n473), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n919), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n975), .A2(new_n956), .A3(new_n977), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n473), .B(new_n504), .C1(new_n991), .C2(new_n985), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n504), .A2(new_n474), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n986), .B1(new_n993), .B2(new_n475), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n990), .B(new_n992), .C1(new_n893), .C2(new_n994), .ZN(G57));
endmodule


