//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981;
  AND2_X1   g000(.A1(G197gat), .A2(G204gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(KEYINPUT73), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n204), .A2(new_n205), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(G183gat), .A3(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n219), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(KEYINPUT25), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n227), .A2(KEYINPUT25), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n214), .A2(KEYINPUT66), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT66), .B1(new_n214), .B2(new_n236), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n216), .B(new_n235), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245));
  AOI21_X1  g044(.A(G190gat), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT28), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT27), .B(G183gat), .ZN(new_n248));
  INV_X1    g047(.A(G190gat), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n248), .A2(KEYINPUT28), .A3(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n220), .B(new_n239), .C1(new_n247), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n234), .A2(new_n251), .B1(new_n255), .B2(new_n252), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n213), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n251), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n255), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n213), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n253), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n260), .B2(new_n253), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT74), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n270), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(KEYINPUT37), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n254), .A2(new_n256), .A3(new_n213), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT37), .B1(new_n277), .B2(new_n265), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT87), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT38), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(KEYINPUT37), .C1(new_n277), .C2(new_n265), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n271), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT37), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n280), .B1(new_n275), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G127gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G127gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT67), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G113gat), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G113gat), .A2(G120gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n290), .B(new_n295), .C1(KEYINPUT1), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n305));
  NAND4_X1  g104(.A1(new_n302), .A2(new_n288), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308));
  AND2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT79), .B(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G155gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n313), .B2(KEYINPUT2), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT77), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G148gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n318), .A3(G141gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n315), .A2(G141gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n319), .B2(new_n322), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n314), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G148gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n321), .A2(new_n330), .B1(new_n309), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n309), .B2(new_n310), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n307), .A2(new_n308), .A3(new_n326), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT81), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n334), .ZN(new_n338));
  INV_X1    g137(.A(new_n325), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n323), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n340), .B2(new_n314), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n341), .A2(KEYINPUT81), .A3(new_n308), .A4(new_n307), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n307), .A2(new_n326), .A3(new_n334), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT4), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n337), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n334), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n301), .A2(new_n306), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n301), .B2(new_n306), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n326), .A2(new_n352), .A3(new_n334), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT82), .B1(new_n345), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n342), .A3(new_n344), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n355), .A4(new_n354), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n301), .A2(new_n306), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT80), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n301), .A2(new_n306), .A3(new_n348), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n355), .B1(new_n365), .B2(new_n343), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n365), .A2(new_n343), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT83), .B(KEYINPUT5), .C1(new_n369), .C2(new_n355), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n357), .A2(new_n360), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n308), .B1(new_n341), .B2(new_n307), .ZN(new_n372));
  INV_X1    g171(.A(new_n335), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT84), .B1(new_n374), .B2(new_n356), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT5), .B1(new_n344), .B2(new_n335), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n355), .A4(new_n354), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n360), .A2(new_n370), .A3(new_n368), .ZN(new_n388));
  INV_X1    g187(.A(new_n356), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n359), .B1(new_n389), .B2(new_n358), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n379), .B(new_n384), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n387), .B(new_n384), .C1(new_n371), .C2(new_n379), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n287), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT31), .B(G50gat), .ZN(new_n396));
  INV_X1    g195(.A(G106gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n209), .A2(new_n255), .A3(new_n212), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n400), .A2(KEYINPUT86), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n352), .B1(new_n400), .B2(KEYINPUT86), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n346), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n353), .A2(new_n255), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n213), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n406), .B(KEYINPUT85), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n206), .A2(new_n208), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n255), .B1(new_n210), .B2(new_n207), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n352), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n346), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n405), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n409), .A2(G22gat), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n416), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n408), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n417), .A2(new_n420), .A3(G78gat), .ZN(new_n421));
  INV_X1    g220(.A(G78gat), .ZN(new_n422));
  OAI21_X1  g221(.A(G22gat), .B1(new_n409), .B2(new_n416), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n418), .A3(new_n408), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n399), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(G78gat), .B1(new_n417), .B2(new_n420), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n422), .A3(new_n424), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n398), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n271), .A2(KEYINPUT30), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n267), .A2(new_n432), .A3(new_n270), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT75), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n273), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n369), .A2(new_n355), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n344), .A2(new_n335), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n355), .B1(new_n439), .B2(new_n354), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  OR3_X1    g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n385), .B1(new_n440), .B2(new_n441), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT40), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(KEYINPUT40), .A3(new_n443), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n437), .A2(new_n386), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n395), .A2(new_n430), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n437), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n391), .A2(new_n387), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n384), .B1(new_n371), .B2(new_n379), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n450), .B1(new_n453), .B2(new_n393), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n426), .A2(new_n429), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n258), .A2(new_n307), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n234), .A2(new_n251), .A3(new_n362), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n457), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n458), .A2(G227gat), .A3(G233gat), .A4(new_n460), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT32), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(new_n457), .C1(new_n459), .C2(new_n461), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G15gat), .B(G43gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT70), .ZN(new_n473));
  XOR2_X1   g272(.A(G71gat), .B(G99gat), .Z(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n471), .B1(new_n469), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n467), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n469), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n470), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n481), .A2(new_n466), .A3(new_n464), .A4(new_n476), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n483), .A2(KEYINPUT72), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n449), .A2(new_n456), .A3(new_n489), .ZN(new_n490));
  AND4_X1   g289(.A1(KEYINPUT88), .A2(new_n426), .A3(new_n429), .A4(new_n483), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n437), .B1(new_n392), .B2(new_n394), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT35), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n426), .A2(KEYINPUT88), .A3(new_n483), .A4(new_n429), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n454), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(G197gat), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT11), .B(G169gat), .Z(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n502), .B(KEYINPUT12), .Z(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  NOR3_X1   g304(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT89), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  INV_X1    g313(.A(G36gat), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n512), .A2(new_n513), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n505), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n505), .A2(new_n519), .ZN(new_n520));
  OAI221_X1 g319(.A(new_n520), .B1(KEYINPUT15), .B2(new_n504), .C1(new_n506), .C2(new_n508), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(G1gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G1gat), .B2(new_n523), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n518), .A2(new_n521), .A3(new_n528), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT13), .Z(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(KEYINPUT92), .A3(new_n529), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n534), .ZN(new_n539));
  INV_X1    g338(.A(new_n530), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n518), .A2(KEYINPUT17), .A3(new_n521), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT91), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n518), .A2(new_n543), .A3(KEYINPUT17), .A4(new_n521), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n529), .B1(new_n522), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g346(.A(new_n539), .B(new_n540), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n538), .B1(new_n548), .B2(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n547), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n534), .A4(new_n530), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n503), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n534), .A3(new_n530), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n537), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n503), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n551), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n498), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  INV_X1    g360(.A(G57gat), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT93), .B1(new_n562), .B2(G64gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n565), .A3(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(G64gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n571), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n569), .ZN(new_n575));
  XNOR2_X1  g374(.A(G57gat), .B(G64gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n528), .B1(new_n561), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT96), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n561), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n586), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n585), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n588), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n582), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n588), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n592), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n581), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(new_n601), .A3(new_n597), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT99), .ZN(new_n607));
  AND2_X1   g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT41), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n607), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT7), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT98), .B1(new_n613), .B2(KEYINPUT7), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT7), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n618), .A2(new_n619), .A3(G85gat), .A4(G92gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n613), .A2(KEYINPUT97), .A3(KEYINPUT7), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n616), .A2(new_n617), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(G85gat), .A2(G92gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(KEYINPUT8), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n622), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n624), .B1(new_n622), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n522), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n610), .B2(new_n609), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n522), .B2(new_n546), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(new_n545), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n606), .A2(KEYINPUT99), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n612), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT100), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n634), .A2(new_n635), .A3(new_n612), .ZN(new_n641));
  OR3_X1    g440(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n637), .B2(new_n641), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n605), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n623), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n573), .A2(new_n578), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n628), .B2(new_n629), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n622), .A2(new_n627), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n623), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n573), .A2(new_n578), .A3(new_n646), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n622), .A2(new_n624), .A3(new_n627), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n654), .A2(KEYINPUT103), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT103), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n648), .A2(new_n653), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT102), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n648), .A2(new_n653), .A3(new_n663), .A4(new_n660), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR4_X1   g464(.A1(new_n628), .A2(new_n629), .A3(new_n660), .A4(new_n579), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n655), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n659), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n668), .A2(KEYINPUT104), .A3(new_n655), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n666), .B1(new_n662), .B2(new_n664), .ZN(new_n678));
  INV_X1    g477(.A(new_n655), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n658), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n675), .B1(new_n681), .B2(new_n672), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT104), .B1(new_n668), .B2(new_n655), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n678), .A2(new_n677), .A3(new_n679), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n659), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n672), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(KEYINPUT105), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n674), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n644), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n560), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n453), .A2(new_n393), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g494(.A1(new_n560), .A2(new_n437), .A3(new_n690), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  AOI21_X1  g498(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n696), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n701), .A2(KEYINPUT42), .A3(new_n699), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT107), .B1(new_n698), .B2(new_n527), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(KEYINPUT106), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n696), .A2(new_n697), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n705), .A2(new_n706), .A3(G8gat), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n703), .A2(new_n709), .ZN(G1325gat));
  OAI21_X1  g509(.A(G15gat), .B1(new_n691), .B2(new_n489), .ZN(new_n711));
  INV_X1    g510(.A(new_n483), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(G15gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n691), .B2(new_n713), .ZN(G1326gat));
  NOR2_X1   g513(.A1(new_n691), .A2(new_n430), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT43), .B(G22gat), .Z(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NAND2_X1  g516(.A1(new_n642), .A2(new_n643), .ZN(new_n718));
  INV_X1    g517(.A(new_n605), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT105), .B1(new_n685), .B2(new_n686), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n681), .A2(new_n675), .A3(new_n672), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n673), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n718), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n560), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n514), .A3(new_n692), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  INV_X1    g526(.A(new_n718), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n490), .B2(new_n497), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(KEYINPUT44), .B(new_n728), .C1(new_n490), .C2(new_n497), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n722), .B(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n554), .A2(new_n555), .ZN(new_n735));
  AND4_X1   g534(.A1(new_n557), .A2(new_n735), .A3(new_n551), .A4(new_n538), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n557), .B1(new_n556), .B2(new_n551), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n734), .A2(new_n738), .A3(new_n719), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(new_n732), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n731), .A2(new_n742), .A3(new_n732), .A4(new_n739), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n741), .A2(new_n692), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n727), .B1(new_n514), .B2(new_n744), .ZN(G1328gat));
  AOI21_X1  g544(.A(G36gat), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n725), .A2(new_n437), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n741), .A2(new_n437), .A3(new_n743), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n515), .B2(new_n750), .ZN(G1329gat));
  NOR3_X1   g550(.A1(new_n724), .A2(G43gat), .A3(new_n712), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G43gat), .B1(new_n740), .B2(new_n489), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(KEYINPUT47), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n489), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n756), .A3(new_n743), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n757), .A2(KEYINPUT111), .A3(G43gat), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT111), .B1(new_n757), .B2(G43gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(new_n752), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n760), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g560(.A1(new_n430), .A2(G50gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT112), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n725), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G50gat), .B1(new_n740), .B2(new_n430), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(KEYINPUT48), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n741), .A2(new_n455), .A3(new_n743), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n767), .A2(G50gat), .B1(new_n725), .B2(new_n763), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n768), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g568(.A1(new_n738), .A2(new_n498), .A3(new_n644), .A4(new_n734), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n692), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n437), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT49), .B(G64gat), .Z(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT113), .ZN(G1333gat));
  NAND2_X1  g576(.A1(new_n770), .A2(new_n756), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n712), .A2(G71gat), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n778), .A2(G71gat), .B1(new_n770), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n770), .A2(new_n455), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n693), .A2(G85gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n498), .A2(KEYINPUT115), .A3(new_n728), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n719), .A2(new_n559), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n729), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AND4_X1   g590(.A1(KEYINPUT51), .A2(new_n785), .A3(new_n786), .A4(new_n790), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n722), .B(new_n784), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n731), .A2(new_n732), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n786), .A2(new_n722), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT114), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n692), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G85gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n793), .A2(new_n799), .ZN(G1336gat));
  NOR2_X1   g599(.A1(new_n450), .A2(G92gat), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n734), .B(new_n801), .C1(new_n791), .C2(new_n792), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n794), .A2(new_n437), .A3(new_n796), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT116), .B1(new_n803), .B2(G92gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1337gat));
  NOR2_X1   g608(.A1(new_n712), .A2(G99gat), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n722), .B(new_n810), .C1(new_n791), .C2(new_n792), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n756), .A3(new_n796), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n794), .A2(KEYINPUT117), .A3(new_n756), .A4(new_n796), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(G99gat), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT118), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n811), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1338gat));
  NOR2_X1   g620(.A1(new_n430), .A2(G106gat), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n734), .B(new_n822), .C1(new_n791), .C2(new_n792), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n797), .A2(new_n455), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G106gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n676), .A2(new_n832), .A3(new_n680), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n686), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT54), .B1(new_n678), .B2(new_n679), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n678), .B2(new_n679), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n678), .A2(new_n836), .A3(new_n679), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n831), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n839), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT54), .B(new_n669), .C1(new_n842), .C2(new_n837), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(KEYINPUT55), .A3(new_n686), .A4(new_n833), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n673), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n534), .B1(new_n550), .B2(new_n530), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n535), .B1(new_n533), .B2(new_n536), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n502), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n558), .A2(new_n848), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n718), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n849), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n722), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT120), .B1(new_n688), .B2(new_n849), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n559), .A2(new_n673), .A3(new_n844), .A4(new_n841), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n850), .B1(new_n856), .B2(new_n728), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n605), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n644), .A2(new_n738), .A3(new_n688), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n693), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND4_X1   g659(.A1(new_n430), .A2(new_n860), .A3(new_n450), .A4(new_n483), .ZN(new_n861));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n559), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n455), .B1(new_n858), .B2(new_n859), .ZN(new_n863));
  AND4_X1   g662(.A1(new_n692), .A2(new_n863), .A3(new_n450), .A4(new_n483), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n738), .A2(new_n296), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(G120gat), .B1(new_n861), .B2(new_n722), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n733), .A2(new_n297), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n864), .B2(new_n868), .ZN(G1341gat));
  NAND3_X1  g668(.A1(new_n861), .A2(new_n291), .A3(new_n719), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n864), .A2(new_n719), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n291), .ZN(G1342gat));
  NAND3_X1  g671(.A1(new_n861), .A2(new_n293), .A3(new_n728), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT56), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n864), .A2(new_n728), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n874), .B(new_n875), .C1(new_n293), .C2(new_n876), .ZN(G1343gat));
  AOI21_X1  g676(.A(new_n430), .B1(new_n858), .B2(new_n859), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n688), .A2(new_n849), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n738), .B1(new_n845), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n841), .A2(new_n844), .A3(KEYINPUT121), .A4(new_n673), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n850), .B1(new_n885), .B2(new_n728), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n886), .A2(new_n605), .B1(new_n738), .B2(new_n690), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n430), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n756), .A2(new_n693), .A3(new_n437), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G141gat), .B1(new_n890), .B2(new_n738), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n489), .A2(KEYINPUT122), .A3(new_n455), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT122), .B1(new_n489), .B2(new_n455), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n437), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n860), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n329), .A3(new_n559), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n859), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n644), .A2(KEYINPUT123), .A3(new_n738), .A4(new_n688), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n886), .B2(new_n605), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n879), .B1(new_n903), .B2(new_n430), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT124), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n906), .B(new_n879), .C1(new_n903), .C2(new_n430), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n722), .A3(new_n889), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n316), .A2(new_n318), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n912), .A3(new_n722), .ZN(new_n913));
  INV_X1    g712(.A(new_n890), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(new_n722), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n911), .B(new_n913), .C1(KEYINPUT59), .C2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n890), .B2(new_n605), .ZN(new_n917));
  INV_X1    g716(.A(G155gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n895), .A2(new_n918), .A3(new_n719), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1346gat));
  OAI21_X1  g719(.A(new_n312), .B1(new_n890), .B2(new_n718), .ZN(new_n921));
  INV_X1    g720(.A(new_n312), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n895), .A2(new_n922), .A3(new_n728), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n692), .A2(new_n450), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n712), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n863), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n738), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n692), .B1(new_n858), .B2(new_n859), .ZN(new_n930));
  AND4_X1   g729(.A1(new_n430), .A2(new_n930), .A3(new_n437), .A4(new_n483), .ZN(new_n931));
  INV_X1    g730(.A(G169gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(new_n559), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(KEYINPUT125), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(KEYINPUT125), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(G1348gat));
  INV_X1    g735(.A(new_n928), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(G176gat), .A3(new_n734), .ZN(new_n938));
  AOI21_X1  g737(.A(G176gat), .B1(new_n931), .B2(new_n722), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1349gat));
  NAND3_X1  g741(.A1(new_n931), .A2(new_n248), .A3(new_n719), .ZN(new_n943));
  OAI21_X1  g742(.A(G183gat), .B1(new_n928), .B2(new_n605), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n249), .A3(new_n728), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n937), .A2(new_n728), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(G190gat), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT61), .B(new_n249), .C1(new_n937), .C2(new_n728), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NOR3_X1   g751(.A1(new_n756), .A2(new_n430), .A3(new_n450), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n930), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n559), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n926), .A2(new_n756), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI22_X1  g757(.A1(new_n904), .A2(KEYINPUT124), .B1(new_n878), .B2(KEYINPUT57), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n907), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n559), .A2(G197gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n734), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n954), .A2(G204gat), .A3(new_n688), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1353gat));
  OR3_X1    g766(.A1(new_n954), .A2(G211gat), .A3(new_n605), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n909), .A2(new_n719), .A3(new_n957), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  INV_X1    g772(.A(G218gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n960), .B2(new_n728), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n954), .A2(G218gat), .A3(new_n718), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n909), .A2(new_n728), .A3(new_n957), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G218gat), .ZN(new_n979));
  INV_X1    g778(.A(new_n976), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n979), .A2(KEYINPUT127), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n977), .A2(new_n981), .ZN(G1355gat));
endmodule


