//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n551, new_n553,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT68), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n478), .B2(G2105), .ZN(G160));
  NOR2_X1   g054(.A1(new_n466), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(new_n465), .A3(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n480), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n495), .A2(new_n465), .A3(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT69), .B1(new_n475), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n493), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .A3(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n507), .A2(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT71), .B(G88), .Z(new_n516));
  OAI21_X1  g091(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n513), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n506), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n517), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  XOR2_X1   g097(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n514), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n510), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n512), .A2(new_n513), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G651), .B1(G52), .B2(new_n510), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n514), .A2(G90), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n506), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n514), .A2(G81), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n510), .A2(G43), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n510), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n533), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(G91), .B2(new_n514), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n510), .A2(G49), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT75), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n518), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n514), .B2(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n512), .B2(new_n513), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n510), .A2(G48), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n507), .A2(new_n509), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n578), .A2(G86), .A3(new_n518), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n506), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n514), .A2(G85), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n510), .A2(G47), .ZN(new_n584));
  NOR3_X1   g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(new_n514), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  AOI22_X1  g166(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n506), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n510), .A2(KEYINPUT78), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n578), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n593), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n591), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g177(.A(new_n601), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G168), .B2(new_n604), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(G168), .B2(new_n604), .ZN(G280));
  INV_X1    g182(.A(new_n600), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT79), .B(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(G860), .B2(new_n609), .ZN(G148));
  NAND2_X1  g185(.A1(new_n548), .A2(new_n604), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n609), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n613), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n481), .A2(G2104), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(KEYINPUT80), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n483), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n465), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT81), .B(G2096), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n618), .B1(KEYINPUT80), .B2(new_n620), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n622), .B(new_n629), .C1(new_n630), .C2(new_n621), .ZN(G156));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT85), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G1341), .ZN(new_n634));
  INV_X1    g209(.A(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT83), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(G2438), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(KEYINPUT83), .ZN(new_n641));
  INV_X1    g216(.A(new_n639), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n640), .A2(new_n643), .A3(new_n645), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT14), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n647), .B2(KEYINPUT14), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n646), .B(new_n653), .C1(new_n649), .C2(new_n650), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n636), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n656), .A3(new_n636), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n663), .B2(KEYINPUT87), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(KEYINPUT87), .B2(new_n663), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n663), .B(KEYINPUT17), .Z(new_n668));
  INV_X1    g243(.A(new_n662), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n665), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n663), .A3(new_n662), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n669), .A3(new_n666), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G1986), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT89), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n683), .B(KEYINPUT19), .ZN(new_n692));
  INV_X1    g267(.A(new_n688), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n687), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n682), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G1981), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n689), .B(KEYINPUT20), .ZN(new_n700));
  INV_X1    g275(.A(new_n697), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(KEYINPUT89), .A3(new_n701), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n699), .B1(new_n698), .B2(new_n702), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n681), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n691), .A2(new_n682), .A3(new_n697), .ZN(new_n709));
  AOI21_X1  g284(.A(KEYINPUT89), .B1(new_n700), .B2(new_n701), .ZN(new_n710));
  OAI21_X1  g285(.A(G1981), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n711), .A2(G1986), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n705), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n708), .B1(new_n705), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n680), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n713), .ZN(new_n717));
  AOI21_X1  g292(.A(G1986), .B1(new_n711), .B2(new_n712), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n707), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n705), .A2(new_n708), .A3(new_n713), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n719), .A2(new_n679), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(new_n721), .ZN(G229));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G23), .ZN(new_n724));
  INV_X1    g299(.A(G288), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT33), .B(G1976), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n723), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n723), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1971), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n723), .A2(G6), .ZN(new_n732));
  INV_X1    g307(.A(G305), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n723), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT32), .B(G1981), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n734), .B(new_n736), .Z(new_n737));
  NOR3_X1   g312(.A1(new_n728), .A2(new_n731), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n481), .A2(G131), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n483), .A2(G119), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n465), .A2(G107), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n742), .B(new_n743), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G25), .B(new_n746), .S(G29), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(G16), .A2(G24), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G290), .B2(new_n723), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n749), .B1(new_n751), .B2(new_n681), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n681), .B2(new_n751), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n740), .A2(new_n741), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(KEYINPUT36), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT30), .B(G28), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n627), .B2(new_n759), .ZN(new_n763));
  NOR2_X1   g338(.A1(G162), .A2(new_n759), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n759), .B2(G35), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT29), .B(G2090), .Z(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n759), .A2(G32), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n470), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(G105), .B2(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(G129), .A2(new_n483), .B1(new_n481), .B2(G141), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(KEYINPUT97), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n774), .A2(new_n778), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n769), .B1(new_n781), .B2(new_n759), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT27), .B(G1996), .Z(new_n783));
  AOI21_X1  g358(.A(new_n768), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n759), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT94), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n481), .A2(G140), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n483), .A2(G128), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n791));
  AND3_X1   g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(new_n759), .ZN(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n759), .A2(G33), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n481), .A2(G139), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT95), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT25), .Z(new_n800));
  AOI22_X1  g375(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n465), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n759), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G2072), .ZN(new_n805));
  NOR2_X1   g380(.A1(G168), .A2(new_n723), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n723), .B2(G21), .ZN(new_n807));
  INV_X1    g382(.A(G1966), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n807), .A2(new_n808), .B1(G2072), .B2(new_n804), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n784), .A2(new_n795), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n759), .A2(G27), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G164), .B2(new_n759), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2078), .ZN(new_n813));
  NAND2_X1  g388(.A1(G160), .A2(G29), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT24), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(G34), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n759), .B1(new_n815), .B2(G34), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n813), .B1(G2084), .B2(new_n819), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n820), .B1(G2084), .B2(new_n819), .C1(new_n782), .C2(new_n783), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n723), .A2(G19), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n549), .B2(new_n723), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G1341), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n723), .A2(G20), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT23), .Z(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G299), .B2(G16), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1956), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n824), .B(new_n828), .C1(new_n808), .C2(new_n807), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n810), .A2(new_n821), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n723), .A2(G5), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G171), .B2(new_n723), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G1961), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT98), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n608), .A2(G16), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G4), .B2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT93), .B(G1348), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n832), .A2(G1961), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n834), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n757), .A2(new_n830), .A3(new_n841), .ZN(G311));
  INV_X1    g417(.A(G311), .ZN(G150));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n533), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n506), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  AOI22_X1  g424(.A1(G93), .A2(new_n514), .B1(new_n510), .B2(G55), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G860), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n849), .A2(new_n855), .A3(new_n850), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n849), .B2(new_n850), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n548), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(KEYINPUT101), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n849), .A2(new_n855), .A3(new_n850), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n549), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n608), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n866), .B2(KEYINPUT39), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n854), .B1(new_n867), .B2(new_n869), .ZN(G145));
  XNOR2_X1  g445(.A(KEYINPUT106), .B(G37), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n481), .A2(G142), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n483), .A2(G130), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(G118), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n875), .A2(KEYINPUT105), .B1(new_n876), .B2(G2105), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(KEYINPUT105), .B2(new_n875), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n777), .A2(new_n779), .A3(new_n792), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n792), .B1(new_n777), .B2(new_n779), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n792), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n780), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(new_n881), .A3(new_n879), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n494), .B1(new_n480), .B2(new_n496), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n475), .A2(new_n498), .A3(KEYINPUT69), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n502), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT103), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n502), .A2(new_n889), .A3(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n493), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n489), .A2(new_n492), .A3(KEYINPUT104), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n893), .A2(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n803), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n502), .A2(new_n889), .A3(new_n894), .A4(new_n890), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n798), .B2(new_n802), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n617), .B(new_n746), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n888), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(new_n887), .A3(new_n884), .A4(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(G160), .B(new_n627), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n487), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n916), .A3(new_n911), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n872), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g494(.A(G288), .B(G303), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n587), .A2(G305), .A3(new_n588), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G305), .B1(new_n587), .B2(new_n588), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n920), .A3(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n558), .A2(new_n562), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n591), .A3(new_n599), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n600), .A2(G299), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n862), .A2(new_n613), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n858), .A2(new_n861), .A3(new_n612), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n932), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n858), .A2(new_n861), .A3(new_n612), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n612), .B1(new_n858), .B2(new_n861), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n939), .B2(new_n943), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n928), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n949));
  INV_X1    g524(.A(new_n928), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n952), .A3(G868), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT107), .B1(new_n851), .B2(new_n604), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n947), .A2(new_n952), .A3(KEYINPUT107), .A4(G868), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(G295));
  AND2_X1   g535(.A1(new_n955), .A2(new_n957), .ZN(G331));
  AOI21_X1  g536(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(new_n935), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n940), .A2(KEYINPUT110), .A3(new_n934), .ZN(new_n965));
  INV_X1    g540(.A(new_n541), .ZN(new_n966));
  NAND3_X1  g541(.A1(G168), .A2(new_n539), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(G286), .B1(new_n540), .B2(new_n541), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n856), .A2(new_n857), .A3(new_n548), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n549), .B1(new_n859), .B2(new_n860), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n858), .A2(new_n861), .A3(new_n968), .A4(new_n967), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n964), .A2(new_n965), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n940), .A3(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n950), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n936), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n940), .A3(new_n973), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n928), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n871), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n972), .A2(new_n973), .B1(new_n935), .B2(new_n933), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n950), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G37), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n980), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n982), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n976), .A2(new_n989), .A3(new_n980), .A4(new_n871), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(G397));
  INV_X1    g568(.A(KEYINPUT60), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n995), .B(new_n471), .C1(new_n478), .C2(G2105), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  INV_X1    g572(.A(new_n493), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n891), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n902), .A2(new_n997), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n635), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n902), .A2(new_n1002), .A3(new_n996), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n902), .A2(new_n996), .A3(KEYINPUT119), .A4(new_n1002), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n600), .B(new_n1005), .C1(new_n1010), .C2(G2067), .ZN(new_n1011));
  AOI21_X1  g586(.A(G2067), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1348), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n608), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n994), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1016), .B(new_n1017), .C1(G164), .C2(G1384), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT113), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n902), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT56), .B(G2072), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1020), .A2(new_n996), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1956), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n997), .B1(new_n902), .B2(new_n1002), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1002), .B1(new_n893), .B2(new_n493), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n996), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n1030));
  XNOR2_X1  g605(.A(G299), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1023), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT61), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1015), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT58), .B(G1341), .Z(new_n1038));
  NAND3_X1  g613(.A1(new_n1008), .A2(new_n1009), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1996), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1020), .A2(new_n1040), .A3(new_n996), .A4(new_n1021), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n548), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1037), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT59), .B1(new_n1042), .B2(KEYINPUT121), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1046), .B(new_n548), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n549), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1046), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(KEYINPUT121), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1037), .A3(KEYINPUT59), .A4(new_n1052), .ZN(new_n1053));
  NOR4_X1   g628(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT60), .A4(new_n600), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1023), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1031), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1054), .B1(new_n1057), .B2(KEYINPUT61), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1036), .A2(new_n1048), .A3(new_n1053), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1033), .B1(new_n1055), .B2(new_n1014), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1020), .A2(new_n1064), .A3(new_n996), .A4(new_n1021), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  INV_X1    g641(.A(G1961), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1065), .A2(new_n1066), .B1(new_n1004), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT45), .B1(new_n902), .B2(new_n1002), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1026), .A2(new_n1017), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G160), .A2(G40), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1066), .A2(G2078), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(G301), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n902), .A2(new_n1002), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1017), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(KEYINPUT123), .A3(new_n996), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1080), .A3(new_n1021), .A4(new_n1073), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1068), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1083), .A2(KEYINPUT124), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(KEYINPUT124), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT54), .B(new_n1075), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1001), .A2(new_n1087), .A3(new_n1003), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(G168), .C1(new_n1072), .C2(G1966), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(G8), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1072), .A2(G1966), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1088), .ZN(new_n1094));
  OAI21_X1  g669(.A(G286), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(G8), .A3(new_n1089), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1096), .B2(KEYINPUT51), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G305), .A2(G1981), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n576), .A2(new_n577), .A3(new_n579), .A4(new_n699), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT49), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(KEYINPUT49), .A3(new_n1099), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1098), .A2(KEYINPUT114), .A3(KEYINPUT49), .A4(new_n1099), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1006), .A2(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n565), .A2(G1976), .A3(new_n567), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1006), .A2(G8), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT52), .ZN(new_n1110));
  INV_X1    g685(.A(G1976), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(G288), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(G8), .A3(new_n1006), .A4(new_n1108), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT115), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1107), .A2(new_n1116), .A3(new_n1113), .A4(new_n1110), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(G303), .A2(G8), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT55), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1016), .B1(new_n1026), .B2(new_n1017), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n999), .A2(KEYINPUT113), .A3(KEYINPUT45), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n996), .B(new_n1021), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1971), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1004), .A2(G2090), .ZN(new_n1127));
  OAI211_X1 g702(.A(G8), .B(new_n1121), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1025), .A2(new_n1027), .A3(G2090), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1130));
  INV_X1    g705(.A(G8), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1120), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1118), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1004), .A2(new_n1067), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1074), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1068), .A2(new_n1081), .A3(G301), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT54), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1097), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1063), .A2(new_n1086), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1384), .B1(new_n898), .B2(new_n892), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1000), .B1(new_n1142), .B2(new_n997), .ZN(new_n1143));
  INV_X1    g718(.A(G2090), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1125), .A2(new_n1124), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1120), .B1(new_n1145), .B2(new_n1131), .ZN(new_n1146));
  AND4_X1   g721(.A1(KEYINPUT63), .A2(new_n1107), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1147));
  NAND2_X1  g722(.A1(G168), .A2(G8), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1070), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1077), .A2(new_n996), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n808), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1151), .B2(new_n1088), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(new_n1128), .A3(new_n1147), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1118), .A2(new_n1128), .A3(new_n1132), .A4(new_n1152), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1156), .A2(KEYINPUT116), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1156), .B2(KEYINPUT116), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1155), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1106), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n725), .A2(new_n1111), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1107), .A2(new_n1163), .B1(new_n699), .B2(new_n733), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1128), .A2(new_n1114), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1089), .A2(G8), .ZN(new_n1167));
  AOI21_X1  g742(.A(G168), .B1(new_n1151), .B2(new_n1088), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT51), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n1169), .B2(new_n1091), .ZN(new_n1170));
  AOI21_X1  g745(.A(G301), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1118), .A2(new_n1128), .A3(new_n1132), .A4(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1097), .A2(new_n1166), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1165), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1141), .A2(new_n1160), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1069), .A2(new_n996), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT111), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1178), .A2(G1996), .A3(new_n780), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1177), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(new_n1040), .A3(new_n781), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n792), .B(new_n794), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT112), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1187));
  INV_X1    g762(.A(new_n748), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n746), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n746), .A2(new_n1188), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1178), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1186), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(G290), .A2(G1986), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n681), .B1(new_n587), .B2(new_n588), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1192), .B1(new_n1180), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1176), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1180), .A2(new_n1040), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT46), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(KEYINPUT125), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1198), .B(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1178), .A2(new_n780), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1199), .A2(KEYINPUT125), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1201), .A2(new_n1202), .A3(new_n1183), .A4(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT47), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1193), .A2(new_n1180), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT48), .Z(new_n1207));
  OAI21_X1  g782(.A(new_n1205), .B1(new_n1192), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1178), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n792), .A2(new_n794), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1197), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g789(.A1(G227), .A2(new_n463), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1216), .B1(new_n659), .B2(new_n660), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n716), .A2(new_n721), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1218), .A2(KEYINPUT126), .ZN(new_n1219));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n1220));
  NAND4_X1  g794(.A1(new_n716), .A2(new_n721), .A3(new_n1217), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g796(.A(new_n918), .B1(new_n988), .B2(new_n990), .ZN(new_n1223));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1224), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
  NAND2_X1  g801(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n1228), .A2(KEYINPUT127), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n1229), .A2(new_n1230), .ZN(G225));
endmodule


