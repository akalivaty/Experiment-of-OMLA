//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n202), .B(new_n205), .C1(new_n206), .C2(KEYINPUT2), .ZN(new_n207));
  AND2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT75), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(new_n211), .A3(new_n202), .ZN(new_n212));
  AND2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n202), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT76), .B1(new_n202), .B2(KEYINPUT2), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n207), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n221));
  INV_X1    g020(.A(G134gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G127gat), .ZN(new_n223));
  INV_X1    g022(.A(G127gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G134gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G113gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(G113gat), .ZN(new_n231));
  INV_X1    g030(.A(G113gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n223), .A2(new_n225), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n240), .B(new_n207), .C1(new_n216), .C2(new_n219), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT77), .B1(new_n220), .B2(KEYINPUT3), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT78), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n241), .A2(new_n239), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .A4(new_n221), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n220), .A2(new_n239), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT4), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n249), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n251), .B1(new_n244), .B2(new_n248), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(KEYINPUT81), .A3(new_n255), .ZN(new_n260));
  INV_X1    g059(.A(new_n231), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n229), .A2(G113gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n226), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n236), .B1(new_n227), .B2(new_n234), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT2), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n208), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n202), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(new_n215), .A3(new_n212), .A4(new_n210), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n270), .A3(new_n207), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT4), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n220), .A2(new_n239), .A3(KEYINPUT4), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(KEYINPUT79), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT79), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n275), .A3(KEYINPUT4), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n254), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n249), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT80), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n264), .B1(new_n207), .B2(new_n270), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n254), .B1(new_n280), .B2(new_n250), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n281), .B2(KEYINPUT5), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n220), .A2(new_n239), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n253), .B1(new_n283), .B2(new_n271), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n284), .A2(KEYINPUT80), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n258), .A2(new_n260), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G1gat), .B(G29gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT0), .ZN(new_n291));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n258), .A2(new_n288), .A3(new_n293), .A4(new_n260), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n289), .A2(KEYINPUT6), .A3(new_n294), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(G211gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G218gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G197gat), .B(G204gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  NAND3_X1  g115(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G183gat), .B2(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT24), .B1(new_n321), .B2(KEYINPUT65), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT23), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT25), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n316), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n329), .B1(KEYINPUT23), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n326), .A2(KEYINPUT25), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n321), .A2(KEYINPUT65), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n320), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  AND2_X1   g138(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n335), .A2(new_n342), .A3(KEYINPUT66), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n325), .A2(KEYINPUT64), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G176gat), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT23), .A4(new_n324), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n337), .ZN(new_n348));
  OR2_X1    g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n317), .ZN(new_n350));
  INV_X1    g149(.A(new_n329), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n332), .A2(KEYINPUT23), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n331), .A2(new_n343), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT27), .B(G183gat), .ZN(new_n358));
  INV_X1    g157(.A(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(KEYINPUT28), .A3(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT26), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n351), .A2(new_n365), .A3(new_n332), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n329), .A2(KEYINPUT26), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n367), .A2(new_n321), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n315), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n314), .B1(new_n357), .B2(new_n369), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n313), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g176(.A(KEYINPUT73), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n368), .A2(new_n366), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n362), .B2(new_n363), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n335), .A2(new_n342), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n381), .A2(new_n316), .B1(new_n355), .B2(new_n354), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n382), .B2(new_n343), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n378), .B1(new_n383), .B2(new_n314), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n373), .A2(KEYINPUT73), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n357), .B2(new_n369), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n312), .B1(new_n387), .B2(new_n315), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n374), .B(new_n377), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT30), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(KEYINPUT74), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n377), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT73), .B1(new_n370), .B2(new_n315), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n378), .B(new_n314), .C1(new_n357), .C2(new_n369), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n388), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n314), .B1(new_n383), .B2(KEYINPUT29), .ZN(new_n400));
  INV_X1    g199(.A(new_n373), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n312), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n396), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n400), .A2(new_n384), .A3(new_n312), .A4(new_n385), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n404), .A2(KEYINPUT30), .A3(new_n374), .A4(new_n377), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n301), .B1(new_n395), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n405), .ZN(new_n408));
  AOI211_X1 g207(.A(KEYINPUT89), .B(new_n408), .C1(new_n393), .C2(new_n394), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n300), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT92), .ZN(new_n411));
  INV_X1    g210(.A(new_n394), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT74), .B1(new_n389), .B2(new_n390), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT89), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n406), .B(new_n301), .C1(new_n412), .C2(new_n413), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n300), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  INV_X1    g219(.A(G50gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT83), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n311), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n308), .B1(new_n305), .B2(new_n306), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n371), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT3), .B1(new_n429), .B2(KEYINPUT84), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n310), .B2(new_n311), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n430), .A2(new_n433), .B1(new_n207), .B2(new_n270), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n241), .A2(new_n371), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n313), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n426), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n220), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n439), .A2(G228gat), .A3(G233gat), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n312), .B1(new_n443), .B2(new_n435), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n241), .A2(KEYINPUT85), .A3(new_n371), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT87), .B(G22gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n438), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n438), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n425), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G22gat), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n438), .B2(new_n449), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n425), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n451), .B(new_n460), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n454), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G15gat), .B(G43gat), .Z(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT69), .ZN(new_n464));
  XNOR2_X1  g263(.A(G71gat), .B(G99gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n383), .A2(new_n239), .ZN(new_n467));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n370), .A2(new_n264), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n474), .A3(new_n476), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n469), .B1(new_n467), .B2(new_n470), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT71), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT34), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n471), .A2(new_n472), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT33), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n480), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n493));
  INV_X1    g292(.A(new_n479), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n493), .B(new_n466), .C1(new_n494), .C2(new_n477), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(new_n490), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n485), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT35), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n462), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n411), .A2(new_n419), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n486), .B1(new_n480), .B2(new_n491), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n495), .A2(new_n496), .A3(new_n485), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n456), .A2(new_n457), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n505), .A2(new_n451), .A3(new_n460), .A4(new_n458), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n506), .B2(new_n454), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n414), .B1(new_n298), .B2(new_n299), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n399), .A2(new_n402), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n377), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n512), .B2(new_n511), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT38), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n400), .A2(new_n401), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n512), .B1(new_n516), .B2(new_n312), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n400), .A2(new_n384), .A3(new_n313), .A4(new_n385), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT38), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n513), .A2(new_n519), .B1(new_n511), .B2(new_n377), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n515), .A2(new_n298), .A3(new_n299), .A4(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT39), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n249), .A2(new_n252), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(new_n254), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n259), .A2(KEYINPUT90), .A3(new_n253), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n523), .A3(new_n254), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT90), .B1(new_n259), .B2(new_n253), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n280), .A2(new_n250), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n522), .B1(new_n530), .B2(new_n253), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n527), .A2(KEYINPUT40), .A3(new_n293), .A4(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n527), .A2(new_n293), .A3(new_n532), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT40), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n415), .A2(new_n538), .A3(new_n295), .A4(new_n416), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n462), .B(new_n521), .C1(new_n535), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n508), .ZN(new_n541));
  INV_X1    g340(.A(new_n462), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n492), .B2(new_n497), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n501), .A2(new_n510), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(G1gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n550), .B(new_n551), .C1(G1gat), .C2(new_n548), .ZN(new_n552));
  NOR2_X1   g351(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT97), .Z(new_n555));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OR3_X1    g356(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n559), .B2(new_n558), .ZN(new_n561));
  INV_X1    g360(.A(G29gat), .ZN(new_n562));
  INV_X1    g361(.A(G36gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n421), .A2(G43gat), .ZN(new_n565));
  INV_X1    g364(.A(G43gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G50gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n567), .A2(KEYINPUT95), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(new_n565), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(KEYINPUT95), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT15), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n575), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n558), .A2(new_n556), .B1(G29gat), .B2(G36gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n570), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT98), .B1(new_n555), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n555), .A2(new_n580), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n554), .B(KEYINPUT97), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584));
  INV_X1    g383(.A(new_n580), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT13), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(KEYINPUT17), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n580), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n554), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n582), .A2(new_n588), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT18), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n587), .A2(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G197gat), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT11), .B(G169gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT12), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n596), .A2(new_n605), .A3(new_n597), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT7), .ZN(new_n609));
  INV_X1    g408(.A(G99gat), .ZN(new_n610));
  INV_X1    g409(.A(G106gat), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT8), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n609), .B(new_n612), .C1(G85gat), .C2(G92gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G99gat), .B(G106gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n590), .A2(new_n592), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n580), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT101), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n620), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT102), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n626), .A2(KEYINPUT102), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G71gat), .B(G78gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G57gat), .B(G64gat), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n634), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n634), .B(new_n633), .C1(new_n637), .C2(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n583), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n645));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n644), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT100), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n648), .B(new_n654), .Z(new_n655));
  NOR2_X1   g454(.A1(new_n632), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n642), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n642), .B1(KEYINPUT103), .B2(new_n614), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n616), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n659), .B2(KEYINPUT10), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G120gat), .B(G148gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT104), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n661), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n662), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n660), .A2(KEYINPUT106), .A3(new_n661), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n672), .A2(new_n673), .B1(new_n668), .B2(new_n659), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n666), .B(KEYINPUT105), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n670), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n656), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n547), .A2(new_n607), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n300), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT107), .B(G1gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1324gat));
  NOR2_X1   g483(.A1(new_n407), .A2(new_n409), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n686), .A2(G8gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n688), .B1(new_n694), .B2(new_n689), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n692), .B1(new_n693), .B2(new_n695), .ZN(G1325gat));
  INV_X1    g495(.A(new_n680), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n545), .A2(new_n543), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n504), .A2(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n697), .B2(new_n700), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n680), .A2(new_n542), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n547), .B2(new_n631), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n462), .A2(new_n498), .A3(new_n499), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(KEYINPUT92), .B2(new_n410), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(new_n419), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n698), .B1(new_n462), .B2(new_n508), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n533), .B(KEYINPUT91), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n712), .A2(new_n685), .A3(new_n295), .A4(new_n538), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n521), .A2(new_n462), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT44), .B(new_n632), .C1(new_n710), .C2(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n706), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n655), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n607), .A2(new_n718), .A3(new_n677), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n300), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n547), .A2(new_n631), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n681), .A2(new_n562), .ZN(new_n724));
  OR3_X1    g523(.A1(new_n723), .A2(KEYINPUT109), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT109), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n721), .B1(new_n728), .B2(new_n729), .ZN(G1328gat));
  OAI21_X1  g529(.A(G36gat), .B1(new_n720), .B2(new_n417), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n723), .A2(G36gat), .A3(new_n417), .ZN(new_n732));
  NAND2_X1  g531(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n735));
  OAI211_X1 g534(.A(new_n731), .B(new_n734), .C1(new_n732), .C2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n698), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n706), .A2(new_n737), .A3(new_n716), .A4(new_n719), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G43gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n504), .A2(G43gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n719), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(new_n741), .A3(KEYINPUT47), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743));
  INV_X1    g542(.A(new_n741), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n739), .B2(KEYINPUT111), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n738), .A2(new_n746), .A3(G43gat), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n743), .B(KEYINPUT47), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n739), .A2(KEYINPUT111), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n747), .A3(new_n741), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT112), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n742), .B1(new_n748), .B2(new_n752), .ZN(G1330gat));
  OAI21_X1  g552(.A(new_n421), .B1(new_n723), .B2(new_n462), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n542), .A2(G50gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n720), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g556(.A(new_n547), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n604), .A2(new_n606), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n632), .A2(new_n678), .A3(new_n759), .A4(new_n655), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n681), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n761), .A2(new_n417), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  NOR3_X1   g568(.A1(new_n761), .A2(G71gat), .A3(new_n504), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n762), .A2(new_n737), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(G71gat), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g572(.A1(new_n761), .A2(new_n462), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT113), .B(G78gat), .Z(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n759), .A2(new_n718), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n722), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n678), .A2(G85gat), .A3(new_n300), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n678), .A2(new_n759), .A3(new_n718), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n717), .A2(new_n681), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G85gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n717), .A2(new_n685), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G92gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n678), .A2(G92gat), .A3(new_n417), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n778), .A2(KEYINPUT114), .A3(new_n779), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n779), .A2(KEYINPUT114), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n722), .A2(new_n777), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n790), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n794), .B2(KEYINPUT115), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n794), .A2(KEYINPUT115), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(new_n780), .B2(new_n789), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n788), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1337gat));
  NAND4_X1  g599(.A1(new_n780), .A2(new_n610), .A3(new_n498), .A4(new_n677), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n717), .A2(new_n737), .A3(new_n783), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n610), .B2(new_n802), .ZN(G1338gat));
  NOR3_X1   g602(.A1(new_n678), .A2(G106gat), .A3(new_n462), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n780), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n706), .A2(new_n542), .A3(new_n716), .A4(new_n783), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n793), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n804), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n807), .A2(new_n809), .B1(new_n811), .B2(new_n806), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n685), .A2(new_n300), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n672), .A2(new_n673), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n660), .B2(new_n661), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n668), .B(new_n657), .C1(new_n659), .C2(KEYINPUT10), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n667), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n670), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT55), .B1(new_n816), .B2(new_n820), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT117), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n816), .A2(new_n820), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n670), .A4(new_n821), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n759), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n587), .A2(new_n589), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n588), .B1(new_n582), .B2(new_n593), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n602), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n606), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n677), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n632), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n606), .B2(new_n833), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n631), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n837), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n824), .A2(new_n839), .A3(new_n829), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n655), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n656), .A2(new_n607), .A3(new_n678), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n814), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n507), .ZN(new_n845));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n759), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n542), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n814), .A2(new_n504), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(new_n232), .A3(new_n607), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n846), .A2(new_n850), .ZN(G1340gat));
  NAND2_X1  g650(.A1(new_n677), .A2(new_n229), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT120), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n677), .A3(new_n848), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(KEYINPUT119), .A3(G120gat), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT119), .B1(new_n855), .B2(G120gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n845), .A2(new_n224), .A3(new_n718), .ZN(new_n859));
  OAI21_X1  g658(.A(G127gat), .B1(new_n849), .B2(new_n655), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1342gat));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n222), .A3(new_n632), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n849), .B2(new_n631), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1343gat));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n814), .A2(new_n737), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n842), .A2(new_n843), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n542), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n542), .A2(KEYINPUT57), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT121), .B1(new_n834), .B2(new_n677), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n607), .A2(new_n822), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n825), .A2(KEYINPUT122), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n825), .A2(KEYINPUT122), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n826), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n834), .A2(KEYINPUT121), .A3(new_n677), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n632), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n655), .B1(new_n881), .B2(new_n841), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n873), .B1(new_n882), .B2(new_n843), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n759), .B(new_n870), .C1(new_n872), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n737), .A2(new_n462), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n607), .A2(G141gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n844), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n869), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g691(.A(new_n868), .B(new_n890), .C1(new_n884), .C2(G141gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(G1344gat));
  INV_X1    g693(.A(new_n822), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n895), .A2(new_n839), .A3(new_n827), .A4(new_n840), .ZN(new_n896));
  INV_X1    g695(.A(new_n874), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n876), .A2(new_n826), .A3(new_n877), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n759), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n897), .B(new_n880), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n900), .B2(new_n631), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n843), .B1(new_n901), .B2(new_n718), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n902), .B2(new_n542), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n873), .B1(new_n842), .B2(new_n843), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n870), .A2(new_n677), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT59), .B(G148gat), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n872), .A2(new_n883), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n677), .A4(new_n870), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n844), .A2(new_n886), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n911), .B2(new_n677), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n907), .B(new_n910), .C1(G148gat), .C2(new_n912), .ZN(G1345gat));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n203), .A3(new_n718), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n908), .A2(new_n718), .A3(new_n870), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n203), .ZN(G1346gat));
  NAND2_X1  g715(.A1(new_n911), .A2(new_n632), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n204), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n631), .A2(new_n204), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n870), .B(new_n919), .C1(new_n872), .C2(new_n883), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n918), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n681), .A2(new_n417), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n871), .A2(new_n507), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n759), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n926), .B(KEYINPUT125), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n847), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(new_n498), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n607), .A2(new_n324), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(G1348gat));
  AOI21_X1  g733(.A(G176gat), .B1(new_n927), .B2(new_n677), .ZN(new_n935));
  AOI211_X1 g734(.A(new_n504), .B(new_n678), .C1(new_n344), .C2(new_n346), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n931), .B2(new_n936), .ZN(G1349gat));
  NAND3_X1  g736(.A1(new_n927), .A2(new_n358), .A3(new_n718), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n847), .A2(new_n498), .A3(new_n718), .A4(new_n930), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G183gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n941), .B(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n359), .A3(new_n632), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n931), .A2(new_n498), .A3(new_n632), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(G190gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n946), .B2(G190gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  AND3_X1   g749(.A1(new_n871), .A2(new_n886), .A3(new_n926), .ZN(new_n951));
  AOI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n759), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n929), .A2(new_n737), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n903), .B2(new_n904), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n759), .A2(G197gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n678), .A2(G204gat), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n951), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(G204gat), .B1(new_n954), .B2(new_n678), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n960), .A2(KEYINPUT62), .A3(new_n962), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(G1353gat));
  NOR2_X1   g767(.A1(new_n655), .A2(new_n302), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n718), .B(new_n953), .C1(new_n903), .C2(new_n904), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  OAI21_X1  g773(.A(G218gat), .B1(new_n954), .B2(new_n631), .ZN(new_n975));
  INV_X1    g774(.A(G218gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n951), .A2(new_n976), .A3(new_n632), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1355gat));
endmodule


