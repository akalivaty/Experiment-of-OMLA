//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n441, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G120), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(new_n441), .A2(G57), .A3(G69), .A4(G108), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  XOR2_X1   g039(.A(KEYINPUT3), .B(G2104), .Z(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n474), .A2(G101), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  OR2_X1    g052(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n474), .B2(new_n476), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(G2104), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n470), .A2(G137), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n478), .A2(new_n479), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n467), .A2(new_n487), .A3(new_n471), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n473), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  OAI21_X1  g065(.A(KEYINPUT71), .B1(new_n481), .B2(new_n483), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(new_n495), .A3(new_n482), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(G136), .A3(new_n475), .ZN(new_n498));
  NOR2_X1   g073(.A1(G100), .A2(G2105), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT72), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n471), .ZN(new_n502));
  INV_X1    g077(.A(G124), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n498), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G162));
  XNOR2_X1  g080(.A(KEYINPUT3), .B(G2104), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n470), .A2(new_n506), .A3(G138), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(G102), .A2(G2105), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n510), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n511));
  INV_X1    g086(.A(G138), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n468), .B2(new_n469), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(KEYINPUT4), .B1(G126), .B2(G2105), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n494), .A2(new_n482), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n509), .B(new_n511), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n521), .A3(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT5), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n524), .B1(new_n531), .B2(new_n518), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT6), .B(G651), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n530), .A2(KEYINPUT74), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT74), .B1(new_n530), .B2(new_n533), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n532), .B1(G88), .B2(new_n536), .ZN(G166));
  AND3_X1   g112(.A1(new_n528), .A2(KEYINPUT5), .A3(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(G543), .B1(new_n528), .B2(KEYINPUT5), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n530), .A2(KEYINPUT74), .A3(new_n533), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G89), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n522), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n533), .A2(KEYINPUT75), .A3(G543), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(new_n549), .A3(G51), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n544), .A2(new_n546), .A3(new_n550), .A4(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  AOI22_X1  g128(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n554), .A2(new_n555), .A3(new_n518), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n554), .B2(new_n518), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n542), .A2(G90), .A3(new_n543), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n548), .A2(new_n549), .A3(G52), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(G301));
  INV_X1    g139(.A(G301), .ZN(G171));
  AND3_X1   g140(.A1(new_n542), .A2(G81), .A3(new_n543), .ZN(new_n566));
  INV_X1    g141(.A(G56), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n527), .B2(new_n529), .ZN(new_n568));
  AND2_X1   g143(.A1(G68), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n548), .A2(new_n549), .ZN(new_n571));
  INV_X1    g146(.A(G43), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  AND3_X1   g150(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G36), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT78), .ZN(G188));
  AOI22_X1  g156(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n518), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(new_n534), .B2(new_n535), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n542), .A2(KEYINPUT80), .A3(new_n543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n583), .B1(new_n587), .B2(G91), .ZN(new_n588));
  INV_X1    g163(.A(G53), .ZN(new_n589));
  NOR3_X1   g164(.A1(new_n522), .A2(KEYINPUT79), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT9), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G166), .ZN(G303));
  NAND2_X1  g168(.A1(new_n587), .A2(G87), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT81), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n523), .A2(G49), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(G288));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n585), .B2(new_n586), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n523), .A2(G48), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n530), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n518), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n542), .A2(new_n543), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT82), .B(G85), .Z(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G47), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n571), .A2(new_n609), .B1(new_n610), .B2(new_n518), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n571), .A2(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n571), .A2(KEYINPUT83), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(G54), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT85), .B(G66), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n530), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT84), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n518), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT10), .B1(new_n587), .B2(G92), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  AOI211_X1 g201(.A(new_n625), .B(new_n626), .C1(new_n585), .C2(new_n586), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n617), .B(new_n623), .C1(new_n624), .C2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n614), .B1(new_n629), .B2(G868), .ZN(G284));
  OAI21_X1  g205(.A(new_n614), .B1(new_n629), .B2(G868), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  INV_X1    g207(.A(G299), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G297));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n629), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n574), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g216(.A1(new_n497), .A2(G123), .A3(new_n471), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n497), .A2(G135), .A3(new_n475), .ZN(new_n643));
  OAI221_X1 g218(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G2096), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NOR4_X1   g222(.A1(new_n465), .A2(G2105), .A3(new_n493), .A4(new_n492), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT13), .B(G2100), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2435), .ZN(new_n661));
  XOR2_X1   g236(.A(G2427), .B(G2438), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT14), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT87), .Z(G401));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2067), .B(G2678), .Z(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(new_n673), .ZN(new_n678));
  INV_X1    g253(.A(new_n672), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n669), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n669), .A3(new_n673), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT18), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n676), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n646), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  INV_X1    g260(.A(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n689), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n693), .A2(KEYINPUT20), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n689), .A3(new_n692), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n696), .B(new_n698), .C1(KEYINPUT20), .C2(new_n693), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT90), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n702), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G35), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G29), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n504), .B2(G29), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI211_X1 g286(.A(KEYINPUT29), .B(new_n708), .C1(new_n504), .C2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(G2090), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G20), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT23), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT23), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G299), .B2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(new_n719), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n713), .B1(G1956), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G1956), .B2(new_n720), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n711), .A2(new_n712), .A3(G2090), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G26), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n491), .A2(G128), .A3(new_n471), .A4(new_n496), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n491), .A2(G140), .A3(new_n475), .A4(new_n496), .ZN(new_n727));
  OAI221_X1 g302(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(new_n724), .ZN(new_n731));
  MUX2_X1   g306(.A(new_n725), .B(new_n731), .S(KEYINPUT28), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  INV_X1    g308(.A(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT96), .B1(new_n734), .B2(G16), .ZN(new_n735));
  OR3_X1    g310(.A1(new_n734), .A2(KEYINPUT96), .A3(G16), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n735), .B(new_n736), .C1(new_n574), .C2(new_n714), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1341), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT94), .B1(G4), .B2(G16), .ZN(new_n740));
  OR3_X1    g315(.A1(KEYINPUT94), .A2(G4), .A3(G16), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n740), .B(new_n741), .C1(new_n628), .C2(new_n714), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT95), .B(G1348), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n722), .A2(new_n723), .A3(new_n739), .A4(new_n744), .ZN(new_n745));
  OR3_X1    g320(.A1(G286), .A2(KEYINPUT102), .A3(new_n714), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  OR2_X1    g322(.A1(G16), .A2(G21), .ZN(new_n748));
  OAI211_X1 g323(.A(KEYINPUT102), .B(new_n748), .C1(G286), .C2(new_n714), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n747), .B1(new_n746), .B2(new_n749), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n642), .A2(new_n643), .A3(G29), .A4(new_n644), .ZN(new_n753));
  INV_X1    g328(.A(G28), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT30), .B2(new_n754), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n751), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT103), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(G5), .A2(G16), .ZN(new_n762));
  OAI211_X1 g337(.A(G1961), .B(new_n762), .C1(G301), .C2(new_n714), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n758), .A2(new_n759), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n746), .A2(new_n749), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G1966), .ZN(new_n766));
  INV_X1    g341(.A(new_n757), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n766), .A2(new_n763), .A3(new_n750), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(KEYINPUT103), .B1(new_n768), .B2(new_n760), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT101), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G29), .B2(G32), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT100), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT26), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n491), .A2(G141), .A3(new_n475), .A4(new_n496), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n491), .A2(G129), .A3(new_n471), .A4(new_n496), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n474), .A2(G105), .A3(new_n475), .A4(new_n476), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT99), .ZN(new_n779));
  AND4_X1   g354(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT27), .B(G1996), .Z(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n780), .A2(G29), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n784), .C1(new_n771), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n771), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n783), .B1(new_n787), .B2(new_n781), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n762), .B1(G301), .B2(new_n714), .ZN(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(KEYINPUT24), .A2(G34), .ZN(new_n792));
  NOR2_X1   g367(.A1(KEYINPUT24), .A2(G34), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n792), .A2(new_n793), .A3(G29), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n489), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2084), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n786), .A2(new_n788), .A3(new_n791), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G29), .A2(G33), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n491), .A2(G139), .A3(new_n475), .A4(new_n496), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n506), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(new_n470), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n470), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n800), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n800), .A2(new_n807), .A3(new_n802), .A4(KEYINPUT97), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n810), .A2(KEYINPUT98), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(KEYINPUT98), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n799), .B1(new_n814), .B2(new_n724), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2072), .ZN(new_n816));
  INV_X1    g391(.A(G2072), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(new_n799), .C1(new_n814), .C2(new_n724), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n797), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n724), .A2(G27), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G164), .B2(new_n724), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT104), .B(G2078), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n770), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT105), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n770), .A2(new_n819), .A3(KEYINPUT105), .A4(new_n823), .ZN(new_n827));
  AOI211_X1 g402(.A(KEYINPUT106), .B(new_n745), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT106), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  INV_X1    g405(.A(new_n745), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n497), .A2(G119), .A3(new_n471), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n497), .A2(G131), .A3(new_n475), .ZN(new_n834));
  OAI221_X1 g409(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n724), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G1991), .ZN(new_n841));
  NOR2_X1   g416(.A1(G25), .A2(G29), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n714), .A2(G24), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n612), .B2(new_n714), .ZN(new_n847));
  INV_X1    g422(.A(G1986), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G1976), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n714), .A2(G23), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G288), .B2(G16), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n587), .A2(G87), .B1(G49), .B2(new_n523), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n714), .B1(new_n855), .B2(new_n596), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n856), .A2(KEYINPUT33), .A3(new_n851), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n850), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n714), .A2(G22), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G303), .B2(G16), .ZN(new_n860));
  INV_X1    g435(.A(G1971), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n852), .A2(new_n853), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT33), .B1(new_n856), .B2(new_n851), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(G1976), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n860), .A2(new_n861), .ZN(new_n866));
  OAI21_X1  g441(.A(G16), .B1(new_n600), .B2(new_n603), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT32), .B(G1981), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n714), .A2(G6), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n867), .B2(new_n870), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n858), .A2(new_n862), .A3(new_n865), .A4(new_n873), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n845), .B(new_n849), .C1(new_n874), .C2(KEYINPUT34), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT93), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(KEYINPUT34), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT92), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT92), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n880), .A3(KEYINPUT34), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n876), .A2(new_n877), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT36), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n879), .A2(new_n881), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n877), .B1(new_n884), .B2(new_n876), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n828), .A2(new_n832), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT36), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n886), .A2(new_n889), .ZN(G311));
  OAI221_X1 g465(.A(new_n888), .B1(new_n885), .B2(new_n883), .C1(new_n828), .C2(new_n832), .ZN(G150));
  NOR2_X1   g466(.A1(new_n628), .A2(new_n636), .ZN(new_n892));
  XOR2_X1   g467(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n573), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n536), .A2(G81), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n542), .A2(G93), .A3(new_n543), .ZN(new_n897));
  INV_X1    g472(.A(G55), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n899));
  OAI22_X1  g474(.A1(new_n571), .A2(new_n898), .B1(new_n899), .B2(new_n518), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n900), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n548), .A2(new_n549), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n530), .A2(G67), .ZN(new_n903));
  NAND2_X1  g478(.A1(G80), .A2(G543), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n902), .A2(G55), .B1(new_n905), .B2(G651), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n536), .A2(G93), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n906), .B(new_n907), .C1(new_n566), .C2(new_n573), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n894), .B(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n911));
  AOI21_X1  g486(.A(G860), .B1(new_n911), .B2(KEYINPUT108), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n912), .B(new_n913), .C1(KEYINPUT108), .C2(new_n911), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n897), .A2(new_n900), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G860), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT37), .Z(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n918), .ZN(G145));
  NAND2_X1  g494(.A1(new_n836), .A2(KEYINPUT109), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n497), .A2(G142), .A3(new_n475), .ZN(new_n921));
  OAI221_X1 g496(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n497), .A2(G130), .A3(new_n471), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n833), .A2(new_n834), .A3(new_n926), .A4(new_n835), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n920), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n920), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n729), .A2(G164), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n516), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(new_n780), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n780), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n934), .A2(new_n935), .B1(new_n812), .B2(new_n813), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n933), .ZN(new_n937));
  INV_X1    g512(.A(new_n780), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n810), .A2(new_n811), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n932), .A2(new_n780), .A3(new_n933), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n936), .A2(new_n650), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n650), .B1(new_n936), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n931), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n650), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT98), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n810), .A2(KEYINPUT98), .A3(new_n811), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n941), .A2(new_n939), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n810), .A2(new_n811), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n934), .A2(new_n935), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n936), .A2(new_n650), .A3(new_n942), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n930), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n945), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G162), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n945), .A2(new_n955), .A3(new_n956), .A4(new_n504), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n645), .B(new_n489), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n961), .A2(new_n962), .A3(G37), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT40), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n963), .B(new_n964), .ZN(G395));
  NAND2_X1  g540(.A1(G288), .A2(G166), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n855), .A2(G303), .A3(new_n596), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n966), .A2(G305), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G305), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(G290), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n604), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(G305), .A3(new_n967), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n612), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n638), .B(new_n909), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n626), .B1(new_n585), .B2(new_n586), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT10), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(G299), .A3(new_n617), .A4(new_n623), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n628), .A2(new_n633), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT41), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT41), .B1(new_n981), .B2(new_n982), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(new_n978), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n977), .B(new_n988), .ZN(new_n989));
  MUX2_X1   g564(.A(new_n916), .B(new_n989), .S(G868), .Z(G295));
  MUX2_X1   g565(.A(new_n916), .B(new_n989), .S(G868), .Z(G331));
  NAND2_X1  g566(.A1(new_n901), .A2(new_n908), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n559), .A2(new_n561), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT77), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G286), .B1(new_n996), .B2(new_n558), .ZN(new_n997));
  OAI211_X1 g572(.A(G286), .B(new_n558), .C1(new_n562), .C2(new_n563), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n992), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G301), .A2(G168), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(new_n909), .A3(new_n998), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n909), .B1(new_n1002), .B2(new_n998), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT112), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n983), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n985), .B2(new_n986), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n975), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT113), .B1(new_n1011), .B2(G37), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1002), .A2(new_n909), .A3(new_n998), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(new_n1005), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT41), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n983), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT41), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n981), .A2(new_n982), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n975), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n970), .A2(new_n974), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n1025));
  INV_X1    g600(.A(G37), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1012), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n987), .A2(new_n1007), .B1(new_n1019), .B2(new_n1009), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1023), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G37), .B1(new_n1021), .B2(new_n975), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(KEYINPUT114), .A3(new_n1023), .ZN(new_n1036));
  AND4_X1   g611(.A1(KEYINPUT43), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT44), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1028), .A2(KEYINPUT43), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1034), .A2(new_n1029), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1043), .ZN(G397));
  XNOR2_X1  g619(.A(G299), .B(KEYINPUT57), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT121), .ZN(new_n1046));
  INV_X1    g621(.A(G1384), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n516), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT45), .ZN(new_n1049));
  AND4_X1   g624(.A1(G40), .A2(new_n473), .A3(new_n486), .A4(new_n488), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n516), .A2(new_n1047), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1049), .A2(new_n1050), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1048), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1050), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1055), .B1(new_n1060), .B2(G1956), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1045), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1049), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1064), .A2(new_n1054), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n628), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1059), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1050), .A2(new_n1070), .A3(new_n1048), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n473), .A2(new_n486), .A3(G40), .A4(new_n488), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT120), .B1(new_n1072), .B2(new_n1051), .ZN(new_n1073));
  INV_X1    g648(.A(G2067), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1046), .A2(new_n1061), .B1(new_n1067), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1996), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1064), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1078), .A2(KEYINPUT122), .A3(new_n1079), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n574), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(KEYINPUT123), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1061), .A2(new_n1045), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT124), .B1(new_n1061), .B2(new_n1045), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1092), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1086), .A2(new_n574), .A3(new_n1089), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT61), .B1(new_n1061), .B2(new_n1045), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1091), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n628), .B1(new_n1076), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT60), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1105), .A2(KEYINPUT125), .A3(new_n628), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1104), .A2(new_n1106), .B1(new_n1101), .B2(new_n1076), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1106), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1076), .A2(new_n1101), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT125), .B1(new_n1105), .B2(new_n628), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1077), .B1(new_n1100), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1050), .A2(new_n1053), .A3(KEYINPUT118), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1049), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n747), .ZN(new_n1119));
  INV_X1    g694(.A(G2084), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1060), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT51), .B(G8), .C1(new_n1122), .C2(G286), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n1124));
  INV_X1    g699(.A(G8), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G168), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1118), .A2(new_n747), .B1(new_n1120), .B2(new_n1060), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1124), .B(new_n1127), .C1(new_n1128), .C2(new_n1125), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1123), .A2(new_n1129), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1063), .A2(new_n861), .ZN(new_n1131));
  INV_X1    g706(.A(G2090), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1057), .A2(new_n1132), .A3(new_n1050), .A4(new_n1058), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1125), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(G303), .A2(G8), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT55), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1063), .B2(G2078), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT126), .B(G1961), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n1059), .A2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1142), .B(G2078), .C1(new_n1048), .C2(KEYINPUT45), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1048), .A2(KEYINPUT115), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1051), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1052), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1150), .A3(new_n472), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n486), .A2(G40), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1143), .B(new_n1145), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G171), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1116), .A2(new_n1146), .A3(new_n1117), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1155), .A2(new_n1143), .A3(G301), .A4(new_n1145), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(KEYINPUT54), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1981), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n604), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n606), .A2(new_n599), .ZN(new_n1160));
  OAI21_X1  g735(.A(G1981), .B1(new_n1160), .B2(new_n603), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(KEYINPUT49), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT116), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT49), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT116), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1159), .A2(new_n1167), .A3(KEYINPUT49), .A4(new_n1161), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1125), .B1(new_n1050), .B2(new_n1048), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1163), .A2(new_n1166), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1169), .ZN(new_n1171));
  NOR2_X1   g746(.A1(G288), .A2(new_n850), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT52), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT52), .B1(G288), .B2(new_n850), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1174), .B(new_n1169), .C1(new_n850), .C2(G288), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1170), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1141), .A2(new_n1157), .A3(new_n1177), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1153), .A2(G171), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1155), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(G171), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT54), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1130), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1113), .A2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1176), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1128), .A2(new_n1125), .A3(G286), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT119), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1185), .A2(new_n1189), .A3(new_n1186), .ZN(new_n1192));
  NOR2_X1   g767(.A1(G288), .A2(G1976), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1170), .A2(new_n1193), .B1(new_n1158), .B2(new_n604), .ZN(new_n1194));
  OAI22_X1  g769(.A1(new_n1194), .A2(new_n1171), .B1(new_n1176), .B2(new_n1138), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT117), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI221_X1 g772(.A(KEYINPUT117), .B1(new_n1176), .B2(new_n1138), .C1(new_n1194), .C2(new_n1171), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1191), .A2(new_n1192), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1181), .B1(new_n1130), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1128), .A2(new_n1127), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT62), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1201), .A2(new_n1204), .A3(new_n1185), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1184), .A2(new_n1199), .A3(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n780), .B(G1996), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n729), .B(new_n1074), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1150), .A2(new_n1072), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n836), .B(new_n841), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n612), .B(new_n848), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1214), .B1(new_n1210), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1206), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1210), .A2(new_n848), .A3(new_n612), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT48), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1219), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1220));
  AOI21_X1  g795(.A(KEYINPUT46), .B1(new_n1210), .B2(new_n1083), .ZN(new_n1221));
  AND3_X1   g796(.A1(new_n1210), .A2(KEYINPUT46), .A3(new_n1083), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1208), .A2(new_n780), .ZN(new_n1223));
  AOI211_X1 g798(.A(new_n1221), .B(new_n1222), .C1(new_n1210), .C2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g799(.A(new_n1224), .B(KEYINPUT47), .ZN(new_n1225));
  AND2_X1   g800(.A1(new_n838), .A2(new_n839), .ZN(new_n1226));
  OR2_X1    g801(.A1(new_n1226), .A2(new_n841), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1211), .ZN(new_n1228));
  OAI22_X1  g803(.A1(new_n1227), .A2(new_n1228), .B1(G2067), .B2(new_n729), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1229), .B(KEYINPUT127), .ZN(new_n1230));
  AOI211_X1 g805(.A(new_n1220), .B(new_n1225), .C1(new_n1210), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1217), .A2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g807(.A(new_n667), .ZN(new_n1234));
  NOR2_X1   g808(.A1(new_n961), .A2(new_n962), .ZN(new_n1235));
  AOI21_X1  g809(.A(new_n1234), .B1(new_n1235), .B2(new_n1026), .ZN(new_n1236));
  OR3_X1    g810(.A1(G227), .A2(new_n462), .A3(G229), .ZN(new_n1237));
  AOI21_X1  g811(.A(new_n1237), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1238));
  AND2_X1   g812(.A1(new_n1236), .A2(new_n1238), .ZN(G308));
  NAND2_X1  g813(.A1(new_n1236), .A2(new_n1238), .ZN(G225));
endmodule


