//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202));
  INV_X1    g001(.A(G8gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT87), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n208), .B2(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n213), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n228), .B(KEYINPUT13), .Z(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n213), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n226), .B1(KEYINPUT88), .B2(KEYINPUT17), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT88), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n224), .A2(new_n225), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(new_n234), .B2(new_n235), .ZN(new_n239));
  INV_X1    g038(.A(new_n236), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n232), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n213), .A2(new_n238), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n228), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n231), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT11), .B(G169gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n242), .A2(KEYINPUT18), .A3(new_n228), .A4(new_n243), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n246), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n246), .B2(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n202), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n251), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(KEYINPUT89), .A3(new_n254), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n262));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G141gat), .B(G148gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT2), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(G141gat), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G141gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G148gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n263), .A2(new_n269), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n273), .A2(new_n275), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G127gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G134gat), .ZN(new_n283));
  INV_X1    g082(.A(G134gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G127gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT68), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G113gat), .B2(G120gat), .ZN(new_n288));
  AND2_X1   g087(.A1(G113gat), .A2(G120gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n279), .B(new_n280), .C1(new_n289), .C2(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n262), .B1(new_n278), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n293), .A3(new_n262), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n295), .A2(KEYINPUT80), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n291), .A2(KEYINPUT77), .A3(new_n292), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n265), .B(new_n264), .C1(new_n267), .C2(KEYINPUT2), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n273), .A2(new_n275), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n276), .A2(new_n265), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT3), .B1(new_n270), .B2(new_n277), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n299), .A2(new_n300), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n295), .B2(KEYINPUT80), .ZN(new_n308));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n297), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n309), .ZN(new_n313));
  INV_X1    g112(.A(new_n296), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(new_n294), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT78), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n295), .A2(new_n296), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n309), .A4(new_n307), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n299), .A2(new_n321), .A3(new_n300), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n278), .A2(new_n293), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n309), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n310), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n312), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G1gat), .B(G29gat), .Z(new_n328));
  XNOR2_X1  g127(.A(G57gat), .B(G85gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  OAI21_X1  g131(.A(KEYINPUT81), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335));
  INV_X1    g134(.A(new_n332), .ZN(new_n336));
  INV_X1    g135(.A(new_n326), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n316), .B2(new_n319), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n336), .C1(new_n338), .C2(new_n312), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n326), .ZN(new_n340));
  INV_X1    g139(.A(new_n312), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n332), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n333), .A2(new_n334), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT6), .B(new_n336), .C1(new_n338), .C2(new_n312), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n347));
  INV_X1    g146(.A(G169gat), .ZN(new_n348));
  INV_X1    g147(.A(G176gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT23), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n350), .A2(KEYINPUT65), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT65), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G190gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(G183gat), .ZN(new_n356));
  INV_X1    g155(.A(G183gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(G190gat), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT24), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n349), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n359), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n347), .B1(new_n354), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n365), .A2(G169gat), .A3(G176gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n351), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n350), .A2(KEYINPUT65), .A3(new_n351), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n357), .A2(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n355), .A2(G183gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n361), .B1(new_n377), .B2(KEYINPUT24), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n374), .A2(KEYINPUT66), .A3(new_n378), .A4(new_n366), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n371), .B1(new_n364), .B2(new_n365), .ZN(new_n380));
  OR2_X1    g179(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n381), .A2(KEYINPUT23), .A3(new_n348), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n359), .A2(new_n380), .A3(new_n362), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n363), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n379), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT27), .B(G183gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n355), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT28), .B1(new_n388), .B2(KEYINPUT67), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391));
  AOI211_X1 g190(.A(new_n390), .B(new_n391), .C1(new_n387), .C2(new_n355), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n364), .A2(KEYINPUT26), .ZN(new_n393));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT26), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n351), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n360), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  OR3_X1    g196(.A1(new_n389), .A2(new_n392), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n386), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n389), .A2(new_n392), .A3(new_n397), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n378), .B(new_n366), .C1(new_n353), .C2(new_n352), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n347), .B1(new_n363), .B2(new_n384), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(new_n379), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n400), .ZN(new_n407));
  XNOR2_X1  g206(.A(G211gat), .B(G218gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G197gat), .B(G204gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT22), .ZN(new_n410));
  INV_X1    g209(.A(G211gat), .ZN(new_n411));
  INV_X1    g210(.A(G218gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n408), .B1(new_n413), .B2(new_n409), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n402), .A2(new_n407), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT72), .B1(new_n399), .B2(new_n401), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT72), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(new_n400), .C1(new_n406), .C2(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n386), .A2(new_n398), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n401), .ZN(new_n425));
  AOI211_X1 g224(.A(KEYINPUT73), .B(new_n400), .C1(new_n386), .C2(new_n398), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n418), .B1(new_n428), .B2(new_n417), .ZN(new_n429));
  XNOR2_X1  g228(.A(G8gat), .B(G36gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  AOI21_X1  g231(.A(new_n346), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n417), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n422), .B2(new_n427), .ZN(new_n435));
  INV_X1    g234(.A(new_n432), .ZN(new_n436));
  NOR4_X1   g235(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n418), .A4(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT74), .ZN(new_n439));
  INV_X1    g238(.A(new_n418), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n426), .B(new_n425), .C1(new_n419), .C2(new_n421), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n439), .B(new_n440), .C1(new_n441), .C2(new_n434), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT74), .B1(new_n435), .B2(new_n418), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT75), .B1(new_n444), .B2(new_n436), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT75), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n446), .B(new_n432), .C1(new_n442), .C2(new_n443), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n345), .B(new_n438), .C1(new_n445), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n293), .ZN(new_n449));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n293), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n386), .A2(new_n452), .A3(new_n398), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G71gat), .B(G99gat), .Z(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(KEYINPUT32), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n454), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n454), .A2(KEYINPUT32), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n454), .A2(new_n458), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n457), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n386), .A2(new_n452), .A3(new_n398), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n452), .B1(new_n386), .B2(new_n398), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n450), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n472), .A2(KEYINPUT71), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n472), .B2(KEYINPUT71), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n465), .A2(new_n476), .A3(new_n468), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n409), .A2(new_n413), .ZN(new_n482));
  INV_X1    g281(.A(new_n408), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT29), .B1(new_n484), .B2(new_n414), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n301), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT29), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n415), .B2(new_n416), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n321), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n305), .A2(new_n488), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n417), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n481), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT82), .B(new_n306), .C1(new_n489), .C2(new_n278), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n321), .C1(new_n485), .C2(KEYINPUT3), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n493), .A2(new_n495), .A3(new_n481), .A4(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(G22gat), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G22gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n486), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n301), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n504), .A2(new_n321), .B1(new_n417), .B2(new_n492), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n501), .B(new_n498), .C1(new_n505), .C2(new_n481), .ZN(new_n506));
  XNOR2_X1  g305(.A(G78gat), .B(G106gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G50gat), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n507), .B(new_n508), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT84), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n509), .A2(KEYINPUT84), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n500), .A2(new_n506), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n511), .B1(new_n500), .B2(new_n506), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n480), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT35), .B1(new_n448), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n465), .A2(new_n476), .A3(new_n468), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n476), .B1(new_n465), .B2(new_n468), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n478), .A2(KEYINPUT85), .A3(new_n479), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n515), .B2(new_n516), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n336), .B1(new_n338), .B2(new_n312), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(new_n334), .A3(new_n342), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(new_n344), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n433), .A2(new_n437), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n428), .A2(new_n417), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n439), .B1(new_n532), .B2(new_n440), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n435), .A2(KEYINPUT74), .A3(new_n418), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n436), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n446), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n444), .A2(KEYINPUT75), .A3(new_n436), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n530), .A2(new_n538), .A3(KEYINPUT86), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT86), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n438), .B1(new_n445), .B2(new_n447), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n519), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n517), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n448), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n480), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n478), .A2(KEYINPUT36), .A3(new_n479), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n325), .B1(new_n297), .B2(new_n308), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n322), .A2(new_n323), .A3(new_n309), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n551), .A2(KEYINPUT39), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n332), .B1(new_n551), .B2(KEYINPUT39), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT40), .ZN(new_n555));
  OR3_X1    g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n527), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n536), .A2(new_n537), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(new_n438), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT38), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n444), .A2(KEYINPUT37), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n432), .B1(new_n429), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n429), .A2(new_n563), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n402), .A2(new_n407), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n563), .B1(new_n567), .B2(new_n417), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(new_n441), .B2(new_n417), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n566), .A2(new_n561), .A3(new_n436), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n429), .A2(new_n432), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n570), .A2(new_n344), .A3(new_n571), .A4(new_n528), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n517), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n546), .B(new_n550), .C1(new_n560), .C2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n261), .B1(new_n544), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT7), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  AOI21_X1  g383(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(new_n587), .B2(new_n586), .ZN(new_n589));
  INV_X1    g388(.A(G64gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(KEYINPUT90), .A3(G57gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(G57gat), .B2(new_n590), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT90), .B1(new_n590), .B2(G57gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G57gat), .B(G64gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI22_X1  g396(.A1(new_n589), .A2(new_n594), .B1(new_n586), .B2(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n584), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n584), .B2(new_n598), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n599), .B(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(new_n604), .B2(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT94), .ZN(new_n606));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n599), .A2(new_n603), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n599), .A2(new_n603), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT10), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n608), .B1(new_n611), .B2(new_n601), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n607), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n614), .A3(new_n610), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n615), .B1(new_n605), .B2(new_n614), .ZN(new_n621));
  INV_X1    g420(.A(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n620), .B1(new_n619), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n282), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n232), .B1(new_n627), .B2(new_n598), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT92), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G155gat), .ZN(new_n636));
  XOR2_X1   g435(.A(G183gat), .B(G211gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G190gat), .B(G218gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n584), .ZN(new_n644));
  NAND2_X1  g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n644), .A2(new_n238), .B1(KEYINPUT41), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n237), .A2(new_n241), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n643), .B(new_n647), .C1(new_n648), .C2(new_n644), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n233), .A2(new_n236), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n239), .A2(new_n240), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n644), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n642), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n646), .A2(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g454(.A(G134gat), .B(G162gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n649), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n649), .B2(new_n654), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n641), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n626), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n575), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n345), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n541), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT16), .B(G8gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT42), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(G8gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT96), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(new_n550), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n523), .A2(new_n524), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n676), .A2(G15gat), .B1(new_n664), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT97), .Z(G1326gat));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n545), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND3_X1  g482(.A1(new_n626), .A2(new_n641), .A3(new_n660), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT98), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n575), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n218), .A3(new_n665), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n660), .A2(KEYINPUT100), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n658), .B2(new_n659), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AOI211_X1 g492(.A(KEYINPUT44), .B(new_n693), .C1(new_n544), .C2(new_n574), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n544), .A2(new_n574), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n660), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT44), .ZN(new_n698));
  INV_X1    g497(.A(new_n660), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n544), .B2(new_n574), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT99), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n694), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n259), .A2(new_n254), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n626), .A2(new_n704), .A3(new_n641), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n703), .A2(new_n345), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n706), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n689), .B1(new_n708), .B2(new_n709), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n686), .A2(G36gat), .A3(new_n538), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n703), .A2(new_n538), .A3(new_n705), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n214), .B2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n677), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n687), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n703), .A2(new_n550), .A3(new_n705), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT47), .B(new_n717), .C1(new_n718), .C2(new_n715), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n718), .B2(new_n715), .ZN(new_n721));
  INV_X1    g520(.A(new_n694), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n697), .B1(new_n696), .B2(KEYINPUT44), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n700), .A2(KEYINPUT99), .A3(new_n701), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n705), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n675), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(KEYINPUT102), .A3(G43gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n721), .A2(new_n728), .A3(new_n717), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n729), .A2(KEYINPUT103), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT103), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n719), .B1(new_n731), .B2(new_n732), .ZN(G1330gat));
  NOR3_X1   g532(.A1(new_n686), .A2(G50gat), .A3(new_n517), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n725), .A2(new_n545), .A3(new_n726), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(G50gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g536(.A(new_n626), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n738), .A2(new_n259), .A3(new_n254), .A4(new_n661), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n574), .B2(new_n544), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n665), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT104), .B(G57gat), .Z(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1332gat));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n740), .B(new_n541), .C1(new_n744), .C2(new_n590), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n590), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1333gat));
  NAND2_X1  g546(.A1(new_n740), .A2(new_n675), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n677), .A2(G71gat), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n748), .A2(G71gat), .B1(new_n740), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n545), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  INV_X1    g553(.A(new_n641), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n704), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n725), .A2(new_n738), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n345), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n700), .A2(KEYINPUT106), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(KEYINPUT107), .B2(KEYINPUT51), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n700), .B2(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT108), .Z(new_n769));
  NAND3_X1  g568(.A1(new_n738), .A2(new_n579), .A3(new_n665), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n758), .B1(new_n769), .B2(new_n771), .ZN(G1336gat));
  NOR2_X1   g571(.A1(new_n538), .A2(G92gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n766), .A2(new_n738), .A3(new_n767), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n538), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n580), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT110), .B1(new_n775), .B2(new_n580), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI221_X1 g578(.A(new_n774), .B1(KEYINPUT110), .B2(KEYINPUT52), .C1(new_n775), .C2(new_n580), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n757), .B2(new_n550), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n626), .A2(G99gat), .A3(new_n677), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n769), .B2(new_n783), .ZN(G1338gat));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n517), .A2(G106gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n766), .A2(new_n738), .A3(new_n767), .A4(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G106gat), .B1(new_n757), .B2(new_n517), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n787), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n789), .B(new_n791), .ZN(G1339gat));
  NOR2_X1   g591(.A1(new_n662), .A2(new_n704), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n605), .B2(new_n614), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n613), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n605), .A2(new_n614), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n618), .B1(new_n797), .B2(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n798), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n801), .A2(new_n619), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n690), .A2(new_n692), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n227), .A2(new_n230), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT112), .Z(new_n806));
  AOI21_X1  g605(.A(new_n228), .B1(new_n242), .B2(new_n243), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n250), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n254), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n803), .A2(new_n804), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n624), .B2(new_n625), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n801), .A2(new_n704), .A3(new_n619), .A4(new_n802), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n814), .B2(new_n804), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n793), .B1(new_n815), .B2(new_n641), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT113), .B1(new_n816), .B2(new_n545), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n716), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n816), .A2(KEYINPUT113), .A3(new_n545), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n538), .A2(new_n665), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n261), .ZN(new_n824));
  NOR4_X1   g623(.A1(new_n816), .A2(new_n345), .A3(new_n541), .A4(new_n518), .ZN(new_n825));
  AOI21_X1  g624(.A(G113gat), .B1(new_n259), .B2(new_n254), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT114), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(G1340gat));
  OAI21_X1  g628(.A(G120gat), .B1(new_n823), .B2(new_n626), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n626), .A2(G120gat), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n823), .B2(new_n641), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n825), .A2(new_n282), .A3(new_n755), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1342gat));
  NAND3_X1  g636(.A1(new_n825), .A2(new_n284), .A3(new_n660), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT116), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n823), .B2(new_n699), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n841), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n517), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n801), .A2(new_n619), .A3(new_n802), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n812), .B1(new_n851), .B2(new_n261), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n699), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n755), .B1(new_n853), .B2(new_n811), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n854), .B2(new_n793), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT119), .B(new_n858), .C1(new_n816), .C2(new_n517), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n804), .B1(new_n812), .B2(new_n813), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n851), .A2(new_n693), .A3(new_n809), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n641), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n793), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n517), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n858), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT120), .B(new_n850), .C1(new_n854), .C2(new_n793), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n857), .A2(new_n859), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n675), .A2(new_n821), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n704), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n550), .A2(new_n545), .A3(new_n538), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n345), .B(new_n873), .C1(new_n863), .C2(new_n864), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n261), .A2(G141gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n848), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n848), .ZN(new_n878));
  INV_X1    g677(.A(new_n261), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n869), .A2(new_n879), .A3(new_n870), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n880), .B2(G141gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n847), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n881), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n871), .A2(G141gat), .B1(new_n874), .B2(new_n875), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n883), .B(KEYINPUT121), .C1(new_n848), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n885), .ZN(G1344gat));
  AND2_X1   g685(.A1(new_n271), .A2(new_n272), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n874), .A2(new_n887), .A3(new_n738), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT122), .Z(new_n889));
  NAND2_X1  g688(.A1(new_n803), .A2(new_n660), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n809), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n853), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n894), .A2(new_n641), .B1(new_n261), .B2(new_n663), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n849), .B1(new_n895), .B2(new_n517), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n865), .A2(new_n866), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n738), .B1(new_n870), .B2(KEYINPUT123), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(KEYINPUT123), .B2(new_n870), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n869), .A2(new_n870), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n887), .B1(new_n903), .B2(new_n738), .ZN(new_n904));
  OAI221_X1 g703(.A(new_n889), .B1(new_n901), .B2(new_n902), .C1(new_n904), .C2(KEYINPUT59), .ZN(G1345gat));
  INV_X1    g704(.A(G155gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n874), .A2(new_n906), .A3(new_n755), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n903), .A2(new_n755), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n906), .ZN(G1346gat));
  AOI21_X1  g708(.A(G162gat), .B1(new_n874), .B2(new_n660), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n804), .A2(G162gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n903), .B2(new_n911), .ZN(G1347gat));
  NOR4_X1   g711(.A1(new_n816), .A2(new_n665), .A3(new_n538), .A4(new_n518), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n348), .A3(new_n704), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT125), .ZN(new_n915));
  INV_X1    g714(.A(new_n820), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n538), .A2(new_n665), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n916), .A2(new_n261), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n919), .B2(new_n348), .ZN(G1348gat));
  AOI21_X1  g719(.A(G176gat), .B1(new_n913), .B2(new_n738), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n916), .A2(new_n918), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n626), .B1(new_n381), .B2(new_n382), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1349gat));
  NAND3_X1  g723(.A1(new_n913), .A2(new_n387), .A3(new_n755), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n916), .A2(new_n641), .A3(new_n918), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n357), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(new_n925), .C1(new_n926), .C2(new_n357), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n355), .A3(new_n804), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n922), .A2(new_n660), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(G190gat), .ZN(new_n935));
  AOI211_X1 g734(.A(KEYINPUT61), .B(new_n355), .C1(new_n922), .C2(new_n660), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1351gat));
  XNOR2_X1  g736(.A(KEYINPUT126), .B(G197gat), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n918), .A2(new_n675), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n896), .B2(new_n897), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n941), .B2(new_n879), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n550), .A2(new_n545), .A3(new_n541), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n816), .A2(new_n665), .A3(new_n943), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(new_n704), .A3(new_n938), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n942), .A2(KEYINPUT127), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT127), .B1(new_n942), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(new_n941), .ZN(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n949), .B2(new_n626), .ZN(new_n950));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n951), .A3(new_n738), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n944), .A2(new_n411), .A3(new_n755), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n941), .A2(new_n755), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n949), .B2(new_n699), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n412), .A3(new_n804), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


