//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G134), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(KEYINPUT11), .A3(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n191), .A2(new_n187), .A3(KEYINPUT11), .A4(G134), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n196), .B2(KEYINPUT11), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT11), .B1(new_n187), .B2(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT66), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n193), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n193), .B2(new_n200), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(KEYINPUT78), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G101), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n207), .A2(new_n210), .A3(new_n214), .A4(new_n211), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n217), .A3(G101), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n222), .A2(KEYINPUT64), .A3(G146), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT64), .B1(new_n222), .B2(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G128), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(KEYINPUT65), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n222), .A2(G146), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n220), .B2(G143), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n222), .A2(KEYINPUT64), .A3(G146), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n229), .B1(new_n234), .B2(new_n226), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n222), .A2(G146), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT0), .A3(G128), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n209), .A2(G104), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n206), .A2(G107), .ZN(new_n242));
  OAI21_X1  g056(.A(G101), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n215), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(KEYINPUT76), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(G143), .B2(new_n220), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n237), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n221), .A2(new_n236), .A3(new_n248), .A4(G128), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n244), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT10), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n219), .A2(new_n240), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n215), .A2(new_n243), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT77), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n249), .A2(new_n245), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n253), .B1(new_n234), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(KEYINPUT10), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n205), .A2(new_n257), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n257), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n190), .A2(new_n192), .ZN(new_n267));
  INV_X1    g081(.A(new_n188), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n198), .B(new_n194), .ZN(new_n270));
  OAI21_X1  g084(.A(G131), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n193), .A2(new_n200), .A3(new_n201), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(G227), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n276), .B(new_n278), .Z(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n282));
  OR3_X1    g096(.A1(new_n263), .A2(new_n244), .A3(KEYINPUT80), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n263), .A2(new_n244), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(new_n255), .A3(KEYINPUT80), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT12), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT12), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n282), .A2(new_n285), .A3(new_n288), .A4(new_n283), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n265), .A2(new_n287), .A3(new_n279), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  OR2_X1    g106(.A1(KEYINPUT82), .A2(G469), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT82), .A2(G469), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n287), .A2(new_n289), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n273), .B(KEYINPUT78), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n266), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n265), .A2(new_n287), .A3(KEYINPUT81), .A4(new_n289), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n280), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n299), .A2(new_n280), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n274), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n295), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT9), .B(G234), .Z(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G475), .ZN(new_n312));
  XNOR2_X1  g126(.A(G113), .B(G122), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(new_n206), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT87), .ZN(new_n315));
  INV_X1    g129(.A(G237), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT68), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G237), .ZN(new_n319));
  AOI21_X1  g133(.A(G953), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(G143), .B1(new_n320), .B2(G214), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(G143), .A3(G214), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n201), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n323), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n325), .A2(G131), .A3(new_n321), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n315), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(KEYINPUT72), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G125), .A3(G140), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n330), .A2(G140), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT73), .B1(new_n335), .B2(new_n328), .ZN(new_n336));
  AND4_X1   g150(.A1(KEYINPUT73), .A2(new_n328), .A3(new_n329), .A4(G125), .ZN(new_n337));
  NOR4_X1   g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .A4(new_n220), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G131), .B1(new_n325), .B2(new_n321), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n322), .A2(new_n201), .A3(new_n323), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT87), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n333), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT19), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(KEYINPUT19), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n220), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n327), .A2(new_n339), .A3(new_n342), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n322), .A2(new_n323), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT18), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n350), .A2(new_n201), .A3(KEYINPUT86), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n351), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n345), .A2(new_n220), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n220), .B2(new_n343), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n314), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n324), .A2(KEYINPUT17), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G146), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n338), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n340), .A2(new_n341), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n358), .B(new_n361), .C1(new_n362), .C2(KEYINPUT17), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n363), .A2(new_n356), .A3(new_n314), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n312), .B(new_n292), .C1(new_n357), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT88), .B1(new_n357), .B2(new_n364), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n365), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n314), .B1(new_n363), .B2(new_n356), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT89), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n364), .A2(KEYINPUT89), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n373), .B(new_n292), .C1(new_n374), .C2(new_n372), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n369), .A2(new_n371), .B1(new_n375), .B2(G475), .ZN(new_n376));
  XOR2_X1   g190(.A(G116), .B(G119), .Z(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT2), .B(G113), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n216), .A3(new_n218), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n381));
  INV_X1    g195(.A(G119), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G116), .ZN(new_n383));
  OAI211_X1 g197(.A(G113), .B(new_n383), .C1(new_n377), .C2(new_n381), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n377), .B2(new_n378), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n380), .B1(new_n260), .B2(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(G110), .B(G122), .Z(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n387), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n389), .B(new_n380), .C1(new_n260), .C2(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n228), .A2(new_n235), .A3(G125), .A4(new_n238), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n263), .A2(new_n330), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G224), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G953), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n394), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n386), .A2(new_n399), .A3(new_n387), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n393), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n390), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n385), .B(new_n258), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n387), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT84), .B1(new_n409), .B2(KEYINPUT7), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n409), .A2(KEYINPUT84), .A3(KEYINPUT7), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n404), .B(new_n408), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n401), .A2(new_n412), .A3(new_n292), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n414), .B(KEYINPUT85), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G214), .B1(G237), .B2(G902), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n401), .A2(new_n412), .A3(new_n292), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(G234), .A2(G237), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(G952), .A3(new_n277), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT21), .B(G898), .Z(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(G902), .A3(G953), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n422), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G478), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT15), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(G116), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n437), .A2(new_n209), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT14), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n436), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT90), .B(new_n436), .C1(new_n434), .C2(new_n439), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n442), .B(new_n443), .C1(KEYINPUT14), .C2(new_n435), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n438), .B1(new_n444), .B2(G107), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n245), .A2(G143), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n222), .A2(G128), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n195), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(KEYINPUT13), .B2(new_n446), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(KEYINPUT13), .B2(new_n446), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G134), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n195), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n437), .A2(new_n209), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n453), .B(new_n454), .C1(new_n438), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G217), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n309), .A2(new_n458), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n450), .A2(new_n456), .A3(new_n459), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT91), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI211_X1 g279(.A(KEYINPUT91), .B(G902), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n432), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n432), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n376), .A2(new_n430), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n311), .A2(KEYINPUT92), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n245), .A2(G119), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n245), .A2(G119), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT23), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT71), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G110), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT71), .ZN(new_n479));
  OAI211_X1 g293(.A(G119), .B(new_n245), .C1(new_n479), .C2(KEYINPUT23), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n481), .A2(KEYINPUT74), .ZN(new_n482));
  INV_X1    g296(.A(new_n475), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n474), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT24), .B(G110), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(KEYINPUT74), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n339), .A3(new_n354), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n477), .A2(new_n480), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G110), .ZN(new_n491));
  OAI221_X1 g305(.A(new_n491), .B1(new_n484), .B2(new_n485), .C1(new_n360), .C2(new_n338), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT22), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(G137), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n492), .A3(new_n496), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n458), .B1(G234), .B2(new_n292), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n292), .A3(new_n499), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT25), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n498), .A2(new_n507), .A3(new_n292), .A4(new_n499), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT32), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n239), .B1(new_n271), .B2(new_n272), .ZN(new_n515));
  OAI21_X1  g329(.A(G131), .B1(new_n196), .B2(new_n188), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n272), .A2(new_n516), .A3(new_n263), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT30), .B(new_n517), .C1(new_n204), .C2(new_n239), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n379), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n379), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(new_n517), .C1(new_n204), .C2(new_n239), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n320), .A2(G210), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n526), .B(new_n527), .Z(new_n528));
  AND4_X1   g342(.A1(new_n513), .A2(new_n521), .A3(new_n523), .A4(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n379), .B1(new_n515), .B2(new_n518), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n523), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n523), .A2(new_n531), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n530), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n513), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n529), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n512), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n521), .A2(new_n523), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n530), .ZN(new_n544));
  INV_X1    g358(.A(new_n523), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n273), .A2(new_n240), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n522), .B1(new_n546), .B2(new_n517), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT28), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n528), .A3(new_n534), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n548), .A2(KEYINPUT29), .A3(new_n528), .A4(new_n534), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n292), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n513), .B2(new_n536), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT32), .B(new_n540), .C1(new_n556), .C2(new_n529), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n542), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n542), .A2(new_n554), .A3(KEYINPUT70), .A4(new_n557), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n511), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT92), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n307), .A2(new_n310), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(new_n471), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n473), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  NOR2_X1   g381(.A1(new_n539), .A2(new_n541), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n292), .B1(new_n556), .B2(new_n529), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(G472), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n511), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n310), .A4(new_n307), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n461), .A2(new_n462), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n462), .B2(KEYINPUT93), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n461), .B(new_n462), .C1(KEYINPUT93), .C2(new_n574), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n431), .B(G902), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n463), .B(new_n464), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n431), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n376), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n430), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT34), .B(G104), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT94), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n583), .B(new_n585), .ZN(G6));
  INV_X1    g400(.A(new_n572), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n365), .A2(KEYINPUT95), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n365), .A2(KEYINPUT95), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n367), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n375), .A2(G475), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n467), .A2(new_n469), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(KEYINPUT20), .A3(new_n589), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n429), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n587), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G107), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G9));
  NAND2_X1  g413(.A1(new_n569), .A2(G472), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n539), .B2(new_n541), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n493), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n502), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n509), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT96), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n509), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n473), .A2(new_n565), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT37), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n478), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G12));
  NAND2_X1  g430(.A1(new_n560), .A2(new_n561), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n421), .B(KEYINPUT99), .Z(new_n618));
  INV_X1    g432(.A(G900), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n426), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n595), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n307), .A2(new_n609), .A3(new_n310), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n617), .A2(new_n621), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  XNOR2_X1  g440(.A(new_n620), .B(KEYINPUT39), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n311), .A2(KEYINPUT40), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n564), .B2(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n418), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n605), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n376), .A2(new_n470), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n530), .B1(new_n521), .B2(new_n523), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n532), .A2(new_n523), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n292), .B1(new_n638), .B2(new_n528), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n542), .A2(new_n557), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n417), .A2(new_n419), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT38), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n636), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n632), .A2(new_n634), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT100), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n632), .A2(new_n648), .A3(new_n645), .A4(new_n634), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n222), .ZN(G45));
  NOR3_X1   g465(.A1(new_n376), .A2(new_n580), .A3(new_n620), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n617), .A2(new_n623), .A3(new_n624), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G146), .ZN(G48));
  INV_X1    g468(.A(new_n582), .ZN(new_n655));
  INV_X1    g469(.A(new_n297), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n303), .A2(new_n656), .B1(new_n275), .B2(new_n280), .ZN(new_n657));
  OAI21_X1  g471(.A(G469), .B1(new_n657), .B2(G902), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n658), .A2(new_n295), .A3(new_n310), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n562), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  NAND4_X1  g476(.A1(new_n617), .A2(new_n596), .A3(new_n571), .A4(new_n659), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G116), .ZN(G18));
  AND3_X1   g478(.A1(new_n659), .A2(new_n623), .A3(new_n428), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n609), .A2(new_n376), .A3(new_n470), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n617), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n617), .A2(KEYINPUT101), .A3(new_n665), .A4(new_n666), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G119), .ZN(G21));
  XNOR2_X1  g486(.A(new_n540), .B(KEYINPUT102), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n537), .A2(new_n538), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n556), .A2(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n673), .B1(new_n678), .B2(new_n529), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n571), .A3(new_n659), .A4(new_n600), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n680), .A2(new_n429), .A3(new_n636), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n433), .ZN(G24));
  AND2_X1   g496(.A1(new_n679), .A2(new_n600), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n659), .A2(new_n623), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n605), .A3(new_n684), .A4(new_n652), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G125), .ZN(G27));
  AOI21_X1  g500(.A(new_n633), .B1(new_n417), .B2(new_n419), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n307), .A2(new_n310), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n376), .A2(new_n580), .A3(KEYINPUT42), .A4(new_n620), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n562), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n652), .A2(new_n558), .A3(new_n571), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT42), .B1(new_n692), .B2(new_n688), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n201), .ZN(G33));
  NAND4_X1  g509(.A1(new_n617), .A2(new_n621), .A3(new_n571), .A4(new_n689), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G134), .ZN(G36));
  NAND2_X1  g511(.A1(new_n302), .A2(new_n304), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n302), .A2(KEYINPUT45), .A3(new_n304), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(G469), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(G469), .A2(G902), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n702), .A2(KEYINPUT46), .A3(new_n703), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n295), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n310), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT104), .B1(new_n709), .B2(new_n627), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n711), .A3(new_n310), .A4(new_n628), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n713));
  INV_X1    g527(.A(new_n580), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n376), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n714), .A2(KEYINPUT43), .A3(new_n376), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n601), .A3(new_n605), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n710), .A2(new_n712), .B1(new_n713), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n713), .ZN(new_n722));
  INV_X1    g536(.A(new_n687), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G137), .ZN(G39));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n708), .A2(new_n727), .A3(new_n310), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n727), .B1(new_n708), .B2(new_n310), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n617), .A2(new_n571), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n652), .A2(new_n687), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n730), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n733), .A3(new_n728), .A4(new_n735), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G140), .ZN(G42));
  INV_X1    g555(.A(new_n715), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n571), .A3(new_n310), .A4(new_n418), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT106), .Z(new_n744));
  NAND2_X1  g558(.A1(new_n658), .A2(new_n295), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(KEYINPUT49), .Z(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n642), .A3(new_n644), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT107), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n729), .A2(new_n730), .B1(new_n310), .B2(new_n745), .ZN(new_n750));
  INV_X1    g564(.A(new_n618), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n717), .B2(new_n718), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n752), .A2(new_n571), .A3(new_n683), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(new_n687), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n633), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n683), .A2(new_n571), .A3(new_n644), .A4(new_n659), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n756), .A2(new_n757), .A3(new_n755), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n750), .A2(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n659), .A2(new_n687), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n571), .A2(new_n422), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n761), .A2(new_n762), .A3(new_n641), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n376), .A3(new_n580), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n761), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n752), .A2(new_n605), .A3(new_n683), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n765), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n749), .B1(new_n760), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n759), .A2(new_n758), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n749), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n770), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n745), .A2(new_n310), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT112), .Z(new_n779));
  OAI21_X1  g593(.A(new_n754), .B1(new_n731), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n759), .A2(new_n775), .A3(new_n758), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n763), .A2(new_n581), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n277), .A2(G952), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n752), .A2(new_n558), .A3(new_n571), .A4(new_n767), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT48), .Z(new_n787));
  AOI211_X1 g601(.A(new_n785), .B(new_n787), .C1(new_n684), .C2(new_n753), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n783), .A2(KEYINPUT115), .A3(new_n784), .A4(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n777), .A2(new_n781), .A3(new_n780), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n788), .B(new_n784), .C1(new_n790), .C2(new_n772), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n376), .A2(new_n470), .A3(new_n622), .A4(new_n605), .ZN(new_n796));
  INV_X1    g610(.A(new_n620), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n311), .A2(new_n796), .A3(new_n797), .A4(new_n641), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n625), .A2(new_n653), .A3(new_n685), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n622), .B1(new_n560), .B2(new_n561), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n801), .B(new_n624), .C1(new_n621), .C2(new_n652), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n685), .A4(new_n798), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n800), .A2(KEYINPUT110), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT109), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n562), .B(new_n659), .C1(new_n655), .C2(new_n596), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n473), .B(new_n565), .C1(new_n562), .C2(new_n611), .ZN(new_n813));
  INV_X1    g627(.A(new_n357), .ZN(new_n814));
  INV_X1    g628(.A(new_n364), .ZN(new_n815));
  AOI21_X1  g629(.A(G475), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n816), .A2(new_n292), .B1(new_n368), .B2(new_n367), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n370), .A2(new_n365), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n592), .B(new_n593), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT108), .B1(new_n819), .B2(new_n429), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT108), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n376), .A2(new_n430), .A3(new_n821), .A4(new_n593), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n572), .B1(new_n823), .B2(new_n582), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n681), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n671), .A2(new_n812), .A3(new_n813), .A4(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n600), .A2(new_n652), .A3(new_n605), .A4(new_n679), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n591), .A2(new_n592), .A3(new_n594), .A4(new_n797), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n564), .A2(new_n828), .A3(new_n610), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n470), .A2(new_n687), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n560), .B2(new_n561), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n827), .A2(new_n689), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n691), .A3(new_n693), .A4(new_n696), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n811), .B1(new_n826), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n660), .A2(new_n663), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n669), .B2(new_n670), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n691), .A2(new_n696), .A3(new_n693), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n831), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n683), .A2(new_n689), .A3(new_n605), .A4(new_n652), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n820), .A2(new_n822), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n587), .B1(new_n842), .B2(new_n655), .ZN(new_n843));
  INV_X1    g657(.A(new_n681), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n813), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n836), .A2(new_n841), .A3(new_n845), .A4(KEYINPUT109), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n809), .A2(new_n810), .A3(new_n834), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n805), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n834), .A2(new_n848), .A3(new_n846), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n850), .A3(KEYINPUT54), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n810), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n826), .A2(new_n833), .A3(new_n810), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n809), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n795), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n834), .A2(new_n810), .A3(new_n846), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n858), .A2(new_n809), .B1(new_n849), .B2(KEYINPUT53), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT111), .B1(new_n859), .B2(KEYINPUT54), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n794), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(G952), .A2(G953), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n748), .B1(new_n861), .B2(new_n862), .ZN(G75));
  AOI22_X1  g677(.A1(new_n849), .A2(new_n810), .B1(new_n809), .B2(new_n854), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n292), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n415), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n391), .A2(new_n400), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(new_n398), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT55), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n866), .A2(KEYINPUT116), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n277), .A2(G952), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT56), .B1(new_n865), .B2(new_n415), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n870), .B1(new_n875), .B2(KEYINPUT116), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(KEYINPUT116), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(G51));
  INV_X1    g692(.A(new_n856), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n864), .A2(new_n853), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n703), .B(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n291), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n864), .A2(new_n292), .A3(new_n702), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n872), .B1(new_n883), .B2(new_n884), .ZN(G54));
  AOI21_X1  g699(.A(KEYINPUT117), .B1(KEYINPUT58), .B2(G475), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(KEYINPUT117), .A2(KEYINPUT58), .A3(G475), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n865), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n357), .A2(new_n364), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n873), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n889), .A2(new_n894), .A3(new_n890), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n891), .B1(new_n893), .B2(new_n895), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT59), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n857), .B2(new_n860), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n576), .A2(new_n577), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n898), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n852), .A2(new_n855), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n856), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n903), .B1(new_n907), .B2(new_n872), .ZN(new_n908));
  OAI211_X1 g722(.A(KEYINPUT119), .B(new_n873), .C1(new_n881), .C2(new_n904), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n902), .A2(new_n908), .A3(new_n909), .ZN(G63));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n912));
  INV_X1    g726(.A(new_n500), .ZN(new_n913));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n864), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n912), .B1(new_n916), .B2(new_n873), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n915), .ZN(new_n919));
  INV_X1    g733(.A(new_n603), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n912), .B1(new_n920), .B2(KEYINPUT121), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n905), .A2(new_n919), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n911), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n917), .A2(new_n925), .A3(KEYINPUT61), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n926), .ZN(G66));
  NAND2_X1  g741(.A1(new_n826), .A2(new_n277), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT122), .Z(new_n929));
  OAI21_X1  g743(.A(G953), .B1(new_n424), .B2(new_n395), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n868), .B1(G898), .B2(new_n277), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  AOI21_X1  g747(.A(new_n277), .B1(G227), .B2(G900), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT126), .Z(new_n936));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n625), .A2(new_n653), .A3(new_n685), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n647), .A2(new_n649), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n819), .B1(new_n376), .B2(new_n580), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n562), .A2(new_n628), .A3(new_n689), .A4(new_n943), .ZN(new_n944));
  AOI22_X1  g758(.A1(new_n721), .A2(new_n724), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(new_n942), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n941), .A2(new_n740), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n277), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n519), .A2(new_n520), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n346), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n937), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n950), .ZN(new_n952));
  AOI211_X1 g766(.A(KEYINPUT124), .B(new_n952), .C1(new_n947), .C2(new_n277), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(G900), .A2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n938), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n721), .B2(new_n724), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n558), .A2(new_n571), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n710), .B2(new_n712), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n636), .A2(new_n622), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n837), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n740), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n955), .B(new_n952), .C1(new_n962), .C2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n936), .B1(new_n954), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n936), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n951), .A2(new_n953), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G72));
  XNOR2_X1  g784(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n971), .B(new_n972), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n947), .B2(new_n826), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n637), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n962), .B2(new_n826), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n543), .A2(new_n528), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n873), .A3(new_n979), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n978), .A2(new_n637), .A3(new_n973), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n859), .B2(new_n981), .ZN(G57));
endmodule


