//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(G116), .B(G119), .Z(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(G134), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .A3(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n198), .A2(G134), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n208), .B1(G134), .B2(new_n198), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n201), .A2(KEYINPUT11), .A3(G137), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n205), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n211), .A3(KEYINPUT67), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n220), .B(G146), .C1(new_n216), .C2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n216), .A2(new_n218), .A3(G143), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n225), .A2(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(KEYINPUT68), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n214), .A2(new_n215), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n219), .A2(new_n221), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G143), .B(G146), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT0), .B(G128), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n211), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT11), .B1(new_n201), .B2(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n208), .A2(new_n198), .A3(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n205), .B1(new_n238), .B2(new_n207), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n234), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n228), .A2(KEYINPUT30), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n204), .A2(new_n225), .A3(new_n211), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n204), .A2(new_n225), .A3(new_n211), .A4(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n196), .B(new_n241), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n196), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n228), .A2(new_n240), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n193), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n246), .A2(new_n196), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n228), .A2(KEYINPUT28), .A3(new_n240), .A4(new_n252), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n193), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n188), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n253), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n228), .A2(KEYINPUT71), .A3(new_n240), .A4(new_n252), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n228), .A2(new_n240), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n196), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT28), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n261), .A2(new_n255), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n257), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G472), .B1(new_n263), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n253), .A2(new_n193), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n251), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n260), .A2(new_n261), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n246), .A2(new_n248), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n241), .A2(new_n196), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n282), .B(new_n275), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT69), .B1(new_n251), .B2(new_n276), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n281), .B1(new_n290), .B2(KEYINPUT31), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n274), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n251), .A2(new_n276), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n282), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n251), .A2(KEYINPUT69), .A3(new_n276), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(KEYINPUT31), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n281), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT32), .B1(new_n303), .B2(new_n292), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n294), .B1(new_n291), .B2(new_n293), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n272), .B(new_n188), .C1(new_n254), .C2(new_n262), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n303), .A2(new_n295), .B1(new_n307), .B2(G472), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT72), .ZN(new_n309));
  INV_X1    g123(.A(G217), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(G234), .B2(new_n188), .ZN(new_n311));
  XOR2_X1   g125(.A(G119), .B(G128), .Z(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT24), .B(G110), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT23), .B1(new_n216), .B2(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n216), .A2(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT73), .B1(new_n318), .B2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(G128), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(KEYINPUT23), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n314), .B1(new_n322), .B2(G110), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G146), .ZN(new_n330));
  XNOR2_X1  g144(.A(G125), .B(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n218), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n322), .A2(G110), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n312), .A2(new_n313), .ZN(new_n335));
  AOI21_X1  g149(.A(G146), .B1(new_n328), .B2(new_n329), .ZN(new_n336));
  INV_X1    g150(.A(new_n330), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G137), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n339), .B(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n333), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n333), .B2(new_n338), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT25), .B1(new_n345), .B2(new_n188), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n347));
  NOR4_X1   g161(.A1(new_n343), .A2(new_n344), .A3(new_n347), .A4(G902), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n311), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n311), .A2(G902), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n305), .A2(new_n309), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n235), .A2(new_n239), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n357), .B2(G107), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G104), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(G107), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n358), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n357), .A2(G107), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n360), .A2(G104), .ZN(new_n366));
  OAI21_X1  g180(.A(G101), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n223), .A2(new_n224), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(KEYINPUT75), .B2(new_n222), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n231), .A2(new_n371), .A3(new_n217), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n225), .B1(new_n364), .B2(new_n367), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n356), .B(KEYINPUT12), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n373), .B2(new_n374), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n222), .A2(KEYINPUT75), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n378), .A2(new_n372), .A3(new_n223), .A4(new_n224), .ZN(new_n379));
  INV_X1    g193(.A(new_n368), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n368), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(KEYINPUT76), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n356), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n375), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n373), .A2(KEYINPUT10), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n358), .A2(new_n361), .A3(new_n363), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G101), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n394), .A3(G101), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n234), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n227), .A4(new_n380), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n390), .A2(new_n396), .A3(new_n355), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n340), .A2(G227), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(KEYINPUT74), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n390), .A2(new_n396), .A3(new_n397), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n356), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n399), .A2(new_n403), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n354), .B(G469), .C1(new_n409), .C2(G902), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n408), .ZN(new_n411));
  INV_X1    g225(.A(new_n398), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n384), .A2(new_n386), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT77), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n412), .B1(new_n416), .B2(new_n375), .ZN(new_n417));
  OAI211_X1 g231(.A(G469), .B(new_n411), .C1(new_n417), .C2(new_n404), .ZN(new_n418));
  NAND2_X1  g232(.A1(G469), .A2(G902), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(KEYINPUT78), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G469), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n405), .B1(new_n416), .B2(new_n375), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n404), .B1(new_n408), .B2(new_n398), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n421), .B(new_n188), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n410), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT9), .B(G234), .ZN(new_n426));
  OAI21_X1  g240(.A(G221), .B1(new_n426), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(G475), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n340), .A3(G214), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n220), .ZN(new_n431));
  AOI21_X1  g245(.A(G143), .B1(new_n189), .B2(G214), .ZN(new_n432));
  OAI21_X1  g246(.A(G131), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n220), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n205), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT83), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT17), .B(G131), .C1(new_n431), .C2(new_n432), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT82), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n436), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT17), .A4(G131), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n337), .A2(new_n336), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n433), .A2(new_n447), .A3(new_n434), .A4(new_n437), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n439), .A2(new_n445), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n357), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n331), .B(new_n218), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n331), .A2(new_n218), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n332), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT18), .A2(G131), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n442), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n442), .A2(new_n458), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n449), .A2(new_n451), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n449), .A2(new_n462), .ZN(new_n465));
  INV_X1    g279(.A(new_n451), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(KEYINPUT84), .B(new_n451), .C1(new_n449), .C2(new_n462), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n428), .B1(new_n469), .B2(new_n188), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT19), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n331), .B1(KEYINPUT81), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(new_n331), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n330), .B1(new_n475), .B2(G146), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n433), .B2(new_n437), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n453), .A2(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n463), .ZN(new_n480));
  NOR2_X1   g294(.A1(G475), .A2(G902), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n481), .ZN(new_n483));
  AOI211_X1 g297(.A(KEYINPUT20), .B(new_n483), .C1(new_n479), .C2(new_n463), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n470), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G478), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT87), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n426), .A2(new_n310), .A3(G953), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G116), .ZN(new_n497));
  INV_X1    g311(.A(G116), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G122), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(G107), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n216), .B2(G143), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n220), .A2(KEYINPUT85), .A3(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n216), .A2(G143), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n201), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT13), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(KEYINPUT13), .A3(new_n504), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n506), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G134), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT86), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n515), .A3(G134), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n508), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n505), .A2(new_n506), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n201), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n360), .B1(new_n497), .B2(KEYINPUT14), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(new_n500), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n495), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n512), .A2(new_n515), .A3(G134), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n515), .B1(new_n512), .B2(G134), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n507), .B(new_n501), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n522), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n494), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n493), .B1(new_n529), .B2(new_n188), .ZN(new_n530));
  AOI211_X1 g344(.A(G902), .B(new_n492), .C1(new_n523), .C2(new_n528), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n486), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n196), .A2(new_n393), .A3(new_n395), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n194), .A2(new_n195), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT5), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n318), .A3(G116), .ZN(new_n537));
  OAI211_X1 g351(.A(G113), .B(new_n537), .C1(new_n194), .C2(new_n536), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n380), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G110), .B(G122), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n539), .A3(new_n541), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(KEYINPUT6), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n225), .A2(new_n326), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n326), .B2(new_n233), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n340), .A2(G224), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT79), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n547), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT6), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n540), .A2(new_n551), .A3(new_n542), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n538), .A2(new_n535), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n368), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n539), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n541), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n558), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n546), .B(new_n560), .C1(new_n326), .C2(new_n233), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n556), .A2(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(G902), .B1(new_n562), .B2(new_n544), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G210), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n553), .A2(new_n565), .A3(new_n563), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G214), .B1(G237), .B2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(G234), .A2(G237), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(G952), .A3(new_n340), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(G902), .A3(G953), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT88), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT21), .B(G898), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n570), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n533), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n425), .A2(new_n427), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n353), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n362), .ZN(G3));
  AOI21_X1  g398(.A(new_n293), .B1(new_n301), .B2(new_n302), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n303), .A2(new_n188), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(G472), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n587), .A2(new_n425), .A3(new_n352), .A4(new_n427), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT89), .Z(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT91), .A2(KEYINPUT33), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n517), .A2(new_n522), .A3(new_n495), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n494), .B1(new_n526), .B2(new_n527), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(KEYINPUT91), .A2(KEYINPUT33), .ZN(new_n594));
  INV_X1    g408(.A(new_n590), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n523), .B(new_n528), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n487), .A2(G902), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n529), .A2(new_n188), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n487), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n486), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n569), .B2(new_n570), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n553), .A2(new_n565), .A3(new_n563), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n565), .B1(new_n553), .B2(new_n563), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n604), .B(new_n570), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n579), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n589), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  AOI22_X1  g428(.A1(KEYINPUT83), .A2(new_n438), .B1(new_n441), .B2(new_n444), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n446), .A2(new_n448), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n478), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT84), .B1(new_n617), .B2(new_n451), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n465), .A2(new_n464), .A3(new_n466), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n618), .A2(new_n619), .B1(new_n451), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g434(.A(G475), .B1(new_n620), .B2(G902), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n479), .A2(new_n463), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT20), .B1(new_n622), .B2(new_n483), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n480), .A2(new_n471), .A3(new_n481), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n532), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n611), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n589), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT92), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  INV_X1    g447(.A(KEYINPUT93), .ZN(new_n634));
  INV_X1    g448(.A(new_n342), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(KEYINPUT36), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n333), .A2(new_n636), .A3(new_n338), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n333), .B2(new_n338), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n634), .B1(new_n639), .B2(new_n351), .ZN(new_n640));
  INV_X1    g454(.A(new_n351), .ZN(new_n641));
  NOR4_X1   g455(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT93), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n349), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n587), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n582), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT37), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  INV_X1    g462(.A(new_n427), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n423), .B1(new_n389), .B2(new_n406), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(G469), .A3(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n418), .A2(new_n419), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n354), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n649), .B1(new_n653), .B2(new_n420), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n606), .A2(new_n607), .ZN(new_n655));
  INV_X1    g469(.A(new_n570), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT90), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n608), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n575), .A2(G900), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n572), .B(KEYINPUT94), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND4_X1   g475(.A1(new_n658), .A2(new_n627), .A3(new_n644), .A4(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n654), .A2(new_n305), .A3(new_n309), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XNOR2_X1  g478(.A(new_n661), .B(KEYINPUT39), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n654), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n299), .A2(new_n300), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n261), .B2(new_n269), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n669), .B2(G902), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n303), .A2(new_n295), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n306), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n655), .B(KEYINPUT38), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n486), .A2(new_n532), .ZN(new_n675));
  INV_X1    g489(.A(new_n644), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n570), .A3(new_n676), .ZN(new_n677));
  OR3_X1    g491(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n667), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n220), .ZN(G45));
  NOR2_X1   g495(.A1(new_n605), .A2(new_n609), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n601), .B(new_n661), .C1(new_n470), .C2(new_n485), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n676), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n654), .A2(new_n305), .A3(new_n309), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT95), .B(G146), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G48));
  NAND2_X1  g501(.A1(new_n611), .A2(new_n603), .ZN(new_n688));
  OAI21_X1  g502(.A(G469), .B1(new_n650), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n424), .A3(new_n427), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT96), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT96), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n689), .A2(new_n424), .A3(new_n692), .A4(new_n427), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n353), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT41), .B(G113), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  AND2_X1   g511(.A1(new_n691), .A2(new_n693), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n305), .A3(new_n309), .A4(new_n352), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT97), .B1(new_n699), .B2(new_n628), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n305), .A2(new_n309), .A3(new_n352), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT97), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n629), .A4(new_n698), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND4_X1   g519(.A1(new_n532), .A2(new_n644), .A3(new_n621), .A4(new_n625), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n427), .A3(new_n424), .A4(new_n689), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n610), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n305), .A3(new_n309), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NAND2_X1  g524(.A1(new_n270), .A2(new_n257), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n261), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n301), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT98), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT98), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n301), .A2(new_n715), .A3(new_n712), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n279), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n292), .ZN(new_n718));
  INV_X1    g532(.A(G472), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n303), .B2(new_n188), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n352), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT99), .B1(new_n486), .B2(new_n532), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT99), .ZN(new_n724));
  OAI221_X1 g538(.A(new_n724), .B1(new_n530), .B2(new_n531), .C1(new_n470), .C2(new_n485), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n723), .A2(new_n725), .B1(new_n657), .B2(new_n608), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(new_n579), .A3(new_n691), .A4(new_n693), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n496), .ZN(G24));
  AOI21_X1  g543(.A(new_n720), .B1(new_n717), .B2(new_n292), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n682), .A2(new_n690), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT100), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n626), .A2(new_n733), .A3(new_n601), .A4(new_n661), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n730), .A2(new_n644), .A3(new_n731), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  XOR2_X1   g551(.A(new_n419), .B(KEYINPUT101), .Z(new_n738));
  NAND3_X1  g552(.A1(new_n418), .A2(new_n424), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n649), .A2(new_n656), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n655), .A2(new_n740), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n732), .A2(new_n739), .A3(new_n734), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n306), .A2(new_n308), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n352), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n743), .B2(new_n352), .ZN(new_n746));
  OAI211_X1 g560(.A(KEYINPUT42), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n742), .A2(new_n305), .A3(new_n309), .A4(new_n352), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT102), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n748), .B2(new_n749), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n747), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND4_X1  g568(.A1(new_n739), .A2(new_n627), .A3(new_n661), .A4(new_n741), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n353), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n201), .ZN(G36));
  OR2_X1    g571(.A1(new_n409), .A2(KEYINPUT45), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n409), .A2(KEYINPUT45), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(G469), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT46), .B1(new_n760), .B2(new_n738), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n651), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(KEYINPUT46), .A3(new_n738), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n649), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n665), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT105), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n626), .A2(new_n602), .ZN(new_n767));
  NOR2_X1   g581(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n768));
  NAND2_X1  g582(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n767), .B2(new_n770), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(new_n644), .C1(new_n585), .C2(new_n720), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT44), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n655), .A2(new_n570), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT107), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n774), .A2(KEYINPUT108), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT108), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n766), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  XNOR2_X1  g594(.A(new_n764), .B(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n305), .A2(new_n309), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n683), .A2(new_n352), .A3(new_n775), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT109), .Z(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n736), .A2(new_n663), .ZN(new_n789));
  INV_X1    g603(.A(new_n661), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n644), .A2(new_n649), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n672), .A2(new_n726), .A3(new_n739), .A4(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n685), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT112), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n663), .A2(new_n736), .A3(new_n685), .A4(new_n792), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n788), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  INV_X1    g615(.A(new_n580), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n627), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n588), .A2(new_n803), .B1(new_n582), .B2(new_n645), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n603), .A2(new_n802), .ZN(new_n805));
  OAI22_X1  g619(.A1(new_n353), .A2(new_n582), .B1(new_n588), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n709), .B1(new_n722), .B2(new_n727), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n695), .A2(new_n809), .ZN(new_n810));
  OAI221_X1 g624(.A(KEYINPUT111), .B1(new_n588), .B2(new_n805), .C1(new_n353), .C2(new_n582), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n704), .A2(new_n808), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n730), .A2(new_n742), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n533), .A2(new_n790), .A3(new_n775), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n305), .A2(new_n309), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n654), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n756), .B1(new_n817), .B2(new_n644), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n753), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n812), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n800), .A2(new_n801), .A3(new_n820), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n704), .A2(new_n808), .A3(new_n811), .A4(new_n810), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n753), .A2(new_n818), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n789), .A2(new_n793), .A3(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n795), .A2(new_n796), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT52), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n798), .A2(new_n822), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(KEYINPUT113), .A3(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n828), .A3(KEYINPUT54), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n808), .A2(KEYINPUT53), .A3(new_n811), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n819), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n704), .A2(new_n810), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n800), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n827), .A2(new_n801), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT114), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n827), .A2(new_n842), .A3(new_n801), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n830), .A2(new_n833), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n772), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n660), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n690), .A2(new_n775), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n730), .A2(new_n644), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n673), .A2(new_n849), .A3(new_n352), .A4(new_n573), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n626), .A3(new_n601), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n722), .A2(new_n847), .A3(new_n660), .ZN(new_n856));
  INV_X1    g670(.A(new_n690), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n656), .A3(new_n674), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n853), .B(new_n855), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n689), .A2(new_n424), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n427), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n781), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n867), .A2(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n856), .A2(new_n776), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n867), .B2(KEYINPUT116), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n864), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n776), .A3(new_n856), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT51), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n851), .B1(new_n745), .B2(new_n746), .ZN(new_n874));
  NOR2_X1   g688(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n603), .ZN(new_n877));
  OAI211_X1 g691(.A(G952), .B(new_n340), .C1(new_n854), .C2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n856), .B2(new_n731), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n876), .B(new_n879), .C1(new_n874), .C2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n871), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n846), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n352), .A2(new_n740), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT110), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n674), .A3(new_n767), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(KEYINPUT49), .B2(new_n865), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(KEYINPUT49), .B2(new_n865), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n672), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n844), .A2(new_n188), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(G210), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n545), .A2(new_n552), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n550), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT55), .Z(new_n896));
  AND3_X1   g710(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n892), .B2(new_n893), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n340), .A2(G952), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G51));
  XOR2_X1   g714(.A(new_n650), .B(KEYINPUT118), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n800), .A2(new_n835), .A3(new_n838), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n827), .A2(new_n842), .A3(new_n801), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n842), .B1(new_n827), .B2(new_n801), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n845), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n738), .B(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n844), .A2(new_n188), .A3(new_n760), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n908), .B2(new_n909), .ZN(G54));
  INV_X1    g724(.A(new_n899), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n622), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n622), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n912), .A2(KEYINPUT119), .A3(new_n622), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n593), .A2(new_n596), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  OR2_X1    g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n911), .B1(new_n906), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n830), .A2(new_n833), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n844), .A2(new_n845), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n919), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT120), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n919), .C1(new_n846), .C2(new_n921), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n923), .B1(new_n928), .B2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT121), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n905), .A2(new_n639), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n905), .A2(KEYINPUT122), .A3(new_n639), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n345), .B1(new_n905), .B2(new_n934), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n899), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n939), .B2(new_n941), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  INV_X1    g759(.A(new_n577), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n340), .B1(new_n946), .B2(G224), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n812), .B2(new_n340), .ZN(new_n948));
  INV_X1    g762(.A(G898), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n894), .B1(new_n949), .B2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  NAND2_X1  g765(.A1(new_n789), .A2(new_n685), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n680), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n603), .A2(new_n627), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n775), .B1(new_n955), .B2(KEYINPUT124), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(KEYINPUT124), .B2(new_n955), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n957), .A2(new_n666), .A3(new_n353), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n954), .A2(new_n779), .A3(new_n786), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n340), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n286), .A2(new_n241), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(new_n475), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n766), .B(new_n726), .C1(new_n745), .C2(new_n746), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n756), .B(new_n952), .C1(new_n781), .C2(new_n785), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n779), .A3(new_n966), .A4(new_n753), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n967), .B2(G953), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n340), .B1(G227), .B2(G900), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT126), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n969), .B(new_n973), .Z(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  OAI211_X1 g790(.A(new_n829), .B(new_n976), .C1(new_n668), .C2(new_n254), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n967), .B2(new_n812), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n251), .A2(new_n253), .A3(new_n261), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n899), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n976), .B1(new_n959), .B2(new_n812), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n261), .B1(new_n251), .B2(new_n253), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n981), .B2(new_n983), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n977), .B(new_n980), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(G57));
endmodule


