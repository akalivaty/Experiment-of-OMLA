//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  XOR2_X1   g035(.A(KEYINPUT66), .B(G2105), .Z(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G137), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n460), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT66), .B(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  OAI221_X1 g045(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n458), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(KEYINPUT67), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n462), .A2(new_n463), .A3(new_n472), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT67), .B1(new_n475), .B2(new_n476), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n461), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n478), .A2(new_n487), .A3(new_n461), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n482), .B1(new_n489), .B2(G124), .ZN(G162));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n479), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G138), .B1(new_n462), .B2(new_n463), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n461), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n475), .A2(new_n476), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n497), .A2(new_n466), .A3(new_n498), .A4(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(G75), .A2(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(G651), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n504), .B2(new_n505), .ZN(new_n511));
  AND2_X1   g086(.A1(G50), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND2_X1  g090(.A1(new_n509), .A2(KEYINPUT69), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n516), .A2(G543), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT70), .B(G89), .Z(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(new_n509), .B1(G63), .B2(G651), .ZN(new_n526));
  INV_X1    g101(.A(new_n505), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n524), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n522), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n504), .A2(new_n505), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n516), .A2(G52), .A3(G543), .A4(new_n520), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(new_n509), .A3(G90), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g118(.A(KEYINPUT72), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n532), .A2(new_n509), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n529), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(G81), .A2(new_n547), .B1(new_n550), .B2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n521), .A2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n516), .A2(G53), .A3(G543), .A4(new_n520), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n503), .B1(new_n509), .B2(KEYINPUT69), .ZN(new_n563));
  XOR2_X1   g138(.A(KEYINPUT73), .B(KEYINPUT9), .Z(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(G53), .A3(new_n520), .A4(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n532), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n568), .B2(new_n534), .ZN(new_n569));
  OAI21_X1  g144(.A(G65), .B1(new_n527), .B2(new_n528), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(KEYINPUT74), .A3(G651), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n569), .A2(new_n573), .B1(G91), .B2(new_n547), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n566), .A2(new_n574), .ZN(G299));
  AND2_X1   g150(.A1(new_n543), .A2(new_n544), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  NAND3_X1  g152(.A1(new_n563), .A2(G49), .A3(new_n520), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n532), .A2(new_n509), .A3(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n529), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G48), .A2(G543), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(G651), .B1(new_n509), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n547), .A2(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n547), .A2(G85), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n516), .A2(G543), .A3(new_n520), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n589), .B1(new_n534), .B2(new_n590), .C1(new_n591), .C2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(new_n592), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n546), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n529), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n600), .A2(new_n603), .B1(G651), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT76), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n595), .B1(new_n594), .B2(new_n609), .ZN(G284));
  XOR2_X1   g185(.A(G284), .B(KEYINPUT77), .Z(G321));
  NAND2_X1  g186(.A1(G299), .A2(new_n594), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n594), .B2(G168), .ZN(G280));
  XOR2_X1   g188(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n615), .B2(G860), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT79), .Z(G148));
  OAI21_X1  g192(.A(KEYINPUT80), .B1(new_n554), .B2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n609), .A2(new_n615), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  MUX2_X1   g195(.A(KEYINPUT80), .B(new_n618), .S(new_n620), .Z(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g197(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n623));
  NOR3_X1   g198(.A1(new_n474), .A2(new_n458), .A3(G2105), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n623), .B(new_n624), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n489), .A2(G123), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n461), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(G2105), .B1(new_n473), .B2(new_n477), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n628), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT84), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(G14), .A3(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n627), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n637), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(KEYINPUT85), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1971), .ZN(new_n695));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n695), .B1(new_n698), .B2(KEYINPUT86), .ZN(new_n699));
  NOR2_X1   g274(.A1(G16), .A2(G23), .ZN(new_n700));
  AND3_X1   g275(.A1(new_n563), .A2(G49), .A3(new_n520), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n579), .A2(new_n580), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT87), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n578), .A2(new_n704), .A3(new_n579), .A4(new_n580), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n699), .B(new_n709), .C1(KEYINPUT86), .C2(new_n698), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n712));
  NOR2_X1   g287(.A1(G25), .A2(G29), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n633), .A2(G131), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(G107), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n461), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n714), .B(new_n717), .C1(new_n489), .C2(G119), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n713), .B1(new_n718), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G24), .B(G290), .S(G16), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1986), .ZN(new_n724));
  INV_X1    g299(.A(new_n719), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n720), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n711), .A2(new_n712), .A3(new_n722), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(KEYINPUT88), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n727), .B(new_n729), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n692), .A2(G4), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n609), .B2(new_n692), .ZN(new_n732));
  INV_X1    g307(.A(G1348), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n692), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n554), .B2(new_n692), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G1341), .Z(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G26), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT28), .Z(new_n740));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n741));
  INV_X1    g316(.A(G140), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n480), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n633), .A2(KEYINPUT89), .A3(G140), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(G2104), .B(new_n746), .C1(new_n466), .C2(G116), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT90), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(KEYINPUT90), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n487), .B1(new_n478), .B2(new_n461), .ZN(new_n751));
  AOI211_X1 g326(.A(KEYINPUT68), .B(new_n466), .C1(new_n473), .C2(new_n477), .ZN(new_n752));
  OAI21_X1  g327(.A(G128), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n745), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n740), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2067), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n734), .A2(new_n737), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT91), .ZN(new_n758));
  OAI21_X1  g333(.A(G129), .B1(new_n751), .B2(new_n752), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(KEYINPUT95), .B(G129), .C1(new_n751), .C2(new_n752), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n633), .A2(G141), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT26), .Z(new_n766));
  INV_X1    g341(.A(G105), .ZN(new_n767));
  INV_X1    g342(.A(new_n459), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n764), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(KEYINPUT96), .B1(new_n763), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n772), .B(new_n769), .C1(new_n761), .C2(new_n762), .ZN(new_n773));
  OAI21_X1  g348(.A(G29), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G32), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(G29), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G5), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G171), .B2(G16), .ZN(new_n780));
  INV_X1    g355(.A(G1961), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G168), .A2(new_n692), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n692), .B2(G21), .ZN(new_n784));
  INV_X1    g359(.A(G1966), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT24), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n738), .B1(new_n787), .B2(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n787), .B2(G34), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G160), .B2(G29), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G2084), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(G28), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n738), .B1(new_n792), .B2(G28), .ZN(new_n794));
  AND2_X1   g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  NOR2_X1   g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n790), .B2(G2084), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n636), .A2(G29), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n786), .A2(new_n791), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n633), .A2(G139), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n497), .A2(G127), .ZN(new_n805));
  AND2_X1   g380(.A1(G115), .A2(G2104), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n461), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  NOR2_X1   g385(.A1(G29), .A2(G33), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT92), .Z(new_n812));
  AOI22_X1  g387(.A1(new_n810), .A2(new_n812), .B1(KEYINPUT94), .B2(G2072), .ZN(new_n813));
  NOR2_X1   g388(.A1(KEYINPUT94), .A2(G2072), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G27), .A2(G29), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G164), .B2(G29), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G2078), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(G2078), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n818), .B(new_n819), .C1(new_n784), .C2(new_n785), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n800), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n692), .A2(G20), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT23), .Z(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G299), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT98), .B(G1956), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G35), .ZN(new_n827));
  OR3_X1    g402(.A1(new_n827), .A2(KEYINPUT97), .A3(G29), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT97), .B1(new_n827), .B2(G29), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n828), .B(new_n829), .C1(G162), .C2(new_n738), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT29), .B(G2090), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  AND4_X1   g407(.A1(new_n782), .A2(new_n821), .A3(new_n826), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n758), .A2(new_n778), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n730), .A2(new_n834), .ZN(G311));
  INV_X1    g410(.A(G311), .ZN(G150));
  NAND2_X1  g411(.A1(new_n609), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT99), .B(G93), .Z(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n529), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n547), .A2(new_n839), .B1(new_n842), .B2(G651), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n521), .A2(G55), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n553), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n551), .A2(new_n843), .A3(new_n552), .A4(new_n844), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n838), .B(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n850), .A2(new_n851), .A3(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n845), .A2(G860), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  XOR2_X1   g430(.A(new_n635), .B(G160), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n496), .A2(new_n499), .ZN(new_n859));
  INV_X1    g434(.A(new_n494), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n489), .A2(G128), .B1(new_n749), .B2(new_n748), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n745), .ZN(new_n863));
  AND4_X1   g438(.A1(new_n861), .A2(new_n745), .A3(new_n750), .A4(new_n753), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n771), .A2(new_n773), .A3(KEYINPUT100), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT95), .B1(new_n489), .B2(G129), .ZN(new_n868));
  INV_X1    g443(.A(G129), .ZN(new_n869));
  AOI211_X1 g444(.A(new_n760), .B(new_n869), .C1(new_n486), .C2(new_n488), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n770), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n772), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n769), .B1(new_n761), .B2(new_n762), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT96), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n867), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n865), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT100), .B1(new_n771), .B2(new_n773), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n867), .A3(new_n874), .ZN(new_n878));
  INV_X1    g453(.A(new_n865), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n809), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n873), .B1(new_n863), .B2(new_n864), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n754), .A2(G164), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n862), .A2(new_n861), .A3(new_n745), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n871), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT101), .B1(new_n886), .B2(new_n808), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n888));
  AOI211_X1 g463(.A(new_n888), .B(new_n809), .C1(new_n882), .C2(new_n885), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n891));
  INV_X1    g466(.A(G118), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n461), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G142), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n480), .A2(KEYINPUT102), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT102), .B1(new_n480), .B2(new_n894), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n489), .A2(new_n898), .A3(G130), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n489), .B2(G130), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n718), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n625), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n718), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n881), .A2(new_n890), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n881), .B2(new_n890), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n858), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n908), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n879), .B1(new_n877), .B2(new_n878), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n913), .A2(new_n914), .A3(new_n808), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n809), .B1(new_n882), .B2(new_n885), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT101), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n912), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n881), .A2(new_n890), .A3(new_n908), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n857), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n911), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n911), .A2(new_n920), .A3(KEYINPUT104), .A4(new_n921), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n924), .A2(KEYINPUT40), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT40), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(G395));
  NAND2_X1  g503(.A1(new_n846), .A2(new_n847), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT105), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n619), .B(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n608), .A2(G299), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n608), .A2(G299), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT41), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n932), .B2(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n933), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n608), .A2(G299), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n931), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n706), .B(G305), .Z(new_n947));
  XNOR2_X1  g522(.A(G290), .B(G166), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n946), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(G868), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n845), .A2(new_n594), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(G295));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n954), .ZN(G331));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g532(.A1(G301), .A2(new_n929), .ZN(new_n958));
  NAND2_X1  g533(.A1(G171), .A2(new_n848), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(G168), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(G171), .A2(new_n848), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n929), .B1(new_n544), .B2(new_n543), .ZN(new_n962));
  OAI21_X1  g537(.A(G286), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n963), .A3(new_n934), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n938), .B1(new_n963), .B2(new_n960), .ZN(new_n966));
  OAI211_X1 g541(.A(KEYINPUT107), .B(new_n949), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n960), .A2(new_n963), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n939), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n947), .B(new_n948), .Z(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n964), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n921), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n969), .B2(new_n964), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(KEYINPUT107), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT108), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n921), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n949), .B1(new_n965), .B2(new_n966), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n977), .A2(new_n980), .A3(new_n981), .A4(new_n967), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n957), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n976), .B2(new_n973), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n976), .C2(new_n973), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n977), .A2(new_n980), .A3(new_n957), .A4(new_n967), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n985), .A2(new_n993), .ZN(G397));
  NAND3_X1  g569(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n995));
  INV_X1    g570(.A(G125), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n475), .B2(new_n476), .ZN(new_n997));
  INV_X1    g572(.A(new_n468), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n461), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G137), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n475), .B2(new_n476), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n466), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n999), .A2(G40), .A3(new_n460), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n995), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(G164), .B2(G1384), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n754), .B(G2067), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n871), .ZN(new_n1012));
  INV_X1    g587(.A(G1996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT127), .B(KEYINPUT46), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1012), .B(new_n1016), .C1(new_n1014), .C2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT47), .Z(new_n1019));
  INV_X1    g594(.A(new_n1010), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1011), .A2(new_n1010), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT111), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1013), .B1(new_n771), .B2(new_n773), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(G1996), .B2(new_n873), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n718), .A2(new_n720), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n754), .A2(G2067), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n718), .A2(new_n720), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1010), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  OR3_X1    g607(.A1(new_n1020), .A2(G1986), .A3(G290), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT48), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1019), .B(new_n1029), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n566), .A2(new_n574), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n547), .A2(G91), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT74), .B1(new_n572), .B2(G651), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n567), .B(new_n534), .C1(new_n570), .C2(new_n571), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n562), .A2(new_n565), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT57), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  INV_X1    g620(.A(G1384), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n861), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1005), .A4(new_n995), .ZN(new_n1049));
  INV_X1    g624(.A(G1956), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n1046), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT56), .B(G2072), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1006), .A2(new_n1009), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1044), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G164), .A2(G1384), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n995), .A3(new_n1005), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G2067), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n733), .B2(new_n1049), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(new_n608), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1044), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1055), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n608), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1059), .B1(KEYINPUT60), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(KEYINPUT60), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1044), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT61), .B1(new_n1067), .B2(new_n1055), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1044), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1061), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1057), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1052), .A2(new_n1009), .A3(new_n1005), .A4(new_n995), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(G1996), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT59), .B1(new_n1078), .B2(new_n553), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1080), .A3(new_n554), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1068), .A2(new_n1073), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1066), .B1(new_n1082), .B2(KEYINPUT119), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(KEYINPUT119), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1062), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1076), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1088), .A2(G1971), .B1(G2090), .B2(new_n1049), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n1090));
  INV_X1    g665(.A(G8), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n508), .B2(new_n513), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT112), .A3(KEYINPUT55), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT112), .B1(new_n1092), .B2(KEYINPUT55), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1095), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT113), .A3(new_n1093), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1092), .A2(KEYINPUT55), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1089), .A2(G8), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT114), .B(G8), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1089), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n703), .A2(G1976), .A3(new_n705), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT115), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n703), .A2(new_n1108), .A3(G1976), .A4(new_n705), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n1057), .A3(new_n1103), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT52), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1057), .A2(new_n1103), .ZN(new_n1112));
  INV_X1    g687(.A(G1976), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT52), .B1(G288), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(new_n1106), .A3(new_n1109), .A4(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT116), .B(G86), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n547), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n586), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G1981), .ZN(new_n1119));
  INV_X1    g694(.A(G1981), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n586), .A2(new_n1120), .A3(new_n587), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT49), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(KEYINPUT49), .A3(new_n1121), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1112), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1111), .A2(new_n1115), .A3(new_n1126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1101), .A2(new_n1104), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1052), .A2(new_n1009), .ZN(new_n1130));
  INV_X1    g705(.A(G2078), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT53), .B(new_n1131), .C1(new_n1003), .C2(KEYINPUT124), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(KEYINPUT124), .B2(new_n1003), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1130), .A2(new_n1133), .B1(new_n1049), .B2(new_n781), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1076), .B2(G2078), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1129), .B(G301), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1133), .A2(new_n1130), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1049), .A2(new_n781), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT125), .B1(new_n1140), .B2(G171), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1009), .A2(new_n1005), .A3(new_n995), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1009), .A2(new_n1145), .A3(new_n1005), .A4(new_n995), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1146), .A3(new_n1052), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1131), .A2(KEYINPUT53), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1139), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(G301), .A2(new_n1136), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT54), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1128), .B1(new_n1142), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1136), .B(new_n1139), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G171), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT123), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1153), .A2(new_n1156), .A3(G171), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1134), .A2(G301), .A3(new_n1136), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G168), .A2(new_n1102), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1143), .A2(KEYINPUT117), .B1(KEYINPUT45), .B2(new_n1056), .ZN(new_n1163));
  AOI21_X1  g738(.A(G1966), .B1(new_n1163), .B2(new_n1146), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1049), .A2(G2084), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1162), .A2(KEYINPUT51), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1147), .B2(new_n785), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1168), .B2(new_n1102), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(KEYINPUT121), .B(new_n1167), .C1(new_n1168), .C2(new_n1102), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n1173));
  OAI21_X1  g748(.A(G8), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1162), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1171), .B(new_n1172), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1166), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1087), .A2(new_n1161), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1126), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1121), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1112), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1089), .A2(G8), .A3(new_n1100), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(new_n1127), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1168), .A2(new_n1102), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1111), .A2(new_n1115), .A3(new_n1126), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1188), .A2(new_n1189), .A3(G168), .A4(new_n1186), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT118), .B1(new_n1190), .B2(new_n1104), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1101), .A2(new_n1127), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1104), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1168), .A2(G286), .A3(new_n1102), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1191), .A2(new_n1192), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1100), .B1(new_n1089), .B2(G8), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1190), .A2(new_n1192), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1187), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1181), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(KEYINPUT126), .B1(new_n1180), .B2(KEYINPUT62), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n1204));
  OAI211_X1 g779(.A(new_n1204), .B(new_n1166), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1206), .A2(new_n1128), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1180), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1202), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1010), .A2(G1986), .A3(G290), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1033), .A2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1213), .B(KEYINPUT110), .Z(new_n1214));
  NAND2_X1  g789(.A1(new_n1032), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1035), .B1(new_n1211), .B2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g791(.A1(new_n924), .A2(new_n925), .ZN(new_n1218));
  INV_X1    g792(.A(G319), .ZN(new_n1219));
  NOR4_X1   g793(.A1(G401), .A2(new_n1219), .A3(G227), .A4(G229), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n1218), .A2(new_n991), .A3(new_n1220), .ZN(G225));
  INV_X1    g795(.A(G225), .ZN(G308));
endmodule


