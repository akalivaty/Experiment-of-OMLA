//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  AOI22_X1  g0004(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n208));
  NAND4_X1  g0008(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT1), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n204), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n211), .B(new_n221), .C1(new_n220), .C2(new_n219), .ZN(G361));
  XOR2_X1   g0022(.A(G238), .B(G244), .Z(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(G226), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(G250), .B(G257), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n227), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G68), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(G50), .B(G58), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  INV_X1    g0039(.A(G33), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT3), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G33), .ZN(new_n243));
  AND2_X1   g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g0044(.A1(G222), .A2(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G223), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n248), .B(new_n249), .C1(G77), .C2(new_n244), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n249), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(G226), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G179), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g0062(.A(new_n262), .B(KEYINPUT69), .Z(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n264), .A2(new_n214), .ZN(new_n265));
  INV_X1    g0065(.A(G58), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT8), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(KEYINPUT8), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n240), .A2(G20), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n269), .A2(new_n270), .B1(G150), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G50), .A2(G58), .ZN(new_n273));
  INV_X1    g0073(.A(G68), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n215), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n265), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G1), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(G50), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n215), .A2(G1), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n278), .A2(new_n215), .A3(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n264), .A2(new_n214), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT67), .B1(new_n284), .B2(new_n285), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n283), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n282), .B1(new_n290), .B2(new_n281), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(KEYINPUT68), .B(new_n282), .C1(new_n290), .C2(new_n281), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n277), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n260), .A2(G169), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n263), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n260), .A2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n260), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n295), .B2(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n299), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  OAI211_X1 g0110(.A(G1), .B(G13), .C1(new_n240), .C2(new_n255), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n253), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(G274), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n310), .A2(new_n312), .B1(new_n313), .B2(new_n253), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n242), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G33), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(G226), .A2(G1698), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n241), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT78), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT78), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n318), .A2(new_n322), .A3(new_n241), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G87), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n318), .A2(G223), .A3(new_n246), .A4(new_n241), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n321), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n314), .B1(new_n326), .B2(new_n249), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n261), .B(new_n314), .C1(new_n326), .C2(new_n249), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n288), .A2(new_n289), .ZN(new_n332));
  INV_X1    g0132(.A(new_n283), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n269), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n269), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n332), .A2(new_n335), .B1(new_n284), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n241), .ZN(new_n339));
  AND2_X1   g0139(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n340));
  NOR2_X1   g0140(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n339), .B1(new_n342), .B2(G33), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT7), .B1(new_n343), .B2(G20), .ZN(new_n344));
  AOI21_X1  g0144(.A(G20), .B1(new_n318), .B2(new_n241), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(G68), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n266), .A2(new_n274), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G58), .A2(G68), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n271), .A2(G159), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n265), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n355));
  INV_X1    g0155(.A(KEYINPUT77), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(new_n240), .C1(new_n340), .C2(new_n341), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n346), .A2(G20), .ZN(new_n358));
  AOI21_X1  g0158(.A(G33), .B1(new_n316), .B2(new_n317), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n243), .A2(KEYINPUT77), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n346), .B1(new_n244), .B2(G20), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n274), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n351), .A2(new_n352), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n355), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n338), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT18), .B1(new_n331), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n326), .A2(new_n249), .ZN(new_n369));
  INV_X1    g0169(.A(new_n314), .ZN(new_n370));
  AOI21_X1  g0170(.A(G200), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g0171(.A(G190), .B(new_n314), .C1(new_n326), .C2(new_n249), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(G68), .B1(new_n345), .B2(new_n346), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n343), .A2(KEYINPUT7), .A3(G20), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n353), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n285), .ZN(new_n377));
  INV_X1    g0177(.A(new_n355), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n361), .A2(new_n362), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  INV_X1    g0180(.A(new_n364), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n337), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n368), .B1(new_n373), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n369), .A2(G179), .A3(new_n370), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n328), .B2(new_n327), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT18), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n369), .A2(new_n389), .A3(new_n370), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G200), .B2(new_n327), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n366), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n367), .A2(new_n384), .A3(new_n388), .A4(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT79), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  INV_X1    g0196(.A(G244), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n312), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G232), .A2(G1698), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n246), .A2(G238), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n244), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n241), .A2(new_n243), .ZN(new_n402));
  INV_X1    g0202(.A(G107), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n311), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI211_X1 g0204(.A(new_n254), .B(new_n398), .C1(new_n401), .C2(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n405), .A2(G169), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n286), .A2(G77), .A3(new_n333), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT15), .B(G87), .ZN(new_n408));
  INV_X1    g0208(.A(new_n270), .ZN(new_n409));
  INV_X1    g0209(.A(G77), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n408), .A2(new_n409), .B1(new_n215), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n271), .B2(new_n269), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n407), .B1(G77), .B2(new_n280), .C1(new_n412), .C2(new_n265), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n405), .A2(new_n261), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n406), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n405), .A2(new_n302), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n413), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(KEYINPUT70), .B1(G190), .B2(new_n405), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT70), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n417), .B2(new_n413), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n416), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n309), .A2(new_n395), .A3(new_n396), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G238), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n312), .B2(KEYINPUT71), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT71), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n258), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(G226), .A2(G1698), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n310), .B2(G1698), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n244), .A2(new_n430), .B1(G33), .B2(G97), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n431), .A2(new_n311), .B1(new_n253), .B2(new_n313), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT13), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n244), .A2(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n254), .B1(new_n436), .B2(new_n249), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT13), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n425), .A2(new_n427), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT72), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n433), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(KEYINPUT72), .B(KEYINPUT13), .C1(new_n428), .C2(new_n432), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(G200), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n284), .A2(new_n274), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT12), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n270), .A2(G77), .B1(G20), .B2(new_n274), .ZN(new_n447));
  INV_X1    g0247(.A(new_n271), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n281), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n286), .A2(G68), .A3(new_n333), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n446), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT73), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT11), .B1(new_n449), .B2(new_n285), .ZN(new_n454));
  OR3_X1    g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n452), .B2(new_n454), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n433), .A2(new_n440), .A3(G190), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n444), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n442), .A2(G169), .A3(new_n443), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT14), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT14), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n442), .A2(new_n463), .A3(G169), .A4(new_n443), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n433), .A2(new_n440), .A3(G179), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n457), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n468), .B(KEYINPUT74), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n423), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n318), .A2(new_n215), .A3(G68), .A4(new_n241), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT19), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n409), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n215), .B1(new_n435), .B2(new_n472), .ZN(new_n475));
  INV_X1    g0275(.A(G87), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(new_n473), .A3(new_n403), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n475), .A2(KEYINPUT83), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT83), .B1(new_n475), .B2(new_n477), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n471), .B(new_n474), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n475), .A2(new_n477), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n471), .A4(new_n474), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n481), .A2(new_n488), .A3(new_n285), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n408), .A2(new_n284), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT85), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n252), .A2(G33), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n265), .A2(new_n280), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n492), .A2(new_n494), .B1(G87), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G238), .A2(G1698), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n397), .B2(G1698), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n343), .A2(new_n500), .B1(G33), .B2(G116), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n311), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n256), .A2(G1), .ZN(new_n503));
  INV_X1    g0303(.A(G250), .ZN(new_n504));
  NOR4_X1   g0304(.A1(new_n249), .A2(KEYINPUT82), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n503), .A2(new_n504), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(new_n311), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n252), .A2(G45), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n505), .A2(new_n508), .B1(new_n313), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n302), .B1(new_n502), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n501), .A2(new_n311), .ZN(new_n512));
  INV_X1    g0312(.A(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(G190), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n489), .A2(new_n493), .A3(new_n490), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n493), .B1(new_n489), .B2(new_n490), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n516), .A2(new_n517), .B1(new_n408), .B2(new_n496), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n512), .A2(new_n261), .A3(new_n513), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n328), .B1(new_n502), .B2(new_n510), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n498), .A2(new_n515), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n318), .A2(new_n241), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n246), .A2(G244), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n526), .A2(new_n524), .B1(new_n504), .B2(new_n246), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n244), .A2(new_n528), .B1(G33), .B2(G283), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n311), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n249), .A2(new_n251), .ZN(new_n531));
  OR2_X1    g0331(.A1(KEYINPUT5), .A2(G41), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT5), .A2(G41), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n509), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT5), .B(G41), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n503), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n311), .ZN(new_n538));
  INV_X1    g0338(.A(G257), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n530), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n261), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n403), .B1(new_n361), .B2(new_n362), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n544), .A2(new_n473), .A3(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(G97), .B(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n215), .B1(new_n410), .B2(new_n448), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n285), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT80), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n280), .B2(G97), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n284), .A2(KEYINPUT80), .A3(new_n473), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n497), .A2(G97), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n328), .B1(new_n530), .B2(new_n540), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n542), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n530), .A2(new_n389), .A3(new_n540), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT81), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n549), .B(new_n553), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n540), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n527), .A2(new_n529), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(G190), .C1(new_n561), .C2(new_n311), .ZN(new_n562));
  OAI21_X1  g0362(.A(G200), .B1(new_n530), .B2(new_n540), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT81), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n556), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n215), .A2(G33), .A3(G116), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n403), .A2(G20), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(KEYINPUT23), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT86), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n567), .B2(KEYINPUT23), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n215), .A2(G87), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n318), .A2(new_n574), .A3(new_n241), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n573), .B1(new_n402), .B2(new_n572), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(new_n569), .A3(KEYINPUT23), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n571), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT24), .ZN(new_n579));
  INV_X1    g0379(.A(new_n577), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n580), .A2(new_n568), .A3(new_n570), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n575), .A4(new_n576), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n265), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT25), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n280), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n403), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n497), .A2(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G250), .A2(G1698), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n539), .B2(G1698), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n318), .A3(new_n241), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G294), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n311), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n537), .A2(G264), .A3(new_n311), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n389), .A3(new_n535), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n537), .A2(new_n313), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n598), .B1(G200), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n593), .A2(new_n594), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n249), .ZN(new_n604));
  INV_X1    g0404(.A(new_n596), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n535), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n261), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n600), .A2(new_n328), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(new_n584), .B2(new_n589), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G270), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n535), .B1(new_n538), .B2(new_n611), .ZN(new_n612));
  MUX2_X1   g0412(.A(G257), .B(G264), .S(G1698), .Z(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n318), .A3(new_n241), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n402), .A2(G303), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n311), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G190), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n284), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n496), .B2(new_n619), .ZN(new_n621));
  NAND2_X1  g0421(.A1(G33), .A2(G283), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n622), .B(new_n215), .C1(G33), .C2(new_n473), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(G20), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n285), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT20), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n626), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n621), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n618), .B(new_n630), .C1(new_n302), .C2(new_n617), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  OAI21_X1  g0432(.A(G169), .B1(new_n612), .B2(new_n616), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(new_n630), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n286), .A2(G116), .A3(new_n495), .ZN(new_n635));
  INV_X1    g0435(.A(new_n629), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n620), .B(new_n635), .C1(new_n636), .C2(new_n627), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n617), .A2(new_n637), .A3(G179), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n534), .A2(new_n249), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(G270), .B1(new_n531), .B2(new_n534), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n614), .A2(new_n615), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n311), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n637), .A3(KEYINPUT21), .A4(G169), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n631), .A2(new_n634), .A3(new_n638), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n565), .A2(new_n610), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n470), .A2(new_n523), .A3(new_n645), .ZN(G372));
  NAND2_X1  g0446(.A1(new_n497), .A2(G87), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n647), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n648));
  INV_X1    g0448(.A(new_n556), .ZN(new_n649));
  INV_X1    g0449(.A(new_n408), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n492), .A2(new_n494), .B1(new_n650), .B2(new_n497), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n648), .B(new_n649), .C1(new_n651), .C2(new_n521), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n602), .B1(new_n559), .B2(new_n564), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n579), .A2(new_n583), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n285), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n606), .A2(G169), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n600), .A2(G179), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n656), .A2(new_n588), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n634), .A2(new_n643), .A3(new_n638), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n556), .B1(new_n654), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT26), .B1(new_n498), .B2(new_n515), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT87), .B1(new_n514), .B2(new_n328), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(KEYINPUT87), .B2(new_n521), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n518), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n470), .B1(new_n653), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n367), .A2(new_n388), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n466), .A2(new_n467), .B1(new_n459), .B2(new_n416), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n384), .A2(new_n392), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n306), .A2(new_n308), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n299), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(G369));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n644), .B(KEYINPUT88), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n279), .A2(new_n215), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(G213), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n679), .B1(new_n630), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n660), .A2(new_n637), .A3(new_n685), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT89), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n678), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n659), .A2(new_n685), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT90), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n602), .B(new_n609), .C1(new_n590), .C2(new_n686), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(KEYINPUT91), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT91), .B1(new_n694), .B2(new_n698), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n698), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n660), .A2(new_n686), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n659), .B2(new_n686), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n218), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  NOR4_X1   g0509(.A1(new_n709), .A2(new_n252), .A3(G116), .A4(new_n477), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n213), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  AOI22_X1  g0512(.A1(new_n498), .A2(new_n515), .B1(new_n666), .B2(new_n518), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT26), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n556), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n652), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(KEYINPUT26), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n649), .B1(new_n498), .B2(new_n515), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n654), .A2(new_n661), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n668), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT92), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT29), .A4(new_n686), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n667), .B1(new_n662), .B2(new_n663), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n685), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n713), .A2(new_n715), .B1(new_n652), .B2(new_n714), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT29), .B(new_n686), .C1(new_n731), .C2(new_n722), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT92), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n726), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n645), .A2(new_n523), .A3(new_n686), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n502), .A2(new_n510), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(new_n597), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n642), .A2(new_n261), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(KEYINPUT30), .A3(new_n738), .A4(new_n541), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n736), .A3(new_n541), .A4(new_n597), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n736), .A2(G179), .A3(new_n617), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n541), .A2(new_n600), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n685), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n740), .A2(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n686), .B1(new_n750), .B2(new_n739), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT31), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n735), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n734), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT93), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n712), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(new_n278), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT94), .B1(new_n758), .B2(G45), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n252), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n758), .A2(KEYINPUT94), .A3(G45), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n709), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n694), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n691), .A2(new_n678), .A3(new_n693), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n763), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n218), .A2(G355), .A3(new_n244), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n708), .A2(new_n343), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G45), .B2(new_n212), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n235), .A2(new_n256), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n768), .B1(G116), .B2(new_n218), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n278), .A2(new_n240), .A3(KEYINPUT95), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT95), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G13), .B2(G33), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n214), .B1(G20), .B2(new_n328), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n767), .B1(new_n772), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n779), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n215), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n389), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n403), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G159), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n785), .B1(new_n789), .B2(KEYINPUT32), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n389), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n215), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G97), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n215), .A2(new_n261), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n389), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n790), .B(new_n794), .C1(new_n281), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n796), .A2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n801), .A2(new_n274), .B1(new_n789), .B2(KEYINPUT32), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n476), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n799), .A2(new_n802), .A3(new_n402), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n795), .A2(G190), .A3(new_n302), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n795), .A2(new_n786), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n806), .A2(new_n266), .B1(new_n807), .B2(new_n410), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT96), .Z(new_n809));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n402), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT97), .Z(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT33), .B(G317), .Z(new_n813));
  INV_X1    g0613(.A(G326), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n801), .A2(new_n813), .B1(new_n798), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n788), .A2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n817), .B2(new_n807), .C1(new_n818), .C2(new_n806), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n792), .A2(new_n820), .B1(new_n784), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n815), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n805), .A2(new_n809), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n778), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n781), .B1(new_n782), .B2(new_n824), .C1(new_n690), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n766), .A2(new_n826), .ZN(G396));
  NOR2_X1   g0627(.A1(new_n415), .A2(new_n685), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n413), .A2(new_n685), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n419), .B2(new_n421), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n829), .B1(new_n831), .B2(new_n416), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n686), .B(new_n833), .C1(new_n669), .C2(new_n653), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT99), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n832), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n836), .B2(new_n729), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n763), .B1(new_n837), .B2(new_n754), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n754), .B2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n776), .A2(new_n779), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n767), .B1(new_n410), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n806), .ZN(new_n842));
  INV_X1    g0642(.A(new_n807), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n842), .A2(G143), .B1(new_n843), .B2(G159), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n844), .B1(new_n798), .B2(new_n845), .C1(new_n846), .C2(new_n801), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT34), .ZN(new_n848));
  INV_X1    g0648(.A(new_n784), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(G68), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n850), .B1(new_n281), .B2(new_n803), .C1(new_n266), .C2(new_n792), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n525), .B(new_n851), .C1(G132), .C2(new_n788), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n800), .A2(G283), .B1(new_n843), .B2(G116), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n810), .B2(new_n798), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT98), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n402), .B1(new_n787), .B2(new_n817), .C1(new_n806), .C2(new_n820), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n794), .B1(new_n403), .B2(new_n803), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(G87), .C2(new_n849), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n848), .A2(new_n852), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n841), .B1(new_n782), .B2(new_n859), .C1(new_n833), .C2(new_n777), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n839), .A2(new_n860), .ZN(G384));
  INV_X1    g0661(.A(new_n547), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n862), .A2(KEYINPUT35), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(KEYINPUT35), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(G116), .A3(new_n216), .A4(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT36), .Z(new_n866));
  OAI211_X1 g0666(.A(new_n213), .B(G77), .C1(new_n266), .C2(new_n274), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n281), .A2(G68), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n252), .B(G13), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT105), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n751), .B2(KEYINPUT31), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n747), .A2(KEYINPUT105), .A3(new_n748), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n735), .A2(new_n872), .A3(new_n873), .A4(new_n752), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n466), .A2(new_n467), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n467), .A2(new_n685), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n459), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n467), .B(new_n685), .C1(new_n466), .C2(new_n460), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n832), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n378), .B1(new_n348), .B2(new_n381), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n337), .B1(new_n377), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n385), .B(new_n683), .C1(new_n328), .C2(new_n327), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT100), .B(new_n337), .C1(new_n377), .C2(new_n883), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n391), .A2(new_n366), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(new_n683), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n383), .B1(new_n386), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n393), .A2(new_n893), .A3(new_n886), .A4(new_n888), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g0702(.A(KEYINPUT101), .B(KEYINPUT38), .C1(new_n897), .C2(new_n898), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n881), .B(new_n882), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n393), .A2(new_n383), .A3(new_n893), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT104), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n393), .A2(new_n908), .A3(new_n383), .A4(new_n893), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n373), .B2(new_n383), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n391), .A2(KEYINPUT102), .A3(new_n366), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n894), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n914), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT103), .B1(new_n914), .B2(KEYINPUT37), .ZN(new_n916));
  INV_X1    g0716(.A(new_n896), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n905), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n880), .B1(new_n919), .B2(new_n899), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n904), .B1(new_n920), .B2(new_n882), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n470), .A2(new_n874), .ZN(new_n923));
  OAI21_X1  g0723(.A(G330), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n875), .A2(new_n685), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT39), .B1(new_n902), .B2(new_n903), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n919), .A2(new_n929), .A3(new_n899), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n877), .A2(new_n878), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n834), .B2(new_n829), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n903), .B2(new_n902), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n671), .A2(new_n893), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n726), .A2(new_n470), .A3(new_n730), .A4(new_n733), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n676), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n925), .A2(new_n941), .B1(new_n252), .B2(new_n758), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n925), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n870), .B1(new_n942), .B2(new_n943), .ZN(G367));
  XNOR2_X1  g0744(.A(new_n762), .B(KEYINPUT109), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n701), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n699), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n686), .B1(new_n549), .B2(new_n553), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n565), .A2(new_n949), .B1(new_n556), .B2(new_n686), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n706), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n706), .A2(new_n950), .ZN(new_n953));
  XOR2_X1   g0753(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n948), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n702), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n698), .B(new_n704), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n694), .B(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n756), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(new_n756), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n709), .B(KEYINPUT41), .Z(new_n965));
  OAI21_X1  g0765(.A(new_n946), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n705), .A2(new_n950), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT42), .Z(new_n968));
  XOR2_X1   g0768(.A(new_n950), .B(KEYINPUT106), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n556), .B1(new_n969), .B2(new_n609), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n686), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n498), .A2(new_n686), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n667), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n713), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n974), .B2(new_n972), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n968), .A2(new_n971), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n976), .B(new_n977), .Z(new_n978));
  INV_X1    g0778(.A(new_n969), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n948), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT107), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n978), .A2(KEYINPUT107), .A3(new_n980), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n966), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n769), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n231), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n780), .B1(new_n218), .B2(new_n408), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n763), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n801), .A2(new_n820), .B1(new_n798), .B2(new_n817), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G107), .B2(new_n793), .ZN(new_n992));
  INV_X1    g0792(.A(new_n803), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(G116), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT46), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n806), .A2(new_n810), .B1(new_n807), .B2(new_n821), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G317), .B2(new_n788), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n784), .A2(new_n473), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(new_n343), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n992), .A2(new_n995), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G159), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n801), .A2(new_n1001), .B1(new_n274), .B2(new_n792), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G143), .B2(new_n797), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n806), .A2(new_n846), .B1(new_n807), .B2(new_n281), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n402), .B(new_n1004), .C1(G137), .C2(new_n788), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n993), .A2(G58), .B1(new_n849), .B2(G77), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT110), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n990), .B1(new_n1010), .B2(new_n779), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n825), .B2(new_n975), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n986), .A2(new_n1012), .ZN(G387));
  INV_X1    g0813(.A(new_n709), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n962), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n756), .B2(new_n961), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n780), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n769), .B1(new_n227), .B2(new_n256), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n477), .A2(G116), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n218), .A2(new_n244), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n269), .A2(new_n281), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT50), .Z(new_n1023));
  AOI21_X1  g0823(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1021), .A2(new_n1025), .B1(new_n403), .B2(new_n708), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n793), .A2(new_n650), .B1(new_n993), .B2(G77), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n1001), .B2(new_n798), .C1(new_n336), .C2(new_n801), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n842), .A2(G50), .B1(new_n843), .B2(G68), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n846), .B2(new_n787), .ZN(new_n1030));
  NOR4_X1   g0830(.A1(new_n1028), .A2(new_n525), .A3(new_n1030), .A4(new_n998), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n842), .A2(G317), .B1(new_n843), .B2(G303), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n798), .B2(new_n818), .C1(new_n817), .C2(new_n801), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n793), .A2(G283), .B1(new_n993), .B2(G294), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT49), .Z(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n525), .B1(new_n619), .B2(new_n784), .C1(new_n814), .C2(new_n787), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n1039), .B2(KEYINPUT111), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1031), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n763), .B1(new_n1017), .B2(new_n1026), .C1(new_n1043), .C2(new_n782), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n703), .B2(new_n778), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n961), .B2(new_n945), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1016), .A2(new_n1046), .ZN(G393));
  OR3_X1    g0847(.A1(new_n959), .A2(KEYINPUT114), .A3(new_n962), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT114), .B1(new_n959), .B2(new_n962), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n709), .A3(new_n963), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n946), .B1(new_n959), .B2(KEYINPUT112), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(KEYINPUT112), .B2(new_n959), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n987), .A2(new_n238), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n780), .B1(new_n473), .B2(new_n218), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n763), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n792), .A2(new_n410), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n801), .A2(new_n281), .B1(new_n803), .B2(new_n274), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G87), .C2(new_n849), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n798), .A2(new_n846), .B1(new_n1001), .B2(new_n806), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n269), .A2(new_n843), .B1(new_n788), .B2(G143), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n343), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G317), .A2(new_n797), .B1(new_n842), .B2(G311), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n993), .A2(G283), .B1(new_n788), .B2(G322), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n244), .B(new_n785), .C1(G294), .C2(new_n843), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G116), .A2(new_n793), .B1(new_n800), .B2(G303), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1063), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1056), .B1(new_n1072), .B2(new_n779), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n979), .B2(new_n825), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1051), .A2(new_n1053), .A3(new_n1074), .ZN(G390));
  NAND3_X1  g0875(.A1(new_n874), .A2(new_n879), .A3(G330), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n933), .B1(new_n754), .B2(new_n832), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT115), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n874), .A2(new_n879), .A3(new_n1079), .A4(G330), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n828), .B1(new_n729), .B2(new_n833), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n753), .A2(new_n932), .A3(G330), .A4(new_n833), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n831), .A2(new_n416), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n686), .B(new_n1086), .C1(new_n731), .C2(new_n722), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1085), .A2(new_n829), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n836), .A2(G330), .A3(new_n874), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n933), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n470), .A2(G330), .A3(new_n874), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n939), .A2(new_n676), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n927), .B1(new_n1082), .B2(new_n933), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n928), .A2(new_n930), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1087), .A2(new_n829), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n932), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n919), .A2(new_n899), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n927), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(new_n1101), .A3(new_n1085), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(KEYINPUT116), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1106), .B(new_n1103), .C1(new_n1097), .C2(new_n1101), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1095), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1103), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1106), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1081), .A2(new_n1083), .B1(new_n1090), .B2(new_n1088), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n939), .A2(new_n676), .A3(new_n1093), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1102), .A4(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1108), .A2(new_n1117), .A3(new_n709), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n928), .A2(new_n930), .A3(new_n776), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n801), .A2(new_n403), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1057), .B(new_n1121), .C1(G283), .C2(new_n797), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n804), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n806), .A2(new_n619), .B1(new_n807), .B2(new_n473), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n244), .B(new_n1124), .C1(G294), .C2(new_n788), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1122), .A2(new_n1123), .A3(new_n850), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n798), .A2(new_n1127), .B1(new_n784), .B2(new_n281), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n801), .A2(new_n845), .B1(new_n1001), .B2(new_n792), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n803), .A2(new_n846), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n402), .B1(new_n842), .B2(G132), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n843), .A2(new_n1136), .B1(new_n788), .B2(G125), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .A4(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n782), .B1(new_n1126), .B2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n767), .B(new_n1139), .C1(new_n336), .C2(new_n840), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1119), .A2(new_n945), .B1(new_n1120), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1118), .A2(new_n1141), .ZN(G378));
  NOR2_X1   g0942(.A1(new_n295), .A2(new_n683), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n309), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n309), .A2(new_n1144), .ZN(new_n1146));
  OR3_X1    g0946(.A1(new_n1145), .A2(new_n1146), .A3(KEYINPUT120), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT120), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1148), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(new_n777), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n343), .A2(G41), .ZN(new_n1154));
  AOI211_X1 g0954(.A(G50), .B(new_n1154), .C1(new_n240), .C2(new_n255), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n801), .A2(new_n473), .B1(new_n798), .B2(new_n619), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G58), .B2(new_n849), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n842), .A2(G107), .B1(new_n843), .B2(new_n650), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n821), .B2(new_n787), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n793), .A2(G68), .B1(new_n993), .B2(G77), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1157), .A2(new_n1154), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT58), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1155), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n800), .A2(G132), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n1127), .B2(new_n806), .C1(new_n845), .C2(new_n807), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G150), .A2(new_n793), .B1(new_n797), .B2(G125), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT118), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(new_n993), .C2(new_n1136), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT59), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1001), .B2(new_n784), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT119), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1164), .B1(new_n1163), .B2(new_n1162), .C1(new_n1171), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n779), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n840), .A2(new_n281), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n763), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1153), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n921), .A2(G330), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n938), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n921), .B(G330), .C1(new_n931), .C2(new_n937), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1152), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1183), .A2(new_n1184), .A3(new_n1152), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1181), .B1(new_n1189), .B2(new_n946), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1183), .A2(new_n1184), .A3(new_n1152), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1152), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1117), .A2(new_n1094), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1014), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1115), .B1(new_n1119), .B2(new_n1116), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1197), .B2(new_n1189), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1190), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(G375));
  INV_X1    g1000(.A(new_n965), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1095), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n945), .B(KEYINPUT121), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n933), .A2(new_n776), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n776), .A2(new_n779), .A3(G68), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n801), .A2(new_n619), .B1(new_n803), .B2(new_n473), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G294), .B2(new_n797), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n806), .A2(new_n821), .B1(new_n807), .B2(new_n403), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n244), .B(new_n1209), .C1(G303), .C2(new_n788), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n793), .A2(new_n650), .B1(new_n849), .B2(G77), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT122), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n806), .A2(new_n845), .B1(new_n807), .B2(new_n846), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G128), .B2(new_n788), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G50), .A2(new_n793), .B1(new_n797), .B2(G132), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n800), .A2(new_n1136), .B1(new_n993), .B2(G159), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n525), .B1(G58), .B2(new_n849), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1214), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n767), .B(new_n1206), .C1(new_n1222), .C2(new_n779), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1092), .A2(new_n1204), .B1(new_n1205), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1203), .A2(new_n1224), .ZN(G381));
  OR2_X1    g1025(.A1(G387), .A2(G390), .ZN(new_n1226));
  OR2_X1    g1026(.A1(G378), .A2(G381), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1228), .B(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OR4_X1    g1031(.A1(G375), .A2(new_n1226), .A3(new_n1227), .A4(new_n1231), .ZN(G407));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1199), .A2(new_n684), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  NOR2_X1   g1035(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1180), .B1(new_n1236), .B2(new_n945), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1187), .A2(KEYINPUT57), .A3(new_n1188), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n709), .B1(new_n1238), .B2(new_n1197), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1195), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G378), .B(new_n1237), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1105), .A2(new_n1107), .A3(new_n1095), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1201), .B1(new_n1242), .B2(new_n1115), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1204), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1189), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1233), .B1(new_n1245), .B2(new_n1180), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G343), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1202), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1014), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1114), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1224), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(G384), .A3(new_n1224), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1247), .A2(new_n1250), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1249), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(KEYINPUT62), .A3(new_n1260), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(KEYINPUT126), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1261), .A2(new_n1267), .A3(new_n1262), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1249), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1260), .B2(KEYINPUT124), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1269), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1271), .A2(new_n1274), .B1(KEYINPUT124), .B2(new_n1260), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n965), .B1(new_n1117), .B2(new_n1094), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1236), .B1(new_n1276), .B2(new_n1204), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G378), .B1(new_n1277), .B2(new_n1181), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G378), .B2(new_n1199), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1279), .B2(new_n1249), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT125), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1260), .A2(KEYINPUT124), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1274), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1269), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(KEYINPUT125), .B(new_n1281), .C1(new_n1264), .C2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1266), .B(new_n1268), .C1(new_n1282), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT127), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1281), .B1(new_n1264), .B2(new_n1286), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1287), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1268), .A4(new_n1266), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(G390), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1226), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1226), .B2(new_n1298), .ZN(new_n1300));
  OR2_X1    g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1290), .A2(new_n1296), .A3(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1261), .B(KEYINPUT63), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1281), .A3(new_n1280), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(G405));
  NAND2_X1  g1106(.A1(G375), .A2(new_n1233), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1241), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1272), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1303), .B(new_n1309), .ZN(G402));
endmodule


