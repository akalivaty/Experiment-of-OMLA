

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XOR2_X1 U322 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n290) );
  NOR2_X1 U323 ( .A1(n539), .A2(n538), .ZN(n564) );
  XNOR2_X1 U324 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U325 ( .A(KEYINPUT48), .B(n505), .Z(n536) );
  XOR2_X1 U326 ( .A(n340), .B(n339), .Z(n532) );
  XNOR2_X1 U327 ( .A(G15GAT), .B(G1GAT), .ZN(n291) );
  XNOR2_X1 U328 ( .A(n291), .B(KEYINPUT69), .ZN(n351) );
  XOR2_X1 U329 ( .A(G50GAT), .B(n351), .Z(n293) );
  NAND2_X1 U330 ( .A1(G229GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U331 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U332 ( .A(n294), .B(G36GAT), .Z(n302) );
  XOR2_X1 U333 ( .A(G141GAT), .B(G197GAT), .Z(n296) );
  XNOR2_X1 U334 ( .A(G169GAT), .B(G22GAT), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U336 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n298) );
  XNOR2_X1 U337 ( .A(G113GAT), .B(G8GAT), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U339 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U340 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U341 ( .A(n303), .B(KEYINPUT29), .Z(n307) );
  XOR2_X1 U342 ( .A(G29GAT), .B(G43GAT), .Z(n305) );
  XNOR2_X1 U343 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n304) );
  XNOR2_X1 U344 ( .A(n305), .B(n304), .ZN(n330) );
  XNOR2_X1 U345 ( .A(n330), .B(KEYINPUT30), .ZN(n306) );
  XNOR2_X1 U346 ( .A(n307), .B(n306), .ZN(n565) );
  XOR2_X1 U347 ( .A(KEYINPUT71), .B(KEYINPUT74), .Z(n309) );
  NAND2_X1 U348 ( .A1(G230GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U349 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U350 ( .A(n310), .B(KEYINPUT70), .Z(n315) );
  XNOR2_X1 U351 ( .A(G71GAT), .B(G57GAT), .ZN(n311) );
  XNOR2_X1 U352 ( .A(n311), .B(KEYINPUT13), .ZN(n350) );
  XOR2_X1 U353 ( .A(G64GAT), .B(G92GAT), .Z(n313) );
  XNOR2_X1 U354 ( .A(G176GAT), .B(G204GAT), .ZN(n312) );
  XNOR2_X1 U355 ( .A(n313), .B(n312), .ZN(n373) );
  XNOR2_X1 U356 ( .A(n350), .B(n373), .ZN(n314) );
  XNOR2_X1 U357 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U358 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n317) );
  XNOR2_X1 U359 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n316) );
  XNOR2_X1 U360 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U361 ( .A(n319), .B(n318), .Z(n323) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U363 ( .A(n320), .B(G148GAT), .ZN(n397) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(G85GAT), .ZN(n321) );
  XNOR2_X1 U365 ( .A(n290), .B(n321), .ZN(n329) );
  XNOR2_X1 U366 ( .A(n397), .B(n329), .ZN(n322) );
  XNOR2_X1 U367 ( .A(n323), .B(n322), .ZN(n569) );
  NOR2_X1 U368 ( .A1(n565), .A2(n569), .ZN(n452) );
  XOR2_X1 U369 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n357) );
  XOR2_X1 U370 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n325) );
  XNOR2_X1 U371 ( .A(KEYINPUT66), .B(KEYINPUT75), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n340) );
  XOR2_X1 U373 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n327) );
  NAND2_X1 U374 ( .A1(G232GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U376 ( .A(n328), .B(KEYINPUT64), .Z(n332) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U378 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U379 ( .A(G36GAT), .B(G190GAT), .Z(n358) );
  XOR2_X1 U380 ( .A(G92GAT), .B(n358), .Z(n334) );
  XOR2_X1 U381 ( .A(G50GAT), .B(G162GAT), .Z(n405) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(n405), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U384 ( .A(n336), .B(n335), .Z(n338) );
  XNOR2_X1 U385 ( .A(G134GAT), .B(G218GAT), .ZN(n337) );
  XNOR2_X1 U386 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U387 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n342) );
  XNOR2_X1 U388 ( .A(G127GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U389 ( .A(n342), .B(n341), .ZN(n355) );
  XNOR2_X1 U390 ( .A(G8GAT), .B(G183GAT), .ZN(n343) );
  XNOR2_X1 U391 ( .A(n343), .B(G211GAT), .ZN(n361) );
  XOR2_X1 U392 ( .A(G22GAT), .B(G155GAT), .Z(n404) );
  XOR2_X1 U393 ( .A(n361), .B(n404), .Z(n345) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U396 ( .A(G64GAT), .B(KEYINPUT76), .Z(n347) );
  XNOR2_X1 U397 ( .A(KEYINPUT14), .B(KEYINPUT77), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U399 ( .A(n349), .B(n348), .Z(n353) );
  XNOR2_X1 U400 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U401 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U402 ( .A(n355), .B(n354), .ZN(n574) );
  NAND2_X1 U403 ( .A1(n532), .A2(n574), .ZN(n356) );
  XNOR2_X1 U404 ( .A(n357), .B(n356), .ZN(n435) );
  XOR2_X1 U405 ( .A(KEYINPUT89), .B(n358), .Z(n360) );
  NAND2_X1 U406 ( .A1(G226GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U407 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U408 ( .A(n362), .B(n361), .Z(n371) );
  XOR2_X1 U409 ( .A(KEYINPUT81), .B(KEYINPUT18), .Z(n364) );
  XNOR2_X1 U410 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n363) );
  XNOR2_X1 U411 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U412 ( .A(n365), .B(KEYINPUT83), .Z(n367) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(KEYINPUT82), .ZN(n366) );
  XNOR2_X1 U414 ( .A(n367), .B(n366), .ZN(n377) );
  XOR2_X1 U415 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n369) );
  XNOR2_X1 U416 ( .A(G197GAT), .B(G218GAT), .ZN(n368) );
  XNOR2_X1 U417 ( .A(n369), .B(n368), .ZN(n398) );
  XNOR2_X1 U418 ( .A(n377), .B(n398), .ZN(n370) );
  XNOR2_X1 U419 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U420 ( .A(n373), .B(n372), .Z(n534) );
  XOR2_X1 U421 ( .A(G127GAT), .B(G134GAT), .Z(n375) );
  XNOR2_X1 U422 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n374) );
  XNOR2_X1 U423 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U424 ( .A(G113GAT), .B(n376), .Z(n418) );
  XNOR2_X1 U425 ( .A(n377), .B(n418), .ZN(n390) );
  XOR2_X1 U426 ( .A(G176GAT), .B(G190GAT), .Z(n379) );
  XNOR2_X1 U427 ( .A(G43GAT), .B(G99GAT), .ZN(n378) );
  XNOR2_X1 U428 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U429 ( .A(KEYINPUT84), .B(G71GAT), .Z(n381) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(G183GAT), .ZN(n380) );
  XNOR2_X1 U431 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U432 ( .A(n383), .B(n382), .Z(n388) );
  XOR2_X1 U433 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n385) );
  NAND2_X1 U434 ( .A1(G227GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U435 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U436 ( .A(KEYINPUT20), .B(n386), .ZN(n387) );
  XNOR2_X1 U437 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U438 ( .A(n390), .B(n389), .ZN(n543) );
  INV_X1 U439 ( .A(n543), .ZN(n471) );
  NOR2_X1 U440 ( .A1(n534), .A2(n471), .ZN(n391) );
  XNOR2_X1 U441 ( .A(KEYINPUT91), .B(n391), .ZN(n410) );
  XOR2_X1 U442 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n393) );
  XNOR2_X1 U443 ( .A(G211GAT), .B(KEYINPUT23), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n409) );
  XOR2_X1 U445 ( .A(KEYINPUT88), .B(G204GAT), .Z(n395) );
  NAND2_X1 U446 ( .A1(G228GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U448 ( .A(n396), .B(KEYINPUT22), .Z(n400) );
  XNOR2_X1 U449 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U450 ( .A(n400), .B(n399), .ZN(n403) );
  XOR2_X1 U451 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n402) );
  XNOR2_X1 U452 ( .A(G141GAT), .B(KEYINPUT87), .ZN(n401) );
  XNOR2_X1 U453 ( .A(n402), .B(n401), .ZN(n419) );
  XOR2_X1 U454 ( .A(n403), .B(n419), .Z(n407) );
  XNOR2_X1 U455 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U456 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U457 ( .A(n409), .B(n408), .Z(n540) );
  NAND2_X1 U458 ( .A1(n410), .A2(n540), .ZN(n411) );
  XOR2_X1 U459 ( .A(KEYINPUT25), .B(n411), .Z(n414) );
  XOR2_X1 U460 ( .A(n534), .B(KEYINPUT27), .Z(n431) );
  NOR2_X1 U461 ( .A1(n540), .A2(n543), .ZN(n412) );
  XNOR2_X1 U462 ( .A(n412), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U463 ( .A1(n431), .A2(n563), .ZN(n413) );
  NAND2_X1 U464 ( .A1(n414), .A2(n413), .ZN(n430) );
  XOR2_X1 U465 ( .A(KEYINPUT1), .B(G57GAT), .Z(n416) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(G148GAT), .ZN(n415) );
  XNOR2_X1 U467 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U468 ( .A(n418), .B(n417), .ZN(n429) );
  XOR2_X1 U469 ( .A(G85GAT), .B(n419), .Z(n421) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(G155GAT), .ZN(n420) );
  XNOR2_X1 U471 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U472 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n423) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U475 ( .A(n425), .B(n424), .Z(n427) );
  XNOR2_X1 U476 ( .A(G162GAT), .B(KEYINPUT6), .ZN(n426) );
  XNOR2_X1 U477 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U478 ( .A(n429), .B(n428), .ZN(n539) );
  INV_X1 U479 ( .A(n539), .ZN(n467) );
  NAND2_X1 U480 ( .A1(n430), .A2(n467), .ZN(n434) );
  XOR2_X1 U481 ( .A(n540), .B(KEYINPUT28), .Z(n488) );
  NAND2_X1 U482 ( .A1(n539), .A2(n431), .ZN(n520) );
  NOR2_X1 U483 ( .A1(n488), .A2(n520), .ZN(n506) );
  XNOR2_X1 U484 ( .A(n506), .B(KEYINPUT90), .ZN(n432) );
  NAND2_X1 U485 ( .A1(n432), .A2(n471), .ZN(n433) );
  NAND2_X1 U486 ( .A1(n434), .A2(n433), .ZN(n449) );
  AND2_X1 U487 ( .A1(n435), .A2(n449), .ZN(n466) );
  NAND2_X1 U488 ( .A1(n452), .A2(n466), .ZN(n436) );
  XNOR2_X1 U489 ( .A(KEYINPUT92), .B(n436), .ZN(n444) );
  NOR2_X1 U490 ( .A1(n444), .A2(n467), .ZN(n438) );
  XNOR2_X1 U491 ( .A(KEYINPUT34), .B(KEYINPUT93), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(n439), .ZN(G1324GAT) );
  NOR2_X1 U494 ( .A1(n534), .A2(n444), .ZN(n440) );
  XOR2_X1 U495 ( .A(KEYINPUT94), .B(n440), .Z(n441) );
  XNOR2_X1 U496 ( .A(G8GAT), .B(n441), .ZN(G1325GAT) );
  NOR2_X1 U497 ( .A1(n444), .A2(n471), .ZN(n443) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(G1326GAT) );
  INV_X1 U500 ( .A(n488), .ZN(n474) );
  NOR2_X1 U501 ( .A1(n444), .A2(n474), .ZN(n445) );
  XOR2_X1 U502 ( .A(G22GAT), .B(n445), .Z(G1327GAT) );
  XOR2_X1 U503 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n447) );
  XNOR2_X1 U504 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT96), .B(KEYINPUT38), .Z(n454) );
  XNOR2_X1 U507 ( .A(KEYINPUT36), .B(KEYINPUT95), .ZN(n448) );
  INV_X1 U508 ( .A(n532), .ZN(n558) );
  XNOR2_X1 U509 ( .A(n448), .B(n558), .ZN(n577) );
  INV_X1 U510 ( .A(n574), .ZN(n529) );
  NAND2_X1 U511 ( .A1(n529), .A2(n449), .ZN(n450) );
  NOR2_X1 U512 ( .A1(n577), .A2(n450), .ZN(n451) );
  XOR2_X1 U513 ( .A(KEYINPUT37), .B(n451), .Z(n480) );
  NAND2_X1 U514 ( .A1(n452), .A2(n480), .ZN(n453) );
  XNOR2_X1 U515 ( .A(n454), .B(n453), .ZN(n463) );
  NAND2_X1 U516 ( .A1(n463), .A2(n539), .ZN(n455) );
  XOR2_X1 U517 ( .A(n456), .B(n455), .Z(G1328GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n458) );
  INV_X1 U519 ( .A(n534), .ZN(n485) );
  NAND2_X1 U520 ( .A1(n463), .A2(n485), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U522 ( .A(G36GAT), .B(n459), .ZN(G1329GAT) );
  XOR2_X1 U523 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n461) );
  NAND2_X1 U524 ( .A1(n463), .A2(n543), .ZN(n460) );
  XNOR2_X1 U525 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U526 ( .A(G43GAT), .B(n462), .ZN(G1330GAT) );
  NAND2_X1 U527 ( .A1(n463), .A2(n488), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n464), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U529 ( .A(n569), .B(KEYINPUT41), .ZN(n523) );
  XNOR2_X1 U530 ( .A(KEYINPUT102), .B(n523), .ZN(n548) );
  INV_X1 U531 ( .A(n565), .ZN(n508) );
  NOR2_X1 U532 ( .A1(n548), .A2(n508), .ZN(n465) );
  XOR2_X1 U533 ( .A(KEYINPUT103), .B(n465), .Z(n481) );
  NAND2_X1 U534 ( .A1(n481), .A2(n466), .ZN(n473) );
  NOR2_X1 U535 ( .A1(n467), .A2(n473), .ZN(n468) );
  XOR2_X1 U536 ( .A(G57GAT), .B(n468), .Z(n469) );
  XNOR2_X1 U537 ( .A(KEYINPUT42), .B(n469), .ZN(G1332GAT) );
  NOR2_X1 U538 ( .A1(n534), .A2(n473), .ZN(n470) );
  XOR2_X1 U539 ( .A(G64GAT), .B(n470), .Z(G1333GAT) );
  NOR2_X1 U540 ( .A1(n471), .A2(n473), .ZN(n472) );
  XOR2_X1 U541 ( .A(G71GAT), .B(n472), .Z(G1334GAT) );
  NOR2_X1 U542 ( .A1(n474), .A2(n473), .ZN(n479) );
  XOR2_X1 U543 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n476) );
  XNOR2_X1 U544 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n475) );
  XNOR2_X1 U545 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U546 ( .A(KEYINPUT104), .B(n477), .ZN(n478) );
  XNOR2_X1 U547 ( .A(n479), .B(n478), .ZN(G1335GAT) );
  XNOR2_X1 U548 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n484) );
  NAND2_X1 U549 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U550 ( .A(n482), .B(KEYINPUT107), .ZN(n489) );
  NAND2_X1 U551 ( .A1(n539), .A2(n489), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n484), .B(n483), .ZN(G1336GAT) );
  NAND2_X1 U553 ( .A1(n485), .A2(n489), .ZN(n486) );
  XNOR2_X1 U554 ( .A(n486), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U555 ( .A1(n489), .A2(n543), .ZN(n487) );
  XNOR2_X1 U556 ( .A(n487), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n491) );
  NAND2_X1 U558 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U559 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(n492), .ZN(G1339GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT112), .B(KEYINPUT47), .Z(n498) );
  XNOR2_X1 U562 ( .A(KEYINPUT110), .B(n574), .ZN(n555) );
  XOR2_X1 U563 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n494) );
  NOR2_X1 U564 ( .A1(n565), .A2(n523), .ZN(n493) );
  XNOR2_X1 U565 ( .A(n494), .B(n493), .ZN(n495) );
  NOR2_X1 U566 ( .A1(n555), .A2(n495), .ZN(n496) );
  NAND2_X1 U567 ( .A1(n496), .A2(n532), .ZN(n497) );
  XNOR2_X1 U568 ( .A(n498), .B(n497), .ZN(n504) );
  XNOR2_X1 U569 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n500) );
  NOR2_X1 U570 ( .A1(n577), .A2(n529), .ZN(n499) );
  XNOR2_X1 U571 ( .A(n500), .B(n499), .ZN(n501) );
  NOR2_X1 U572 ( .A1(n501), .A2(n569), .ZN(n502) );
  NAND2_X1 U573 ( .A1(n565), .A2(n502), .ZN(n503) );
  NAND2_X1 U574 ( .A1(n504), .A2(n503), .ZN(n505) );
  NAND2_X1 U575 ( .A1(n543), .A2(n506), .ZN(n507) );
  NOR2_X1 U576 ( .A1(n536), .A2(n507), .ZN(n517) );
  NAND2_X1 U577 ( .A1(n508), .A2(n517), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n509), .B(KEYINPUT114), .ZN(n510) );
  XNOR2_X1 U579 ( .A(G113GAT), .B(n510), .ZN(G1340GAT) );
  INV_X1 U580 ( .A(n517), .ZN(n511) );
  NOR2_X1 U581 ( .A1(n548), .A2(n511), .ZN(n513) );
  XNOR2_X1 U582 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n512) );
  XNOR2_X1 U583 ( .A(n513), .B(n512), .ZN(G1341GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n515) );
  NAND2_X1 U585 ( .A1(n517), .A2(n555), .ZN(n514) );
  XNOR2_X1 U586 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U587 ( .A(G127GAT), .B(n516), .ZN(G1342GAT) );
  XOR2_X1 U588 ( .A(G134GAT), .B(KEYINPUT51), .Z(n519) );
  NAND2_X1 U589 ( .A1(n517), .A2(n558), .ZN(n518) );
  XNOR2_X1 U590 ( .A(n519), .B(n518), .ZN(G1343GAT) );
  NOR2_X1 U591 ( .A1(n536), .A2(n520), .ZN(n521) );
  NAND2_X1 U592 ( .A1(n521), .A2(n563), .ZN(n531) );
  NOR2_X1 U593 ( .A1(n565), .A2(n531), .ZN(n522) );
  XOR2_X1 U594 ( .A(G141GAT), .B(n522), .Z(G1344GAT) );
  NOR2_X1 U595 ( .A1(n523), .A2(n531), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n525) );
  XNOR2_X1 U597 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n524) );
  XNOR2_X1 U598 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U599 ( .A(KEYINPUT52), .B(n526), .ZN(n527) );
  XNOR2_X1 U600 ( .A(n528), .B(n527), .ZN(G1345GAT) );
  NOR2_X1 U601 ( .A1(n529), .A2(n531), .ZN(n530) );
  XOR2_X1 U602 ( .A(G155GAT), .B(n530), .Z(G1346GAT) );
  NOR2_X1 U603 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U604 ( .A(G162GAT), .B(n533), .Z(G1347GAT) );
  XNOR2_X1 U605 ( .A(n534), .B(KEYINPUT118), .ZN(n535) );
  NOR2_X1 U606 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U607 ( .A(KEYINPUT54), .B(n537), .Z(n538) );
  NAND2_X1 U608 ( .A1(n564), .A2(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n541) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n554), .A2(n565), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G169GAT), .B(n545), .ZN(n546) );
  INV_X1 U613 ( .A(n546), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT120), .B(n547), .ZN(G1348GAT) );
  NOR2_X1 U615 ( .A1(n548), .A2(n554), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n550) );
  XNOR2_X1 U617 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(KEYINPUT56), .B(n551), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1349GAT) );
  XOR2_X1 U621 ( .A(G183GAT), .B(KEYINPUT123), .Z(n557) );
  INV_X1 U622 ( .A(n554), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n559), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(n562), .B(G190GAT), .Z(G1351GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n576) );
  NOR2_X1 U630 ( .A1(n565), .A2(n576), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U635 ( .A(n576), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n573), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(G218GAT), .B(n580), .Z(G1355GAT) );
endmodule

