//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006;
  OAI21_X1  g000(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT14), .ZN(new_n203));
  NOR3_X1   g002(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n202), .A2(KEYINPUT14), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G43gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(G50gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT88), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(KEYINPUT88), .A3(KEYINPUT15), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n209), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n205), .A2(new_n208), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT89), .B1(new_n223), .B2(new_n214), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT17), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n220), .A2(new_n224), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n221), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT16), .A3(new_n232), .ZN(new_n233));
  OAI221_X1 g032(.A(new_n233), .B1(KEYINPUT91), .B2(G8gat), .C1(new_n232), .C2(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235));
  INV_X1    g034(.A(G8gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n226), .A2(new_n230), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT92), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n222), .A2(new_n225), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT93), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n234), .A2(new_n237), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n234), .A2(new_n237), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n238), .A2(KEYINPUT93), .A3(new_n239), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n241), .A2(new_n244), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT94), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT18), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT18), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(KEYINPUT94), .A3(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n250), .B(new_n249), .C1(new_n222), .C2(new_n225), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n243), .B(KEYINPUT13), .Z(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n255), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G113gat), .B(G141gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G169gat), .B(G197gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n257), .A3(new_n261), .A4(new_n268), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G197gat), .A2(G204gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276));
  NAND2_X1  g075(.A1(G211gat), .A2(G218gat), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G211gat), .ZN(new_n280));
  INV_X1    g079(.A(G218gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n277), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n282), .B2(new_n277), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n279), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n286), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n278), .A3(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G155gat), .ZN(new_n292));
  INV_X1    g091(.A(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT78), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G162gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n293), .A2(KEYINPUT78), .ZN(new_n304));
  OAI21_X1  g103(.A(G155gat), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT79), .B1(new_n305), .B2(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n293), .A2(KEYINPUT78), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(G162gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n292), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n301), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(G155gat), .B2(G162gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n299), .B2(KEYINPUT77), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n297), .B2(new_n298), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n296), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n294), .A2(KEYINPUT76), .A3(new_n295), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n313), .A2(new_n314), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n291), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n287), .A2(new_n326), .A3(new_n289), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n314), .A2(new_n328), .B1(new_n313), .B2(new_n324), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT82), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G228gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT78), .B(G162gat), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT79), .B(KEYINPUT2), .C1(new_n335), .C2(new_n292), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n300), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n316), .A2(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT3), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n290), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n328), .A2(new_n314), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n338), .B2(new_n337), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n333), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n330), .B(new_n332), .C1(new_n343), .C2(KEYINPUT82), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n327), .A2(new_n329), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n345), .B(new_n331), .C1(new_n346), .C2(new_n333), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G22gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(G22gat), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT31), .B(G50gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  AOI21_X1  g154(.A(G22gat), .B1(new_n344), .B2(new_n347), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n350), .A2(new_n357), .A3(new_n351), .A4(new_n355), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G15gat), .B(G43gat), .Z(new_n362));
  XNOR2_X1  g161(.A(G71gat), .B(G99gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G113gat), .ZN(new_n370));
  INV_X1    g169(.A(G113gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G120gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n373), .A2(KEYINPUT67), .ZN(new_n374));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT1), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n376), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n374), .A2(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n382), .A2(new_n383), .B1(G169gat), .B2(G176gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385));
  INV_X1    g184(.A(G169gat), .ZN(new_n386));
  INV_X1    g185(.A(G176gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G183gat), .B(G190gat), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n384), .B(new_n390), .C1(new_n383), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(new_n397), .B2(KEYINPUT24), .ZN(new_n398));
  INV_X1    g197(.A(G183gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G190gat), .ZN(new_n400));
  INV_X1    g199(.A(G190gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G183gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n398), .B1(new_n403), .B2(KEYINPUT24), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT25), .A3(new_n390), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n394), .A2(new_n395), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n395), .B1(new_n394), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT26), .B1(new_n386), .B2(new_n387), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n409), .A2(new_n396), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT26), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n397), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(G190gat), .B1(new_n399), .B2(KEYINPUT27), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT65), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT27), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(KEYINPUT65), .A2(KEYINPUT27), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n399), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n415), .B1(new_n420), .B2(KEYINPUT66), .ZN(new_n421));
  AND2_X1   g220(.A1(KEYINPUT65), .A2(KEYINPUT27), .ZN(new_n422));
  NOR2_X1   g221(.A1(KEYINPUT65), .A2(KEYINPUT27), .ZN(new_n423));
  OAI21_X1  g222(.A(G183gat), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT66), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT28), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n417), .A2(G183gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n414), .A2(KEYINPUT28), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n413), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n381), .B1(new_n408), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n392), .A2(new_n393), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT25), .B1(new_n404), .B2(new_n390), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT64), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n394), .A2(new_n395), .A3(new_n405), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n431), .A2(new_n435), .A3(new_n381), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n368), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n366), .B1(new_n439), .B2(KEYINPUT32), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n435), .A3(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(new_n381), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n437), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT33), .B1(new_n444), .B2(new_n368), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT70), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n366), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n367), .B1(new_n443), .B2(new_n437), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT32), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT70), .B1(new_n452), .B2(new_n445), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT71), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT34), .B1(new_n444), .B2(new_n368), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT34), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n443), .A2(new_n457), .A3(new_n367), .A4(new_n437), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n439), .A2(KEYINPUT32), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n366), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n454), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n447), .B1(new_n440), .B2(new_n446), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n452), .A2(KEYINPUT70), .A3(new_n445), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n459), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n361), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G226gat), .ZN(new_n472));
  INV_X1    g271(.A(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n431), .A2(new_n435), .A3(new_n474), .A4(new_n436), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(KEYINPUT29), .ZN(new_n476));
  INV_X1    g275(.A(new_n413), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT28), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n414), .B1(new_n424), .B2(new_n425), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n418), .A2(new_n419), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT66), .B1(new_n480), .B2(G183gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n477), .B1(new_n482), .B2(new_n429), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n433), .A2(new_n434), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n475), .A2(new_n485), .A3(new_n291), .ZN(new_n486));
  XOR2_X1   g285(.A(G8gat), .B(G36gat), .Z(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT73), .ZN(new_n488));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(new_n429), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n491), .A2(new_n413), .B1(new_n394), .B2(new_n405), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n441), .A2(new_n476), .B1(new_n492), .B2(new_n474), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n486), .B(new_n490), .C1(new_n493), .C2(new_n291), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT74), .ZN(new_n495));
  INV_X1    g294(.A(new_n476), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n408), .B2(new_n431), .ZN(new_n497));
  NOR4_X1   g296(.A1(new_n483), .A2(new_n484), .A3(new_n472), .A4(new_n473), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n290), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT74), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n486), .A4(new_n490), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n490), .B1(new_n499), .B2(new_n486), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n495), .A2(new_n501), .B1(new_n502), .B2(KEYINPUT30), .ZN(new_n503));
  INV_X1    g302(.A(new_n490), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n441), .A2(new_n476), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n492), .A2(new_n474), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n291), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n486), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n486), .B1(new_n493), .B2(new_n291), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT75), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n504), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n503), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G1gat), .B(G29gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT0), .ZN(new_n519));
  XNOR2_X1  g318(.A(G57gat), .B(G85gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(new_n520), .Z(new_n521));
  INV_X1    g320(.A(KEYINPUT5), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n442), .B1(new_n337), .B2(new_n338), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n313), .A2(new_n324), .A3(new_n381), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G225gat), .A2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n522), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT3), .B1(new_n337), .B2(new_n338), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n325), .A2(new_n529), .A3(new_n442), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n313), .A2(KEYINPUT4), .A3(new_n324), .A4(new_n381), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n530), .A2(new_n532), .A3(new_n526), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT80), .B1(new_n534), .B2(KEYINPUT5), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n534), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n521), .B(new_n535), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT80), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n522), .A4(new_n526), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n544), .A2(new_n536), .B1(new_n534), .B2(new_n528), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n521), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n548));
  INV_X1    g347(.A(new_n521), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(KEYINPUT6), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n517), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT35), .B1(new_n471), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n547), .A2(new_n551), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n456), .A2(new_n458), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n454), .B2(new_n465), .ZN(new_n558));
  AOI211_X1 g357(.A(new_n556), .B(new_n464), .C1(new_n448), .C2(new_n453), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n512), .A2(new_n513), .A3(new_n504), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n513), .B1(new_n512), .B2(new_n504), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT30), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n495), .A2(new_n501), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n502), .A2(KEYINPUT30), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT84), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT84), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n503), .A2(new_n515), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n555), .A2(new_n361), .A3(new_n560), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n527), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n574), .B(KEYINPUT39), .C1(new_n527), .C2(new_n525), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT39), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n576), .A3(new_n527), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n575), .A2(KEYINPUT40), .A3(new_n521), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT40), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n521), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT39), .B1(new_n525), .B2(new_n527), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n527), .B2(new_n573), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n579), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(new_n546), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n569), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n493), .B2(new_n291), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n475), .A2(new_n485), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n290), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT38), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n494), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n591), .A2(KEYINPUT85), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT85), .B1(new_n591), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT6), .B1(new_n545), .B2(new_n521), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n548), .A2(new_n549), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n510), .A2(new_n514), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n499), .A2(KEYINPUT37), .A3(new_n486), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n596), .A2(new_n599), .A3(new_n550), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n361), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n516), .B1(new_n599), .B2(new_n550), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n469), .A2(new_n556), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n454), .A2(new_n557), .A3(new_n465), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT36), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n460), .B1(new_n454), .B2(new_n465), .ZN(new_n611));
  AOI211_X1 g410(.A(new_n459), .B(new_n464), .C1(new_n448), .C2(new_n453), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI221_X1 g413(.A(new_n606), .B1(new_n607), .B2(new_n361), .C1(new_n610), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n273), .B1(new_n572), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G85gat), .A2(G92gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT7), .ZN(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  INV_X1    g420(.A(G85gat), .ZN(new_n622));
  INV_X1    g421(.A(G92gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(KEYINPUT8), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G99gat), .B(G106gat), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n620), .A3(new_n624), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n629), .A2(new_n632), .B1(new_n627), .B2(new_n625), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n226), .A2(new_n230), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n245), .B2(new_n633), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n618), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT101), .ZN(new_n643));
  XOR2_X1   g442(.A(G134gat), .B(G162gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n635), .A2(new_n639), .A3(new_n618), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n640), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n635), .A2(new_n639), .A3(KEYINPUT103), .A4(new_n618), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI211_X1 g452(.A(KEYINPUT104), .B(new_n645), .C1(new_n649), .C2(new_n650), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(KEYINPUT105), .B(new_n647), .C1(new_n653), .C2(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT21), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n661));
  INV_X1    g460(.A(G57gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(G64gat), .ZN(new_n663));
  INV_X1    g462(.A(G64gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n663), .B(new_n665), .C1(G57gat), .C2(new_n664), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT97), .ZN(new_n667));
  XOR2_X1   g466(.A(G71gat), .B(G78gat), .Z(new_n668));
  AOI21_X1  g467(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(G57gat), .B(G64gat), .Z(new_n672));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n673), .B2(new_n672), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n249), .B(new_n250), .C1(new_n660), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT100), .ZN(new_n679));
  XNOR2_X1  g478(.A(G127gat), .B(G155gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NAND2_X1  g480(.A1(G231gat), .A2(G233gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT98), .Z(new_n683));
  XOR2_X1   g482(.A(new_n681), .B(new_n683), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n679), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n677), .A2(new_n660), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G183gat), .B(G211gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n685), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G230gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n473), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n629), .A2(new_n632), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n627), .B(KEYINPUT106), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n625), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n698), .A2(new_n671), .A3(new_n676), .A4(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT10), .ZN(new_n702));
  INV_X1    g501(.A(new_n677), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n633), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n697), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n701), .B1(new_n703), .B2(new_n633), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n697), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(G120gat), .B(G148gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(G176gat), .B(G204gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n711), .B(new_n712), .Z(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n707), .A2(new_n709), .A3(new_n713), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  AND4_X1   g517(.A1(new_n616), .A2(new_n659), .A3(new_n695), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n554), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G1gat), .ZN(G1324gat));
  INV_X1    g520(.A(new_n570), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n236), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n719), .A2(new_n722), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G8gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n725), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n727), .B1(new_n730), .B2(KEYINPUT42), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1325gat));
  INV_X1    g532(.A(G15gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n734), .A3(new_n560), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n614), .B2(new_n610), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n470), .A2(KEYINPUT36), .A3(new_n466), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n737), .B(new_n738), .C1(new_n560), .C2(KEYINPUT36), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n719), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n735), .B1(new_n742), .B2(new_n734), .ZN(G1326gat));
  NAND2_X1  g542(.A1(new_n359), .A2(new_n360), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n719), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT43), .B(G22gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1327gat));
  NAND2_X1  g546(.A1(new_n572), .A2(new_n615), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n659), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n694), .A2(new_n718), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n273), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n361), .B2(new_n607), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n552), .A2(KEYINPUT110), .A3(new_n744), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n755), .A2(new_n606), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n740), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n659), .B1(new_n758), .B2(new_n572), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n751), .B(new_n753), .C1(new_n759), .C2(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT111), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n757), .A2(new_n740), .B1(new_n553), .B2(new_n571), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n749), .B1(new_n762), .B2(new_n659), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(new_n764), .A3(new_n751), .A4(new_n753), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n554), .ZN(new_n767));
  OAI21_X1  g566(.A(G29gat), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n659), .A2(new_n752), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n616), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n206), .A3(new_n554), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n773), .ZN(G1328gat));
  OAI21_X1  g573(.A(G36gat), .B1(new_n766), .B2(new_n570), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n770), .A2(G36gat), .A3(new_n570), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1329gat));
  INV_X1    g577(.A(new_n560), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n770), .A2(G43gat), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n761), .A2(new_n741), .A3(new_n765), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(G43gat), .ZN(new_n782));
  INV_X1    g581(.A(new_n760), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n210), .B1(new_n783), .B2(new_n741), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n782), .A2(KEYINPUT47), .B1(new_n784), .B2(new_n786), .ZN(G1330gat));
  OAI21_X1  g586(.A(G50gat), .B1(new_n760), .B2(new_n361), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n770), .A2(G50gat), .A3(new_n361), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(KEYINPUT48), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n761), .A2(new_n744), .A3(new_n765), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G50gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n790), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n789), .B1(new_n793), .B2(G50gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n798), .A2(KEYINPUT112), .A3(KEYINPUT48), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n791), .B1(new_n797), .B2(new_n799), .ZN(G1331gat));
  NAND4_X1  g599(.A1(new_n659), .A2(new_n695), .A3(new_n273), .A4(new_n717), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n762), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n554), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g603(.A1(new_n762), .A2(new_n570), .A3(new_n801), .ZN(new_n805));
  NOR2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  AND2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n805), .B2(new_n806), .ZN(G1333gat));
  NAND2_X1  g608(.A1(new_n802), .A2(new_n741), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n779), .A2(G71gat), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n810), .A2(G71gat), .B1(new_n802), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g612(.A1(new_n802), .A2(new_n744), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g614(.A1(new_n273), .A2(new_n694), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n762), .A2(new_n659), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n820), .A2(new_n622), .A3(new_n554), .A4(new_n717), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n763), .A2(new_n751), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n816), .A2(new_n718), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n825), .B2(new_n767), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G85gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n825), .A2(new_n822), .A3(new_n767), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n821), .B1(new_n827), .B2(new_n828), .ZN(G1336gat));
  NAND3_X1  g628(.A1(new_n823), .A2(new_n722), .A3(new_n824), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT114), .B1(new_n830), .B2(G92gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n570), .A2(G92gat), .A3(new_n718), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n820), .A2(new_n833), .B1(G92gat), .B2(new_n830), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n832), .B(new_n834), .ZN(G1337gat));
  NOR3_X1   g634(.A1(new_n779), .A2(G99gat), .A3(new_n718), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G99gat), .B1(new_n825), .B2(new_n740), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1338gat));
  NOR3_X1   g638(.A1(new_n361), .A2(G106gat), .A3(new_n718), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n820), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n744), .A3(new_n824), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G106gat), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT115), .B(new_n840), .C1(new_n818), .C2(new_n819), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT53), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT53), .B1(new_n820), .B2(new_n840), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G106gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(new_n851), .ZN(G1339gat));
  NAND3_X1  g651(.A1(new_n704), .A2(new_n697), .A3(new_n705), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n707), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n713), .B1(new_n706), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(KEYINPUT55), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n716), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT55), .B1(new_n854), .B2(new_n856), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n259), .A2(new_n260), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n244), .B1(new_n241), .B2(new_n252), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n267), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n860), .A2(new_n271), .A3(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n657), .A2(new_n658), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n272), .A2(new_n860), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n271), .A2(new_n717), .A3(new_n863), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n657), .A2(new_n658), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n694), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n659), .A2(new_n695), .A3(new_n273), .A4(new_n718), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n779), .A2(new_n744), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n871), .A2(new_n554), .A3(new_n872), .A4(new_n570), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n371), .A3(new_n273), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n767), .B1(new_n869), .B2(new_n870), .ZN(new_n875));
  INV_X1    g674(.A(new_n471), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n722), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n272), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n874), .B1(new_n879), .B2(new_n371), .ZN(G1340gat));
  NOR3_X1   g679(.A1(new_n873), .A2(new_n369), .A3(new_n718), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n717), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n369), .ZN(G1341gat));
  INV_X1    g682(.A(G127gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n878), .A2(new_n884), .A3(new_n695), .ZN(new_n885));
  OAI21_X1  g684(.A(G127gat), .B1(new_n873), .B2(new_n694), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1342gat));
  NOR2_X1   g686(.A1(new_n659), .A2(new_n722), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT117), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n877), .A2(new_n889), .A3(G134gat), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n892));
  OAI21_X1  g691(.A(G134gat), .B1(new_n873), .B2(new_n659), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G1343gat));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n361), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT119), .B1(new_n858), .B2(new_n859), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n272), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n858), .A2(KEYINPUT119), .A3(new_n859), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n867), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n659), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n865), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n659), .A2(new_n901), .A3(KEYINPUT120), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n695), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n870), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n897), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n361), .B1(new_n869), .B2(new_n870), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT118), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n866), .A2(new_n867), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n659), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n657), .A2(new_n658), .A3(new_n864), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n695), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n744), .B1(new_n914), .B2(new_n907), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n896), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n908), .A2(new_n910), .A3(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n741), .A2(new_n767), .A3(new_n722), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n272), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G141gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n875), .A2(new_n744), .A3(new_n740), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n722), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n273), .A2(G141gat), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT121), .Z(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT58), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n921), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1344gat));
  INV_X1    g730(.A(G148gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n923), .A2(new_n932), .A3(new_n717), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(KEYINPUT59), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n717), .ZN(new_n936));
  XOR2_X1   g735(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n937));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n717), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n695), .B1(new_n902), .B2(new_n913), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n744), .B1(new_n939), .B2(new_n907), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n896), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n871), .A2(new_n897), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n932), .B1(new_n943), .B2(KEYINPUT123), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n937), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n933), .B1(new_n936), .B2(new_n946), .ZN(G1345gat));
  NAND3_X1  g746(.A1(new_n918), .A2(new_n695), .A3(new_n919), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G155gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n923), .A2(new_n292), .A3(new_n695), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1346gat));
  INV_X1    g754(.A(new_n659), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n335), .B1(new_n935), .B2(new_n956), .ZN(new_n957));
  NOR4_X1   g756(.A1(new_n922), .A2(new_n889), .A3(new_n303), .A4(new_n304), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n570), .A2(new_n554), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n961), .B1(new_n869), .B2(new_n870), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n872), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n963), .A2(new_n386), .A3(new_n273), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n876), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n272), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n964), .B1(new_n967), .B2(new_n386), .ZN(G1348gat));
  NAND3_X1  g767(.A1(new_n966), .A2(new_n387), .A3(new_n717), .ZN(new_n969));
  OAI21_X1  g768(.A(G176gat), .B1(new_n963), .B2(new_n718), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1349gat));
  OAI21_X1  g770(.A(G183gat), .B1(new_n963), .B2(new_n694), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n399), .A2(KEYINPUT27), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n695), .A2(new_n973), .A3(new_n428), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n966), .A2(new_n401), .A3(new_n956), .ZN(new_n977));
  OAI21_X1  g776(.A(G190gat), .B1(new_n963), .B2(new_n659), .ZN(new_n978));
  XNOR2_X1  g777(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n978), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(G1351gat));
  NOR2_X1   g782(.A1(new_n741), .A2(new_n961), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n909), .A2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(G197gat), .B1(new_n986), .B2(new_n272), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n941), .A2(new_n942), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n984), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n272), .A2(G197gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(G1352gat));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g792(.A(G204gat), .B1(new_n993), .B2(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n986), .A2(new_n717), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n995), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g796(.A(G204gat), .B1(new_n989), .B2(new_n718), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(G1353gat));
  NAND3_X1  g798(.A1(new_n986), .A2(new_n280), .A3(new_n695), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n990), .A2(new_n695), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n1001), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(KEYINPUT63), .B1(new_n1001), .B2(G211gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(G1354gat));
  OAI21_X1  g803(.A(G218gat), .B1(new_n989), .B2(new_n659), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n281), .A3(new_n956), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1355gat));
endmodule


