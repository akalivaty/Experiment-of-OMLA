//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n545, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT65), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n465), .A2(new_n467), .A3(G137), .A4(new_n463), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n465), .A2(new_n467), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(new_n475), .B2(new_n463), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n478), .A2(new_n484), .A3(new_n486), .ZN(G162));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n465), .A2(new_n467), .A3(G126), .A4(G2105), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT70), .A2(G138), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n467), .A3(new_n492), .A4(new_n463), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n481), .A2(KEYINPUT4), .A3(new_n463), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n500), .B(new_n502), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n504), .A2(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT71), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(new_n506), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n499), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n511), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(new_n509), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n500), .A2(new_n502), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(G168));
  AND2_X1   g103(.A1(G77), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n515), .B2(G64), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n499), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(G90), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G52), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n522), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(new_n522), .A2(G43), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n503), .A2(G81), .A3(new_n515), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n499), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT74), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n543), .A2(new_n547), .ZN(G188));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n509), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(KEYINPUT75), .B1(new_n503), .B2(new_n515), .ZN(new_n551));
  OAI21_X1  g126(.A(G91), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n522), .A2(G53), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n522), .A2(new_n555), .A3(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  OAI21_X1  g134(.A(G65), .B1(new_n507), .B2(new_n508), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n559), .B1(new_n562), .B2(G651), .ZN(new_n563));
  AOI211_X1 g138(.A(KEYINPUT76), .B(new_n499), .C1(new_n560), .C2(new_n561), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n558), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n509), .A2(new_n549), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n503), .A2(KEYINPUT75), .A3(new_n515), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G91), .B1(new_n554), .B2(new_n556), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT76), .B1(new_n572), .B2(new_n499), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n562), .A2(new_n559), .A3(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT77), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND2_X1  g155(.A1(new_n570), .A2(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n522), .A2(G49), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  AOI22_X1  g159(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n499), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n522), .A2(G48), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n570), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n520), .A2(G85), .B1(G47), .B2(new_n522), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n499), .B2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(G92), .B1(new_n550), .B2(new_n551), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n515), .A2(G66), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n499), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(G54), .B2(new_n522), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n570), .A2(new_n602), .A3(G92), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n597), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n577), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n577), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g192(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2100), .Z(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n624), .B(new_n625), .C1(G111), .C2(new_n463), .ZN(new_n626));
  INV_X1    g201(.A(new_n476), .ZN(new_n627));
  INV_X1    g202(.A(G135), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G123), .B2(new_n483), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n621), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(KEYINPUT14), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n639), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n636), .A2(new_n637), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n640), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n640), .B2(new_n645), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  NOR3_X1   g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n648), .B1(new_n646), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT82), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n654), .B(new_n648), .C1(new_n646), .C2(new_n647), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT83), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  OAI21_X1  g240(.A(KEYINPUT17), .B1(new_n659), .B2(new_n663), .ZN(new_n666));
  AOI22_X1  g241(.A1(new_n666), .A2(new_n660), .B1(new_n659), .B2(new_n663), .ZN(new_n667));
  OAI211_X1 g242(.A(KEYINPUT17), .B(new_n661), .C1(new_n659), .C2(new_n663), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT84), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n676), .A2(new_n677), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n678), .A3(new_n680), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n683), .B(new_n685), .C1(new_n680), .C2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G33), .ZN(new_n695));
  NAND2_X1  g270(.A1(G115), .A2(G2104), .ZN(new_n696));
  INV_X1    g271(.A(G127), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n475), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G2105), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT25), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n476), .A2(G139), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT92), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n698), .A2(G2105), .B1(new_n476), .B2(G139), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n701), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n695), .B1(new_n709), .B2(new_n694), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G2072), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(new_n694), .ZN(new_n714));
  INV_X1    g289(.A(G160), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n694), .ZN(new_n716));
  INV_X1    g291(.A(G2084), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n483), .A2(G129), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT26), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n481), .A2(G141), .A3(new_n463), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n724));
  AND3_X1   g299(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G29), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n718), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n711), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT94), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G4), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n606), .B2(new_n734), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1348), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n711), .A2(new_n738), .A3(new_n731), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n716), .A2(new_n717), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g316(.A1(G164), .A2(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G27), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT30), .B(G28), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n743), .A2(new_n744), .B1(new_n694), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n741), .B(new_n746), .C1(new_n744), .C2(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(G168), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G16), .B2(G21), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  NOR2_X1   g325(.A1(G5), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G171), .B2(G16), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n749), .A2(new_n750), .B1(new_n752), .B2(G1961), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n733), .A2(new_n737), .A3(new_n739), .A4(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n734), .A2(KEYINPUT23), .A3(G20), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT23), .ZN(new_n757));
  INV_X1    g332(.A(G20), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G16), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n759), .C1(new_n577), .C2(new_n734), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT96), .B(G1956), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n729), .A2(new_n730), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n736), .A2(G1348), .B1(G1961), .B2(new_n752), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n630), .A2(G29), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n541), .A2(new_n734), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n734), .B2(G19), .ZN(new_n767));
  INV_X1    g342(.A(G1341), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n768), .B2(new_n767), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n764), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n755), .A2(new_n762), .A3(new_n763), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G35), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G162), .B2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT29), .B(G2090), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n694), .A2(G25), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n475), .A2(new_n479), .A3(new_n463), .ZN(new_n779));
  AOI21_X1  g354(.A(KEYINPUT69), .B1(new_n481), .B2(G2105), .ZN(new_n780));
  OAI21_X1  g355(.A(G119), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n463), .A2(G107), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n782), .A2(new_n783), .A3(KEYINPUT87), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT87), .B1(new_n782), .B2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n476), .A2(G131), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n781), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n778), .B1(new_n788), .B2(new_n694), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT35), .B(G1991), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT88), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G24), .B(G290), .S(G16), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1986), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n792), .B(new_n794), .C1(KEYINPUT90), .C2(KEYINPUT36), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n734), .A2(G23), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G288), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT33), .ZN(new_n798));
  INV_X1    g373(.A(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT89), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G166), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G16), .B2(G22), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1971), .Z(new_n807));
  NOR2_X1   g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n800), .A2(KEYINPUT34), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(KEYINPUT34), .B1(new_n800), .B2(new_n808), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n795), .B1(KEYINPUT90), .B2(KEYINPUT36), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n795), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g387(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n773), .A2(new_n777), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n694), .A2(G26), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n483), .A2(G128), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n476), .A2(G140), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n819));
  NOR2_X1   g394(.A1(G104), .A2(G2105), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT91), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n816), .B1(new_n823), .B2(new_n694), .ZN(new_n824));
  MUX2_X1   g399(.A(new_n816), .B(new_n824), .S(KEYINPUT28), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2067), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n749), .A2(new_n750), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n815), .A2(new_n826), .A3(new_n828), .ZN(G311));
  AND3_X1   g404(.A1(new_n773), .A2(new_n811), .A3(new_n814), .ZN(new_n830));
  INV_X1    g405(.A(new_n826), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n830), .A2(new_n831), .A3(new_n827), .A4(new_n777), .ZN(G150));
  NAND2_X1  g407(.A1(new_n522), .A2(G55), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT97), .B(G93), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n503), .A2(new_n515), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n835), .C1(new_n836), .C2(new_n499), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n604), .B(KEYINPUT78), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n612), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n541), .A2(new_n837), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n833), .A2(new_n835), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n515), .A2(G67), .ZN(new_n845));
  NAND2_X1  g420(.A1(G80), .A2(G543), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n499), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n540), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT39), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n842), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n839), .B1(new_n852), .B2(G860), .ZN(G145));
  NAND2_X1  g428(.A1(new_n483), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n476), .A2(G142), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n781), .A2(new_n786), .A3(new_n787), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n788), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT100), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n859), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n788), .A2(new_n861), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n863), .A2(new_n619), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n619), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n864), .B2(new_n865), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n495), .A2(new_n496), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n489), .A2(new_n490), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n491), .A2(KEYINPUT98), .A3(new_n495), .A4(new_n496), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n726), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n726), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n823), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n708), .A2(KEYINPUT99), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n704), .A2(new_n883), .A3(new_n707), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n876), .A2(new_n877), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n727), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n823), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n878), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n881), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n881), .A2(new_n889), .B1(new_n883), .B2(new_n709), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n868), .B(new_n872), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n889), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n888), .B1(new_n887), .B2(new_n878), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n884), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n881), .A2(new_n885), .A3(new_n889), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n870), .A2(new_n871), .A3(new_n869), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n619), .B1(new_n863), .B2(new_n867), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n630), .B(new_n715), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G162), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n892), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n892), .B2(new_n899), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G37), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  NOR4_X1   g482(.A1(new_n840), .A2(G559), .A3(new_n849), .A4(new_n843), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n850), .B1(new_n606), .B2(new_n612), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n604), .B1(new_n567), .B2(new_n576), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n566), .B1(new_n558), .B2(new_n565), .ZN(new_n912));
  INV_X1    g487(.A(G92), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(new_n568), .B2(new_n569), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT10), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n571), .A2(new_n575), .A3(KEYINPUT77), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n912), .A2(new_n915), .A3(new_n916), .A4(new_n601), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n567), .A2(new_n576), .A3(new_n604), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n912), .A2(new_n916), .B1(new_n915), .B2(new_n601), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT41), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n911), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(KEYINPUT101), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n911), .A2(new_n917), .A3(new_n926), .A4(new_n923), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n919), .B1(new_n928), .B2(new_n910), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n930));
  XNOR2_X1  g505(.A(G288), .B(G290), .ZN(new_n931));
  XNOR2_X1  g506(.A(G305), .B(G166), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n919), .B(new_n934), .C1(new_n928), .C2(new_n910), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n930), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n930), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g514(.A(new_n938), .B1(G868), .B2(new_n848), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n941));
  AOI21_X1  g516(.A(G168), .B1(KEYINPUT102), .B2(G301), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n541), .A2(new_n837), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n848), .A2(new_n540), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n531), .A2(new_n946), .A3(new_n532), .A4(new_n534), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n946), .B(G171), .C1(new_n843), .C2(new_n849), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n942), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n925), .A2(new_n927), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n933), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n918), .B1(new_n953), .B2(new_n950), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n954), .B1(new_n922), .B2(new_n924), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n933), .B1(new_n961), .B2(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n905), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n941), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(KEYINPUT103), .A3(new_n905), .A4(new_n962), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT104), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n956), .A2(new_n959), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n933), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n971), .A2(new_n905), .A3(new_n965), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n964), .A2(new_n975), .A3(KEYINPUT43), .A4(new_n966), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n905), .A4(new_n965), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n973), .B1(new_n960), .B2(new_n963), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n969), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(G397));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT45), .B1(new_n886), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n468), .A2(new_n469), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(G2105), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n471), .A2(new_n472), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(G40), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(G160), .A2(KEYINPUT105), .A3(G40), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n983), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(G1996), .A3(new_n726), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT106), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n823), .B(G2067), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G1996), .B2(new_n726), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n992), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n859), .A2(new_n791), .ZN(new_n999));
  OAI22_X1  g574(.A1(new_n998), .A2(new_n999), .B1(G2067), .B2(new_n888), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n992), .ZN(new_n1001));
  INV_X1    g576(.A(new_n992), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1002), .A2(G1986), .A3(G290), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT48), .Z(new_n1004));
  INV_X1    g579(.A(new_n998), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n859), .B(new_n791), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n992), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n992), .A2(KEYINPUT46), .A3(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT126), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1002), .B1(new_n727), .B2(new_n995), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n992), .B2(new_n1010), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT125), .Z(new_n1016));
  AOI21_X1  g591(.A(new_n1009), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1014), .A2(new_n1009), .A3(new_n1016), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1001), .B(new_n1008), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT108), .B(G8), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n982), .B1(new_n874), .B2(new_n875), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n991), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n503), .A2(G86), .A3(new_n515), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n587), .B(new_n1026), .C1(new_n585), .C2(new_n499), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G1981), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT110), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n589), .A2(new_n590), .A3(new_n690), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1031), .A3(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1029), .A2(new_n1030), .A3(KEYINPUT49), .A4(new_n1032), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1025), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G288), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n799), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1030), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(G1976), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1025), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT109), .B(G1976), .Z(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1025), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1037), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(G166), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT55), .B(G8), .C1(new_n511), .C2(new_n518), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n886), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT45), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n989), .A2(new_n990), .B1(new_n1023), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1971), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n497), .A2(new_n1062), .A3(new_n982), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n991), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(G2090), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1056), .B(G8), .C1(new_n1060), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1025), .A2(new_n1040), .B1(new_n1048), .B2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT112), .B(KEYINPUT63), .Z(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1047), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1021), .B1(new_n1065), .B2(new_n1060), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1064), .A2(G2084), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1024), .A2(KEYINPUT45), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1966), .B1(new_n1059), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(G286), .B(new_n1022), .C1(new_n1075), .C2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .A4(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1048), .A2(new_n1079), .A3(new_n1074), .A4(new_n1066), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT111), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1069), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1065), .A2(new_n1060), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT113), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT113), .B(G8), .C1(new_n1065), .C2(new_n1060), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1073), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AND4_X1   g663(.A1(KEYINPUT63), .A2(new_n1088), .A3(new_n1070), .A4(new_n1079), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1068), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT118), .B1(new_n1091), .B2(G8), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1064), .A2(G2084), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT118), .B(G8), .C1(new_n1093), .C2(new_n1077), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G168), .A2(new_n1022), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(new_n1021), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n1096), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1098), .A2(new_n1101), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1059), .A2(new_n744), .A3(new_n1076), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1059), .A2(KEYINPUT119), .A3(new_n744), .A4(new_n1076), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT53), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1057), .A2(new_n1059), .A3(new_n744), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT120), .B(G1961), .Z(new_n1111));
  AOI22_X1  g686(.A1(new_n1109), .A2(new_n1110), .B1(new_n1064), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT122), .B1(new_n1113), .B2(G171), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n1115));
  AOI211_X1 g690(.A(new_n1115), .B(G301), .C1(new_n1108), .C2(new_n1112), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1102), .B1(new_n1103), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1057), .A2(new_n1059), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n558), .B2(new_n565), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n571), .A2(new_n575), .A3(KEYINPUT57), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1064), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1057), .A2(new_n1059), .A3(KEYINPUT114), .A4(new_n1119), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1122), .A2(new_n1126), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1348), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT105), .B1(G160), .B2(G40), .ZN(new_n1133));
  INV_X1    g708(.A(G40), .ZN(new_n1134));
  NOR4_X1   g709(.A1(new_n470), .A2(new_n473), .A3(new_n988), .A4(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1131), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G2067), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n991), .A2(new_n1138), .A3(new_n1024), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n604), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1130), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1122), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1124), .A2(KEYINPUT115), .A3(new_n1125), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT115), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT116), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1141), .A2(new_n1149), .A3(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1146), .A2(new_n1130), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n1139), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1153), .A2(KEYINPUT117), .A3(new_n604), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n604), .B1(new_n1153), .B2(KEYINPUT117), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1154), .A2(new_n1155), .B1(KEYINPUT117), .B2(new_n1153), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1157), .A2(KEYINPUT60), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1152), .A2(KEYINPUT61), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1142), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT61), .B1(new_n1160), .B2(new_n1130), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1057), .A2(new_n1059), .A3(new_n1010), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT58), .B(G1341), .Z(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1136), .B2(new_n1023), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n540), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT59), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1151), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1113), .A2(G301), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT53), .B1(KEYINPUT123), .B2(G2078), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n983), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n987), .B1(KEYINPUT123), .B2(G2078), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1057), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1112), .A2(new_n1173), .A3(G171), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1169), .A2(KEYINPUT54), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1112), .A2(new_n1173), .A3(G301), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(KEYINPUT124), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1114), .A2(new_n1116), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT54), .B1(new_n1176), .B2(KEYINPUT124), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1118), .B1(new_n1168), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(new_n1102), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1090), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(G290), .B(G1986), .Z(new_n1186));
  OAI211_X1 g761(.A(new_n1005), .B(new_n1007), .C1(new_n1002), .C2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1020), .B1(new_n1185), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g763(.A1(new_n656), .A2(new_n673), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1190), .B1(new_n904), .B2(new_n905), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G229), .A2(new_n461), .ZN(new_n1192));
  NAND4_X1  g766(.A1(new_n1191), .A2(new_n978), .A3(new_n979), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  XNOR2_X1  g768(.A(new_n1193), .B(new_n1194), .ZN(G308));
  XNOR2_X1  g769(.A(new_n1193), .B(KEYINPUT127), .ZN(G225));
endmodule


