//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n203));
  MUX2_X1   g002(.A(G183gat), .B(new_n203), .S(G190gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n207), .B2(KEYINPUT24), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(KEYINPUT64), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n204), .A2(new_n208), .A3(new_n213), .A4(new_n210), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT23), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220));
  OR2_X1    g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n212), .A2(new_n214), .A3(new_n217), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT24), .B1(new_n206), .B2(KEYINPUT68), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(KEYINPUT68), .B2(new_n206), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n204), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n229), .B(new_n218), .C1(new_n221), .C2(new_n220), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n218), .B1(new_n221), .B2(new_n220), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n224), .B1(new_n221), .B2(new_n220), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n228), .A2(new_n230), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT71), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT71), .A3(G134gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G113gat), .ZN(new_n243));
  INV_X1    g042(.A(G113gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G120gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT1), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT72), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT72), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n248), .A2(new_n238), .A3(new_n249), .A4(new_n240), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n236), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT27), .B(G183gat), .Z(new_n254));
  OAI21_X1  g053(.A(KEYINPUT28), .B1(new_n254), .B2(G190gat), .ZN(new_n255));
  INV_X1    g054(.A(G183gat), .ZN(new_n256));
  OR3_X1    g055(.A1(new_n256), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT27), .B1(new_n256), .B2(KEYINPUT69), .ZN(new_n258));
  NOR2_X1   g057(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n255), .A2(new_n263), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n221), .A2(KEYINPUT26), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n219), .B1(KEYINPUT26), .B2(new_n221), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n207), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n235), .A2(new_n253), .A3(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n247), .A2(new_n250), .B1(new_n246), .B2(new_n236), .ZN(new_n272));
  INV_X1    g071(.A(new_n234), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n223), .B2(new_n224), .ZN(new_n274));
  INV_X1    g073(.A(new_n269), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n262), .B2(new_n264), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G227gat), .ZN(new_n279));
  INV_X1    g078(.A(G233gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n279), .A2(new_n280), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n271), .A2(new_n277), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G15gat), .B(G43gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT33), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT73), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n271), .A2(new_n277), .A3(new_n284), .A4(new_n289), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT73), .B1(new_n293), .B2(new_n290), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n283), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n283), .A2(new_n296), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n300));
  INV_X1    g099(.A(G50gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G228gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(new_n280), .ZN(new_n307));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n313), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT3), .B1(new_n318), .B2(KEYINPUT82), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n313), .B(new_n314), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(KEYINPUT29), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n325), .B1(new_n328), .B2(KEYINPUT2), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT77), .B1(new_n330), .B2(G141gat), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(G148gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n330), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n325), .B(new_n328), .C1(new_n336), .C2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n324), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n316), .B1(new_n342), .B2(new_n317), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n307), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n346), .A2(new_n307), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n340), .B2(new_n318), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(new_n343), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n345), .A2(G22gat), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G22gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n349), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n340), .B1(new_n319), .B2(new_n323), .ZN(new_n353));
  OAI22_X1  g152(.A1(new_n353), .A2(new_n343), .B1(new_n306), .B2(new_n280), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n305), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(G22gat), .B1(new_n345), .B2(new_n349), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT84), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n354), .A3(new_n351), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n360), .A2(new_n362), .A3(new_n304), .A4(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT83), .B(new_n305), .C1(new_n350), .C2(new_n355), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n299), .A2(KEYINPUT88), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n342), .A2(new_n346), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT78), .B1(new_n370), .B2(new_n272), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n253), .A2(new_n372), .A3(new_n346), .A4(new_n342), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n272), .A2(new_n375), .A3(new_n340), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n272), .A2(KEYINPUT79), .A3(new_n375), .A4(new_n340), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n272), .A2(new_n340), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n253), .A2(new_n338), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n380), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n386), .B2(new_n369), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  AOI21_X1  g191(.A(KEYINPUT5), .B1(new_n381), .B2(new_n376), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT80), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n388), .A2(new_n394), .ZN(new_n397));
  INV_X1    g196(.A(new_n392), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n383), .A2(new_n387), .B1(new_n374), .B2(new_n393), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n392), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n396), .A2(new_n399), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n217), .A2(new_n222), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(KEYINPUT65), .B2(new_n211), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT25), .B1(new_n408), .B2(new_n214), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n270), .B1(new_n409), .B2(new_n273), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n410), .A2(new_n317), .B1(G226gat), .B2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(G226gat), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n412), .B(new_n280), .C1(new_n235), .C2(new_n270), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n320), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n274), .A2(new_n276), .ZN(new_n415));
  OAI22_X1  g214(.A1(new_n415), .A2(KEYINPUT29), .B1(new_n412), .B2(new_n280), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(G226gat), .A3(G233gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n316), .ZN(new_n418));
  XOR2_X1   g217(.A(G8gat), .B(G36gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT75), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n414), .A2(new_n418), .A3(KEYINPUT30), .A4(new_n423), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n424), .A2(KEYINPUT76), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n411), .A2(new_n413), .A3(new_n320), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n316), .B1(new_n416), .B2(new_n417), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT76), .A3(new_n424), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n423), .A3(new_n418), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n425), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n406), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n299), .A2(new_n366), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n202), .B(new_n367), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n358), .A2(new_n364), .A3(new_n365), .ZN(new_n437));
  INV_X1    g236(.A(new_n282), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n281), .B(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(new_n292), .C1(new_n295), .C2(new_n294), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n283), .A2(new_n296), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n430), .A2(new_n431), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n444), .A2(KEYINPUT76), .A3(new_n424), .A4(new_n428), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n404), .A2(new_n405), .B1(new_n445), .B2(new_n425), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n443), .B(new_n446), .C1(KEYINPUT88), .C2(KEYINPUT35), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n371), .A2(new_n373), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n381), .A2(new_n376), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n368), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT85), .B(KEYINPUT39), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n392), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n385), .A2(new_n368), .A3(new_n380), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT39), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n455), .B2(KEYINPUT39), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n451), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n448), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  OR3_X1    g259(.A1(new_n451), .A2(new_n457), .A3(new_n458), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n398), .B1(new_n451), .B2(new_n452), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(KEYINPUT40), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n463), .A3(new_n399), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n366), .B1(new_n433), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n414), .A2(new_n466), .A3(new_n418), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n426), .B2(new_n427), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n422), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n470), .B2(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n414), .A2(new_n418), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n423), .B1(new_n472), .B2(KEYINPUT37), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT38), .ZN(new_n477));
  INV_X1    g276(.A(new_n430), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n467), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n480), .B2(new_n473), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n481), .A2(new_n404), .A3(new_n405), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n465), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n297), .B2(new_n298), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n440), .A2(KEYINPUT36), .A3(new_n441), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n446), .B2(new_n366), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n436), .B(new_n447), .C1(new_n483), .C2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT16), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(G1gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G1gat), .B2(new_n490), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(G8gat), .Z(new_n494));
  INV_X1    g293(.A(G43gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(new_n301), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT91), .B(G50gat), .ZN(new_n497));
  AOI211_X1 g296(.A(KEYINPUT15), .B(new_n496), .C1(new_n497), .C2(new_n495), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(G29gat), .A2(G36gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT14), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT90), .B(G29gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(G36gat), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT15), .B1(new_n496), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n498), .B2(new_n499), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n504), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n510), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(KEYINPUT17), .ZN(new_n516));
  AOI211_X1 g315(.A(KEYINPUT93), .B(new_n512), .C1(new_n508), .C2(new_n510), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n494), .B(new_n513), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n494), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT18), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n515), .A2(new_n494), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n519), .B(KEYINPUT13), .Z(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT94), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n518), .A2(KEYINPUT18), .A3(new_n519), .A4(new_n521), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT12), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n524), .A2(new_n532), .A3(new_n533), .A4(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n489), .A2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G57gat), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n557), .A2(G64gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(G64gat), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n554), .B(new_n556), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n549), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n553), .A2(new_n549), .A3(new_n560), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT21), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT97), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G183gat), .B(G211gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n569), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n553), .A2(new_n549), .A3(new_n560), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n576), .A2(new_n561), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(new_n520), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT100), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n575), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT102), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G99gat), .ZN(new_n588));
  INV_X1    g387(.A(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT102), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT7), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT7), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(G85gat), .A3(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G85gat), .ZN(new_n600));
  INV_X1    g399(.A(G92gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n587), .A2(new_n593), .A3(new_n599), .A4(new_n602), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n513), .B(new_n606), .C1(new_n516), .C2(new_n517), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  AND2_X1   g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n511), .A2(new_n608), .B1(KEYINPUT41), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n584), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n607), .A2(new_n584), .A3(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G134gat), .B(G162gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT101), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT110), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n606), .B1(new_n576), .B2(new_n561), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT104), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n606), .B(new_n628), .C1(new_n576), .C2(new_n561), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n608), .A2(new_n562), .A3(new_n563), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n606), .A2(new_n576), .A3(new_n561), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT105), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n630), .A2(new_n646), .A3(new_n633), .A4(new_n635), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT106), .B1(new_n631), .B2(new_n646), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n649), .A3(KEYINPUT10), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT107), .B1(new_n652), .B2(new_n637), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654));
  AOI211_X1 g453(.A(new_n654), .B(new_n638), .C1(new_n647), .C2(new_n651), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n645), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT108), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n645), .B(new_n658), .C1(new_n653), .C2(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n637), .B(KEYINPUT109), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n643), .B1(new_n662), .B2(new_n639), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n625), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  AOI211_X1 g464(.A(KEYINPUT110), .B(new_n663), .C1(new_n657), .C2(new_n659), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n582), .A2(new_n624), .A3(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n546), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n406), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  INV_X1    g472(.A(new_n433), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n675), .A2(G8gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT42), .B2(new_n678), .ZN(G1325gat));
  INV_X1    g479(.A(G15gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n670), .A2(new_n681), .A3(new_n299), .ZN(new_n682));
  INV_X1    g481(.A(new_n487), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n670), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n684), .B2(new_n681), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n437), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT111), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  AND4_X1   g488(.A1(new_n546), .A2(new_n624), .A3(new_n582), .A4(new_n667), .ZN(new_n690));
  INV_X1    g489(.A(new_n503), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n671), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n436), .A2(new_n447), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT112), .B1(new_n483), .B2(new_n488), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n460), .A2(new_n399), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n697), .A2(new_n445), .A3(new_n425), .A4(new_n463), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n479), .B1(new_n471), .B2(new_n475), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n481), .A2(new_n404), .A3(new_n405), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n698), .B(new_n366), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n434), .A2(new_n437), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .A4(new_n487), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n695), .B1(new_n696), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n694), .B1(new_n705), .B2(new_n623), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n489), .A2(KEYINPUT44), .A3(new_n624), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n581), .A2(new_n668), .A3(new_n544), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n503), .B1(new_n710), .B2(new_n406), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n711), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n690), .A2(new_n713), .A3(new_n674), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT46), .Z(new_n715));
  OAI21_X1  g514(.A(G36gat), .B1(new_n710), .B2(new_n433), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  NAND2_X1  g516(.A1(new_n683), .A2(G43gat), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n690), .A2(new_n299), .ZN(new_n719));
  OAI22_X1  g518(.A1(new_n710), .A2(new_n718), .B1(new_n719), .B2(G43gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g520(.A(new_n497), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n710), .B2(new_n366), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n690), .A2(new_n437), .A3(new_n497), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT48), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n723), .B(new_n724), .C1(new_n726), .C2(KEYINPUT48), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  NAND3_X1  g529(.A1(new_n581), .A2(new_n544), .A3(new_n623), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n705), .A2(new_n667), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n671), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n674), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT49), .B(G64gat), .Z(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n732), .A2(new_n739), .A3(new_n299), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n732), .A2(new_n683), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n739), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n437), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n705), .A2(new_n623), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n581), .A2(new_n545), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT51), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  INV_X1    g548(.A(new_n747), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n705), .A2(new_n749), .A3(new_n623), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OR4_X1    g551(.A1(G85gat), .A2(new_n752), .A3(new_n406), .A4(new_n667), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n750), .A2(new_n667), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n706), .A2(new_n707), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n706), .A2(KEYINPUT114), .A3(new_n707), .A4(new_n754), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n757), .A2(new_n671), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(new_n600), .B2(new_n759), .ZN(G1336gat));
  NOR2_X1   g559(.A1(new_n433), .A2(G92gat), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n668), .B(new_n761), .C1(new_n748), .C2(new_n751), .ZN(new_n762));
  OAI21_X1  g561(.A(G92gat), .B1(new_n755), .B2(new_n433), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n757), .A2(new_n674), .A3(new_n758), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n762), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n764), .ZN(G1337gat));
  AND4_X1   g568(.A1(G99gat), .A2(new_n757), .A3(new_n683), .A4(new_n758), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n299), .B(new_n668), .C1(new_n748), .C2(new_n751), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n588), .B2(new_n771), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n437), .A3(new_n758), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(G106gat), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n667), .A2(G106gat), .A3(new_n366), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT115), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n748), .B2(new_n751), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT116), .B(new_n776), .C1(new_n748), .C2(new_n751), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n774), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G106gat), .B1(new_n755), .B2(new_n366), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  INV_X1    g583(.A(new_n775), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n783), .B(new_n784), .C1(new_n752), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(G1339gat));
  NOR3_X1   g586(.A1(new_n674), .A2(new_n406), .A3(new_n442), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n669), .A2(new_n544), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT54), .B1(new_n652), .B2(new_n661), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n652), .A2(new_n637), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n654), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n652), .A2(KEYINPUT107), .A3(new_n637), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n644), .B1(new_n662), .B2(KEYINPUT54), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n796), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n653), .A2(new_n655), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n798), .B(KEYINPUT55), .C1(new_n799), .C2(new_n791), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n660), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n544), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n519), .B1(new_n518), .B2(new_n521), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n526), .A2(new_n527), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n539), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n543), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n665), .B2(new_n666), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n624), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n811));
  NOR4_X1   g610(.A1(new_n810), .A2(new_n801), .A3(new_n811), .A4(new_n623), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n582), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n789), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT118), .B1(new_n814), .B2(new_n366), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n816), .B(new_n437), .C1(new_n789), .C2(new_n813), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n788), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT119), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n788), .C1(new_n815), .C2(new_n817), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n819), .A2(G113gat), .A3(new_n545), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n406), .B1(new_n789), .B2(new_n813), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n435), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n433), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n244), .B1(new_n826), .B2(new_n544), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n822), .A2(new_n827), .ZN(G1340gat));
  NAND4_X1  g627(.A1(new_n819), .A2(G120gat), .A3(new_n668), .A4(new_n821), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n242), .B1(new_n826), .B2(new_n667), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(G1341gat));
  AND3_X1   g630(.A1(new_n819), .A2(new_n581), .A3(new_n821), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n581), .A2(new_n239), .ZN(new_n833));
  OAI22_X1  g632(.A1(new_n832), .A2(new_n239), .B1(new_n826), .B2(new_n833), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n674), .A2(new_n623), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n825), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT56), .Z(new_n838));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n624), .A3(new_n821), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G134gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1343gat));
  XOR2_X1   g640(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n842));
  NOR2_X1   g641(.A1(new_n674), .A2(new_n406), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n487), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n366), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n793), .A2(new_n794), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n658), .B1(new_n847), .B2(new_n645), .ZN(new_n848));
  INV_X1    g647(.A(new_n659), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n664), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT110), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n660), .A2(new_n625), .A3(new_n664), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n806), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n544), .A2(new_n801), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT120), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n802), .A2(new_n808), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n623), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n812), .B1(new_n858), .B2(KEYINPUT121), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n855), .A2(new_n860), .A3(new_n623), .A4(new_n857), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n581), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n789), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n846), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n814), .A2(new_n437), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n845), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n844), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n332), .B1(new_n867), .B2(new_n545), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n824), .A2(KEYINPUT122), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n683), .A2(new_n366), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n823), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n544), .A2(G141gat), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n874), .A2(new_n674), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n842), .B1(new_n868), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n869), .A2(new_n873), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n433), .A3(new_n875), .ZN(new_n880));
  INV_X1    g679(.A(new_n842), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n544), .B(new_n844), .C1(new_n864), .C2(new_n866), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n881), .C1(new_n882), .C2(new_n332), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n885), .A3(new_n668), .ZN(new_n886));
  INV_X1    g685(.A(new_n812), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n581), .B1(new_n858), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n437), .B1(new_n863), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n889), .A2(new_n845), .B1(new_n814), .B2(new_n846), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n668), .A2(new_n843), .A3(new_n487), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT59), .B(G148gat), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n874), .A2(new_n674), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n885), .B1(new_n893), .B2(new_n668), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n886), .B(new_n892), .C1(new_n894), .C2(G148gat), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n326), .A3(new_n581), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n867), .A2(new_n581), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n326), .ZN(G1346gat));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n327), .A3(new_n836), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n867), .A2(new_n624), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n327), .ZN(G1347gat));
  AOI21_X1  g700(.A(new_n671), .B1(new_n789), .B2(new_n813), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n435), .A2(new_n433), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n545), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n671), .A2(new_n433), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n442), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n814), .A2(new_n366), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n816), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n814), .A2(KEYINPUT118), .A3(new_n366), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n544), .A2(new_n216), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n906), .B1(new_n914), .B2(new_n915), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n905), .B2(new_n668), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n667), .A2(new_n215), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n914), .B2(new_n918), .ZN(G1349gat));
  OR3_X1    g718(.A1(new_n904), .A2(new_n254), .A3(new_n582), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n581), .B(new_n909), .C1(new_n815), .C2(new_n817), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(new_n256), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT60), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n920), .B(new_n925), .C1(new_n922), .C2(new_n256), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1350gat));
  INV_X1    g726(.A(G190gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n905), .A2(new_n928), .A3(new_n624), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n624), .ZN(new_n930));
  NOR2_X1   g729(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1351gat));
  NAND2_X1  g734(.A1(new_n870), .A2(new_n674), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT125), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n902), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n545), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n890), .A2(new_n683), .A3(new_n908), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n545), .A2(G197gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n938), .A2(new_n943), .A3(new_n668), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n940), .A2(new_n668), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n947), .B(new_n949), .C1(new_n950), .C2(new_n943), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n310), .A3(new_n581), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n908), .A2(new_n683), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n889), .A2(new_n845), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n814), .A2(new_n846), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n581), .B(new_n953), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  AOI21_X1  g758(.A(G218gat), .B1(new_n938), .B2(new_n624), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n624), .A2(G218gat), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n940), .B2(new_n962), .ZN(G1355gat));
endmodule


